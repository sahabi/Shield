module shield(clock, l1, l2, l3, l1__1, l2__1, l3__1);
  input clock;
  input l1;
  input l2;
  input l3;
  output l1__1;
  output l2__1;
  output l3__1;

  wire s0n;
  wire s1n;
  wire s2n;
  wire s3n;
  wire tmp1;
  wire tmp2;
  wire tmp3;
  wire tmp4;
  wire tmp5;
  wire tmp6;
  wire tmp7;
  wire tmp8;
  wire tmp9;
  wire tmp10;
  wire tmp11;
  wire tmp12;
  wire tmp13;
  wire tmp14;
  wire tmp15;
  wire tmp16;
  wire tmp17;
  wire tmp18;
  wire tmp19;
  wire tmp20;
  wire tmp21;
  wire tmp22;
  wire tmp23;
  wire tmp24;
  wire tmp25;
  wire tmp26;
  wire tmp27;
  wire tmp28;
  wire tmp29;
  wire tmp30;
  wire tmp31;
  wire tmp32;
  wire tmp33;
  wire tmp34;
  wire tmp35;
  wire tmp36;
  wire tmp37;
  wire tmp38;
  wire tmp39;
  wire tmp40;
  wire tmp41;
  wire tmp42;
  wire tmp43;
  wire tmp44;
  wire tmp45;
  wire tmp46;
  wire tmp47;
  wire tmp48;
  wire tmp49;
  wire tmp50;
  wire tmp51;
  wire tmp52;
  wire tmp53;
  wire tmp54;
  wire tmp55;
  wire tmp56;
  wire tmp57;
  wire tmp58;
  wire tmp59;
  wire tmp60;
  wire tmp61;
  wire tmp62;
  wire tmp63;
  wire tmp64;
  wire tmp65;
  wire tmp66;
  wire tmp67;
  wire tmp68;
  wire tmp69;
  wire tmp70;
  wire tmp71;
  wire tmp72;
  wire tmp73;
  wire tmp74;
  wire tmp75;
  wire tmp76;
  wire tmp77;
  wire tmp78;
  wire tmp79;
  wire tmp80;
  wire tmp81;
  wire tmp82;
  wire tmp83;
  wire tmp84;
  wire tmp85;
  wire tmp86;
  wire tmp87;

  reg s0;
  reg s1;
  reg s2;
  reg s3;

  assign tmp1 = l1 ? 1 : 0;
  assign l1__1 = tmp1;

  assign tmp4 = l2 ? 1 : 0;
  assign tmp3 = l1 ? tmp4 : 1;
  assign tmp8 = l1 ? 1 : tmp4;
  assign tmp7 = s0 ? tmp8 : tmp3;
  assign tmp10 = ~(l2 ? 1 : 0);
  assign tmp9 = ~(l1 ? 1 : tmp10);
  assign tmp6 = s1 ? tmp7 : tmp9;
  assign tmp12 = s0 ? tmp4 : tmp8;
  assign tmp14 = ~(l1 ? tmp4 : 0);
  assign tmp13 = ~(s0 ? 1 : tmp14);
  assign tmp11 = s1 ? tmp12 : tmp13;
  assign tmp5 = s2 ? tmp6 : tmp11;
  assign tmp2 = s3 ? tmp3 : tmp5;
  assign l2__1 = tmp2;

  assign tmp20 = l2 ? 1 : 0;
  assign tmp19 = ~(l1 ? tmp20 : 1);
  assign tmp18 = s0 ? 1 : tmp19;
  assign tmp22 = l3 ? 1 : 0;
  assign tmp21 = l1 ? tmp22 : 1;
  assign tmp17 = s1 ? tmp18 : tmp21;
  assign tmp27 = ~(l3 ? 1 : 0);
  assign tmp26 = ~(l2 ? 1 : tmp27);
  assign tmp25 = l1 ? 1 : tmp26;
  assign tmp24 = s0 ? tmp25 : 0;
  assign tmp29 = l1 ? 1 : tmp27;
  assign tmp31 = l2 ? 1 : tmp27;
  assign tmp30 = l1 ? tmp31 : 1;
  assign tmp28 = ~(s0 ? tmp29 : tmp30);
  assign tmp23 = s1 ? tmp24 : tmp28;
  assign tmp16 = s2 ? tmp17 : tmp23;
  assign tmp15 = s3 ? 1 : tmp16;
  assign l3__1 = tmp15;

  assign tmp34 = l2 ? 1 : 0;
  assign tmp33 = l1 ? tmp34 : 0;
  assign tmp38 = l1 ? 1 : 0;
  assign tmp37 = s0 ? tmp38 : 0;
  assign tmp36 = s1 ? tmp37 : 0;
  assign tmp40 = s0 ? tmp33 : 0;
  assign tmp39 = s1 ? tmp40 : 0;
  assign tmp35 = s2 ? tmp36 : tmp39;
  assign tmp32 = s3 ? tmp33 : tmp35;
  assign s3n = tmp32;

  assign tmp42 = l1 ? 1 : 0;
  assign tmp48 = l3 ? 1 : 0;
  assign tmp47 = ~(l2 ? 1 : tmp48);
  assign tmp46 = l1 ? 1 : tmp47;
  assign tmp50 = ~(l2 ? 1 : 0);
  assign tmp49 = l1 ? 1 : tmp50;
  assign tmp45 = s0 ? tmp46 : tmp49;
  assign tmp53 = ~(l3 ? 1 : 0);
  assign tmp52 = l1 ? 1 : tmp53;
  assign tmp51 = s0 ? tmp52 : 1;
  assign tmp44 = s1 ? tmp45 : tmp51;
  assign tmp43 = s2 ? tmp42 : tmp44;
  assign tmp41 = ~(s3 ? tmp42 : tmp43);
  assign s2n = tmp41;

  assign tmp56 = l2 ? 1 : 0;
  assign tmp55 = l1 ? tmp56 : 0;
  assign tmp61 = ~(l2 ? 1 : 0);
  assign tmp60 = l1 ? 1 : tmp61;
  assign tmp59 = s0 ? tmp60 : 0;
  assign tmp63 = l3 ? 1 : 0;
  assign tmp62 = ~(l1 ? tmp63 : tmp56);
  assign tmp58 = s1 ? tmp59 : tmp62;
  assign tmp66 = l1 ? tmp56 : tmp61;
  assign tmp67 = ~(l1 ? 1 : tmp56);
  assign tmp65 = s0 ? tmp66 : tmp67;
  assign tmp70 = l2 ? 1 : tmp63;
  assign tmp69 = ~(l1 ? tmp70 : 0);
  assign tmp68 = s0 ? 1 : tmp69;
  assign tmp64 = s1 ? tmp65 : tmp68;
  assign tmp57 = s2 ? tmp58 : tmp64;
  assign tmp54 = ~(s3 ? tmp55 : tmp57);
  assign s1n = tmp54;

  assign tmp73 = l2 ? 1 : 0;
  assign tmp72 = l1 ? tmp73 : 0;
  assign tmp77 = l1 ? 1 : 0;
  assign tmp78 = l1 ? tmp73 : 1;
  assign tmp76 = s0 ? tmp77 : tmp78;
  assign tmp75 = s1 ? tmp76 : 0;
  assign tmp83 = ~(l3 ? 1 : 0);
  assign tmp82 = l2 ? 1 : tmp83;
  assign tmp81 = l1 ? tmp73 : tmp82;
  assign tmp80 = s0 ? tmp81 : 1;
  assign tmp86 = l3 ? 1 : 0;
  assign tmp85 = l1 ? 1 : tmp86;
  assign tmp87 = ~(l1 ? tmp73 : 1);
  assign tmp84 = ~(s0 ? tmp85 : tmp87);
  assign tmp79 = s1 ? tmp80 : tmp84;
  assign tmp74 = s2 ? tmp75 : tmp79;
  assign tmp71 = ~(s3 ? tmp72 : tmp74);
  assign s0n = tmp71;

  initial
   begin
    s0 = 0;
    s1 = 0;
    s2 = 0;
    s3 = 0;
   end

  always @(posedge clock)
   begin
    s0 = s0n;
    s1 = s1n;
    s2 = s2n;
    s3 = s3n;
   end
endmodule

