/**************************************
* Simulation for inputfiles   
*    "inputfiles/uav/map_16_states/map.dfa",
*    "inputfiles/uav/map_16_states/communication.dfa",
*    "inputfiles/uav/map_16_states/roz.dfa"
*
***************************************/

module main;
  // Input of DUT:
  reg clk;
  reg l4;
  reg l3;
  reg l2;
  reg l1;
  
  // Output of the DUT:
  wire l4__1;
  wire l3__1;
  wire l2__1;
  wire l1__1;

  //Instantiate the DUT:
  shield s(clk, l1, l2, l3, l4, l1__1, l2__1, l3__1, l4__1);
  
  // make clock toggle:
  always #5 clk = ~clk;
  
  // Sequence of input stimuli to test with:
  initial begin
    clk = 0;
    l4 = 0;
    l3 = 0;
    l2 = 0;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d", 
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1);

    $display("Go to location 12: 1 -> 6 -> 3 -> 11 -> 12 -> 12 ");    

    //time=11 -------------------------------------------------
    #9
    l4 = 0;
    l3 = 1;
    l2 = 0;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d",  
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1);

    //time=21 -------------------------------------------------
    #9
    l4 = 0;
    l3 = 0;
    l2 = 1;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d",  
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1);
 
    //time=31 -------------------------------------------------
    #9
    l4 = 1;
    l3 = 0;
    l2 = 1;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d", 
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1);

    //time=61 -------------------------------------------------
    #9
    l4 = 1;
    l3 = 0;
    l2 = 1;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d", 
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1); 

    //time=71 -------------------------------------------------
    #9
    l4 = 1;
    l3 = 0;
    l2 = 1;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d (Error by Design, ROZ)",  
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1);

    //time=81 -------------------------------------------------
    #9
    l4 = 1;
    l3 = 1;
    l2 = 0;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d", 
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1); 

    //time=91 -------------------------------------------------
    #9
    l4 = 1;
    l3 = 1;
    l2 = 0;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d%d, loc_shield=%d%d%d%d", 
             $time, 
             l4, l3, l2, l1, l4__1, l3__1, l2__1, l1__1); 

    #1 $finish;         
  end
endmodule


module shield(clock, l1, l2, l3, l4, l1__1, l2__1, l3__1, l4__1, recovery__1, recovery__2);  
  input clock;
  input l1;
  input l2;
  input l3;
  input l4;
  output l1__1;
  output l2__1;
  output l3__1;
  output l4__1;
  output recovery__1;
  output recovery__2;

  wire s0n;
  wire s1n;
  wire s2n;
  wire s3n;
  wire s4n;
  wire s5n;
  wire s6n;
  wire s7n;
  wire s8n;
  wire s9n;
  wire s10n;
  wire s11n;
  wire s12n;
  wire s13n;
  wire s14n;
  wire s15n;
  wire s16n;
  wire s17n;
  wire s18n;
  wire tmp1;
  wire tmp2;
  wire tmp3;
  wire tmp4;
  wire tmp5;
  wire tmp6;
  wire tmp7;
  wire tmp8;
  wire tmp9;
  wire tmp10;
  wire tmp11;
  wire tmp12;
  wire tmp13;
  wire tmp14;
  wire tmp15;
  wire tmp16;
  wire tmp17;
  wire tmp18;
  wire tmp19;
  wire tmp20;
  wire tmp21;
  wire tmp22;
  wire tmp23;
  wire tmp24;
  wire tmp25;
  wire tmp26;
  wire tmp27;
  wire tmp28;
  wire tmp29;
  wire tmp30;
  wire tmp31;
  wire tmp32;
  wire tmp33;
  wire tmp34;
  wire tmp35;
  wire tmp36;
  wire tmp37;
  wire tmp38;
  wire tmp39;
  wire tmp40;
  wire tmp41;
  wire tmp42;
  wire tmp43;
  wire tmp44;
  wire tmp45;
  wire tmp46;
  wire tmp47;
  wire tmp48;
  wire tmp49;
  wire tmp50;
  wire tmp51;
  wire tmp52;
  wire tmp53;
  wire tmp54;
  wire tmp55;
  wire tmp56;
  wire tmp57;
  wire tmp58;
  wire tmp59;
  wire tmp60;
  wire tmp61;
  wire tmp62;
  wire tmp63;
  wire tmp64;
  wire tmp65;
  wire tmp66;
  wire tmp67;
  wire tmp68;
  wire tmp69;
  wire tmp70;
  wire tmp71;
  wire tmp72;
  wire tmp73;
  wire tmp74;
  wire tmp75;
  wire tmp76;
  wire tmp77;
  wire tmp78;
  wire tmp79;
  wire tmp80;
  wire tmp81;
  wire tmp82;
  wire tmp83;
  wire tmp84;
  wire tmp85;
  wire tmp86;
  wire tmp87;
  wire tmp88;
  wire tmp89;
  wire tmp90;
  wire tmp91;
  wire tmp92;
  wire tmp93;
  wire tmp94;
  wire tmp95;
  wire tmp96;
  wire tmp97;
  wire tmp98;
  wire tmp99;
  wire tmp100;
  wire tmp101;
  wire tmp102;
  wire tmp103;
  wire tmp104;
  wire tmp105;
  wire tmp106;
  wire tmp107;
  wire tmp108;
  wire tmp109;
  wire tmp110;
  wire tmp111;
  wire tmp112;
  wire tmp113;
  wire tmp114;
  wire tmp115;
  wire tmp116;
  wire tmp117;
  wire tmp118;
  wire tmp119;
  wire tmp120;
  wire tmp121;
  wire tmp122;
  wire tmp123;
  wire tmp124;
  wire tmp125;
  wire tmp126;
  wire tmp127;
  wire tmp128;
  wire tmp129;
  wire tmp130;
  wire tmp131;
  wire tmp132;
  wire tmp133;
  wire tmp134;
  wire tmp135;
  wire tmp136;
  wire tmp137;
  wire tmp138;
  wire tmp139;
  wire tmp140;
  wire tmp141;
  wire tmp142;
  wire tmp143;
  wire tmp144;
  wire tmp145;
  wire tmp146;
  wire tmp147;
  wire tmp148;
  wire tmp149;
  wire tmp150;
  wire tmp151;
  wire tmp152;
  wire tmp153;
  wire tmp154;
  wire tmp155;
  wire tmp156;
  wire tmp157;
  wire tmp158;
  wire tmp159;
  wire tmp160;
  wire tmp161;
  wire tmp162;
  wire tmp163;
  wire tmp164;
  wire tmp165;
  wire tmp166;
  wire tmp167;
  wire tmp168;
  wire tmp169;
  wire tmp170;
  wire tmp171;
  wire tmp172;
  wire tmp173;
  wire tmp174;
  wire tmp175;
  wire tmp176;
  wire tmp177;
  wire tmp178;
  wire tmp179;
  wire tmp180;
  wire tmp181;
  wire tmp182;
  wire tmp183;
  wire tmp184;
  wire tmp185;
  wire tmp186;
  wire tmp187;
  wire tmp188;
  wire tmp189;
  wire tmp190;
  wire tmp191;
  wire tmp192;
  wire tmp193;
  wire tmp194;
  wire tmp195;
  wire tmp196;
  wire tmp197;
  wire tmp198;
  wire tmp199;
  wire tmp200;
  wire tmp201;
  wire tmp202;
  wire tmp203;
  wire tmp204;
  wire tmp205;
  wire tmp206;
  wire tmp207;
  wire tmp208;
  wire tmp209;
  wire tmp210;
  wire tmp211;
  wire tmp212;
  wire tmp213;
  wire tmp214;
  wire tmp215;
  wire tmp216;
  wire tmp217;
  wire tmp218;
  wire tmp219;
  wire tmp220;
  wire tmp221;
  wire tmp222;
  wire tmp223;
  wire tmp224;
  wire tmp225;
  wire tmp226;
  wire tmp227;
  wire tmp228;
  wire tmp229;
  wire tmp230;
  wire tmp231;
  wire tmp232;
  wire tmp233;
  wire tmp234;
  wire tmp235;
  wire tmp236;
  wire tmp237;
  wire tmp238;
  wire tmp239;
  wire tmp240;
  wire tmp241;
  wire tmp242;
  wire tmp243;
  wire tmp244;
  wire tmp245;
  wire tmp246;
  wire tmp247;
  wire tmp248;
  wire tmp249;
  wire tmp250;
  wire tmp251;
  wire tmp252;
  wire tmp253;
  wire tmp254;
  wire tmp255;
  wire tmp256;
  wire tmp257;
  wire tmp258;
  wire tmp259;
  wire tmp260;
  wire tmp261;
  wire tmp262;
  wire tmp263;
  wire tmp264;
  wire tmp265;
  wire tmp266;
  wire tmp267;
  wire tmp268;
  wire tmp269;
  wire tmp270;
  wire tmp271;
  wire tmp272;
  wire tmp273;
  wire tmp274;
  wire tmp275;
  wire tmp276;
  wire tmp277;
  wire tmp278;
  wire tmp279;
  wire tmp280;
  wire tmp281;
  wire tmp282;
  wire tmp283;
  wire tmp284;
  wire tmp285;
  wire tmp286;
  wire tmp287;
  wire tmp288;
  wire tmp289;
  wire tmp290;
  wire tmp291;
  wire tmp292;
  wire tmp293;
  wire tmp294;
  wire tmp295;
  wire tmp296;
  wire tmp297;
  wire tmp298;
  wire tmp299;
  wire tmp300;
  wire tmp301;
  wire tmp302;
  wire tmp303;
  wire tmp304;
  wire tmp305;
  wire tmp306;
  wire tmp307;
  wire tmp308;
  wire tmp309;
  wire tmp310;
  wire tmp311;
  wire tmp312;
  wire tmp313;
  wire tmp314;
  wire tmp315;
  wire tmp316;
  wire tmp317;
  wire tmp318;
  wire tmp319;
  wire tmp320;
  wire tmp321;
  wire tmp322;
  wire tmp323;
  wire tmp324;
  wire tmp325;
  wire tmp326;
  wire tmp327;
  wire tmp328;
  wire tmp329;
  wire tmp330;
  wire tmp331;
  wire tmp332;
  wire tmp333;
  wire tmp334;
  wire tmp335;
  wire tmp336;
  wire tmp337;
  wire tmp338;
  wire tmp339;
  wire tmp340;
  wire tmp341;
  wire tmp342;
  wire tmp343;
  wire tmp344;
  wire tmp345;
  wire tmp346;
  wire tmp347;
  wire tmp348;
  wire tmp349;
  wire tmp350;
  wire tmp351;
  wire tmp352;
  wire tmp353;
  wire tmp354;
  wire tmp355;
  wire tmp356;
  wire tmp357;
  wire tmp358;
  wire tmp359;
  wire tmp360;
  wire tmp361;
  wire tmp362;
  wire tmp363;
  wire tmp364;
  wire tmp365;
  wire tmp366;
  wire tmp367;
  wire tmp368;
  wire tmp369;
  wire tmp370;
  wire tmp371;
  wire tmp372;
  wire tmp373;
  wire tmp374;
  wire tmp375;
  wire tmp376;
  wire tmp377;
  wire tmp378;
  wire tmp379;
  wire tmp380;
  wire tmp381;
  wire tmp382;
  wire tmp383;
  wire tmp384;
  wire tmp385;
  wire tmp386;
  wire tmp387;
  wire tmp388;
  wire tmp389;
  wire tmp390;
  wire tmp391;
  wire tmp392;
  wire tmp393;
  wire tmp394;
  wire tmp395;
  wire tmp396;
  wire tmp397;
  wire tmp398;
  wire tmp399;
  wire tmp400;
  wire tmp401;
  wire tmp402;
  wire tmp403;
  wire tmp404;
  wire tmp405;
  wire tmp406;
  wire tmp407;
  wire tmp408;
  wire tmp409;
  wire tmp410;
  wire tmp411;
  wire tmp412;
  wire tmp413;
  wire tmp414;
  wire tmp415;
  wire tmp416;
  wire tmp417;
  wire tmp418;
  wire tmp419;
  wire tmp420;
  wire tmp421;
  wire tmp422;
  wire tmp423;
  wire tmp424;
  wire tmp425;
  wire tmp426;
  wire tmp427;
  wire tmp428;
  wire tmp429;
  wire tmp430;
  wire tmp431;
  wire tmp432;
  wire tmp433;
  wire tmp434;
  wire tmp435;
  wire tmp436;
  wire tmp437;
  wire tmp438;
  wire tmp439;
  wire tmp440;
  wire tmp441;
  wire tmp442;
  wire tmp443;
  wire tmp444;
  wire tmp445;
  wire tmp446;
  wire tmp447;
  wire tmp448;
  wire tmp449;
  wire tmp450;
  wire tmp451;
  wire tmp452;
  wire tmp453;
  wire tmp454;
  wire tmp455;
  wire tmp456;
  wire tmp457;
  wire tmp458;
  wire tmp459;
  wire tmp460;
  wire tmp461;
  wire tmp462;
  wire tmp463;
  wire tmp464;
  wire tmp465;
  wire tmp466;
  wire tmp467;
  wire tmp468;
  wire tmp469;
  wire tmp470;
  wire tmp471;
  wire tmp472;
  wire tmp473;
  wire tmp474;
  wire tmp475;
  wire tmp476;
  wire tmp477;
  wire tmp478;
  wire tmp479;
  wire tmp480;
  wire tmp481;
  wire tmp482;
  wire tmp483;
  wire tmp484;
  wire tmp485;
  wire tmp486;
  wire tmp487;
  wire tmp488;
  wire tmp489;
  wire tmp490;
  wire tmp491;
  wire tmp492;
  wire tmp493;
  wire tmp494;
  wire tmp495;
  wire tmp496;
  wire tmp497;
  wire tmp498;
  wire tmp499;
  wire tmp500;
  wire tmp501;
  wire tmp502;
  wire tmp503;
  wire tmp504;
  wire tmp505;
  wire tmp506;
  wire tmp507;
  wire tmp508;
  wire tmp509;
  wire tmp510;
  wire tmp511;
  wire tmp512;
  wire tmp513;
  wire tmp514;
  wire tmp515;
  wire tmp516;
  wire tmp517;
  wire tmp518;
  wire tmp519;
  wire tmp520;
  wire tmp521;
  wire tmp522;
  wire tmp523;
  wire tmp524;
  wire tmp525;
  wire tmp526;
  wire tmp527;
  wire tmp528;
  wire tmp529;
  wire tmp530;
  wire tmp531;
  wire tmp532;
  wire tmp533;
  wire tmp534;
  wire tmp535;
  wire tmp536;
  wire tmp537;
  wire tmp538;
  wire tmp539;
  wire tmp540;
  wire tmp541;
  wire tmp542;
  wire tmp543;
  wire tmp544;
  wire tmp545;
  wire tmp546;
  wire tmp547;
  wire tmp548;
  wire tmp549;
  wire tmp550;
  wire tmp551;
  wire tmp552;
  wire tmp553;
  wire tmp554;
  wire tmp555;
  wire tmp556;
  wire tmp557;
  wire tmp558;
  wire tmp559;
  wire tmp560;
  wire tmp561;
  wire tmp562;
  wire tmp563;
  wire tmp564;
  wire tmp565;
  wire tmp566;
  wire tmp567;
  wire tmp568;
  wire tmp569;
  wire tmp570;
  wire tmp571;
  wire tmp572;
  wire tmp573;
  wire tmp574;
  wire tmp575;
  wire tmp576;
  wire tmp577;
  wire tmp578;
  wire tmp579;
  wire tmp580;
  wire tmp581;
  wire tmp582;
  wire tmp583;
  wire tmp584;
  wire tmp585;
  wire tmp586;
  wire tmp587;
  wire tmp588;
  wire tmp589;
  wire tmp590;
  wire tmp591;
  wire tmp592;
  wire tmp593;
  wire tmp594;
  wire tmp595;
  wire tmp596;
  wire tmp597;
  wire tmp598;
  wire tmp599;
  wire tmp600;
  wire tmp601;
  wire tmp602;
  wire tmp603;
  wire tmp604;
  wire tmp605;
  wire tmp606;
  wire tmp607;
  wire tmp608;
  wire tmp609;
  wire tmp610;
  wire tmp611;
  wire tmp612;
  wire tmp613;
  wire tmp614;
  wire tmp615;
  wire tmp616;
  wire tmp617;
  wire tmp618;
  wire tmp619;
  wire tmp620;
  wire tmp621;
  wire tmp622;
  wire tmp623;
  wire tmp624;
  wire tmp625;
  wire tmp626;
  wire tmp627;
  wire tmp628;
  wire tmp629;
  wire tmp630;
  wire tmp631;
  wire tmp632;
  wire tmp633;
  wire tmp634;
  wire tmp635;
  wire tmp636;
  wire tmp637;
  wire tmp638;
  wire tmp639;
  wire tmp640;
  wire tmp641;
  wire tmp642;
  wire tmp643;
  wire tmp644;
  wire tmp645;
  wire tmp646;
  wire tmp647;
  wire tmp648;
  wire tmp649;
  wire tmp650;
  wire tmp651;
  wire tmp652;
  wire tmp653;
  wire tmp654;
  wire tmp655;
  wire tmp656;
  wire tmp657;
  wire tmp658;
  wire tmp659;
  wire tmp660;
  wire tmp661;
  wire tmp662;
  wire tmp663;
  wire tmp664;
  wire tmp665;
  wire tmp666;
  wire tmp667;
  wire tmp668;
  wire tmp669;
  wire tmp670;
  wire tmp671;
  wire tmp672;
  wire tmp673;
  wire tmp674;
  wire tmp675;
  wire tmp676;
  wire tmp677;
  wire tmp678;
  wire tmp679;
  wire tmp680;
  wire tmp681;
  wire tmp682;
  wire tmp683;
  wire tmp684;
  wire tmp685;
  wire tmp686;
  wire tmp687;
  wire tmp688;
  wire tmp689;
  wire tmp690;
  wire tmp691;
  wire tmp692;
  wire tmp693;
  wire tmp694;
  wire tmp695;
  wire tmp696;
  wire tmp697;
  wire tmp698;
  wire tmp699;
  wire tmp700;
  wire tmp701;
  wire tmp702;
  wire tmp703;
  wire tmp704;
  wire tmp705;
  wire tmp706;
  wire tmp707;
  wire tmp708;
  wire tmp709;
  wire tmp710;
  wire tmp711;
  wire tmp712;
  wire tmp713;
  wire tmp714;
  wire tmp715;
  wire tmp716;
  wire tmp717;
  wire tmp718;
  wire tmp719;
  wire tmp720;
  wire tmp721;
  wire tmp722;
  wire tmp723;
  wire tmp724;
  wire tmp725;
  wire tmp726;
  wire tmp727;
  wire tmp728;
  wire tmp729;
  wire tmp730;
  wire tmp731;
  wire tmp732;
  wire tmp733;
  wire tmp734;
  wire tmp735;
  wire tmp736;
  wire tmp737;
  wire tmp738;
  wire tmp739;
  wire tmp740;
  wire tmp741;
  wire tmp742;
  wire tmp743;
  wire tmp744;
  wire tmp745;
  wire tmp746;
  wire tmp747;
  wire tmp748;
  wire tmp749;
  wire tmp750;
  wire tmp751;
  wire tmp752;
  wire tmp753;
  wire tmp754;
  wire tmp755;
  wire tmp756;
  wire tmp757;
  wire tmp758;
  wire tmp759;
  wire tmp760;
  wire tmp761;
  wire tmp762;
  wire tmp763;
  wire tmp764;
  wire tmp765;
  wire tmp766;
  wire tmp767;
  wire tmp768;
  wire tmp769;
  wire tmp770;
  wire tmp771;
  wire tmp772;
  wire tmp773;
  wire tmp774;
  wire tmp775;
  wire tmp776;
  wire tmp777;
  wire tmp778;
  wire tmp779;
  wire tmp780;
  wire tmp781;
  wire tmp782;
  wire tmp783;
  wire tmp784;
  wire tmp785;
  wire tmp786;
  wire tmp787;
  wire tmp788;
  wire tmp789;
  wire tmp790;
  wire tmp791;
  wire tmp792;
  wire tmp793;
  wire tmp794;
  wire tmp795;
  wire tmp796;
  wire tmp797;
  wire tmp798;
  wire tmp799;
  wire tmp800;
  wire tmp801;
  wire tmp802;
  wire tmp803;
  wire tmp804;
  wire tmp805;
  wire tmp806;
  wire tmp807;
  wire tmp808;
  wire tmp809;
  wire tmp810;
  wire tmp811;
  wire tmp812;
  wire tmp813;
  wire tmp814;
  wire tmp815;
  wire tmp816;
  wire tmp817;
  wire tmp818;
  wire tmp819;
  wire tmp820;
  wire tmp821;
  wire tmp822;
  wire tmp823;
  wire tmp824;
  wire tmp825;
  wire tmp826;
  wire tmp827;
  wire tmp828;
  wire tmp829;
  wire tmp830;
  wire tmp831;
  wire tmp832;
  wire tmp833;
  wire tmp834;
  wire tmp835;
  wire tmp836;
  wire tmp837;
  wire tmp838;
  wire tmp839;
  wire tmp840;
  wire tmp841;
  wire tmp842;
  wire tmp843;
  wire tmp844;
  wire tmp845;
  wire tmp846;
  wire tmp847;
  wire tmp848;
  wire tmp849;
  wire tmp850;
  wire tmp851;
  wire tmp852;
  wire tmp853;
  wire tmp854;
  wire tmp855;
  wire tmp856;
  wire tmp857;
  wire tmp858;
  wire tmp859;
  wire tmp860;
  wire tmp861;
  wire tmp862;
  wire tmp863;
  wire tmp864;
  wire tmp865;
  wire tmp866;
  wire tmp867;
  wire tmp868;
  wire tmp869;
  wire tmp870;
  wire tmp871;
  wire tmp872;
  wire tmp873;
  wire tmp874;
  wire tmp875;
  wire tmp876;
  wire tmp877;
  wire tmp878;
  wire tmp879;
  wire tmp880;
  wire tmp881;
  wire tmp882;
  wire tmp883;
  wire tmp884;
  wire tmp885;
  wire tmp886;
  wire tmp887;
  wire tmp888;
  wire tmp889;
  wire tmp890;
  wire tmp891;
  wire tmp892;
  wire tmp893;
  wire tmp894;
  wire tmp895;
  wire tmp896;
  wire tmp897;
  wire tmp898;
  wire tmp899;
  wire tmp900;
  wire tmp901;
  wire tmp902;
  wire tmp903;
  wire tmp904;
  wire tmp905;
  wire tmp906;
  wire tmp907;
  wire tmp908;
  wire tmp909;
  wire tmp910;
  wire tmp911;
  wire tmp912;
  wire tmp913;
  wire tmp914;
  wire tmp915;
  wire tmp916;
  wire tmp917;
  wire tmp918;
  wire tmp919;
  wire tmp920;
  wire tmp921;
  wire tmp922;
  wire tmp923;
  wire tmp924;
  wire tmp925;
  wire tmp926;
  wire tmp927;
  wire tmp928;
  wire tmp929;
  wire tmp930;
  wire tmp931;
  wire tmp932;
  wire tmp933;
  wire tmp934;
  wire tmp935;
  wire tmp936;
  wire tmp937;
  wire tmp938;
  wire tmp939;
  wire tmp940;
  wire tmp941;
  wire tmp942;
  wire tmp943;
  wire tmp944;
  wire tmp945;
  wire tmp946;
  wire tmp947;
  wire tmp948;
  wire tmp949;
  wire tmp950;
  wire tmp951;
  wire tmp952;
  wire tmp953;
  wire tmp954;
  wire tmp955;
  wire tmp956;
  wire tmp957;
  wire tmp958;
  wire tmp959;
  wire tmp960;
  wire tmp961;
  wire tmp962;
  wire tmp963;
  wire tmp964;
  wire tmp965;
  wire tmp966;
  wire tmp967;
  wire tmp968;
  wire tmp969;
  wire tmp970;
  wire tmp971;
  wire tmp972;
  wire tmp973;
  wire tmp974;
  wire tmp975;
  wire tmp976;
  wire tmp977;
  wire tmp978;
  wire tmp979;
  wire tmp980;
  wire tmp981;
  wire tmp982;
  wire tmp983;
  wire tmp984;
  wire tmp985;
  wire tmp986;
  wire tmp987;
  wire tmp988;
  wire tmp989;
  wire tmp990;
  wire tmp991;
  wire tmp992;
  wire tmp993;
  wire tmp994;
  wire tmp995;
  wire tmp996;
  wire tmp997;
  wire tmp998;
  wire tmp999;
  wire tmp1000;
  wire tmp1001;
  wire tmp1002;
  wire tmp1003;
  wire tmp1004;
  wire tmp1005;
  wire tmp1006;
  wire tmp1007;
  wire tmp1008;
  wire tmp1009;
  wire tmp1010;
  wire tmp1011;
  wire tmp1012;
  wire tmp1013;
  wire tmp1014;
  wire tmp1015;
  wire tmp1016;
  wire tmp1017;
  wire tmp1018;
  wire tmp1019;
  wire tmp1020;
  wire tmp1021;
  wire tmp1022;
  wire tmp1023;
  wire tmp1024;
  wire tmp1025;
  wire tmp1026;
  wire tmp1027;
  wire tmp1028;
  wire tmp1029;
  wire tmp1030;
  wire tmp1031;
  wire tmp1032;
  wire tmp1033;
  wire tmp1034;
  wire tmp1035;
  wire tmp1036;
  wire tmp1037;
  wire tmp1038;
  wire tmp1039;
  wire tmp1040;
  wire tmp1041;
  wire tmp1042;
  wire tmp1043;
  wire tmp1044;
  wire tmp1045;
  wire tmp1046;
  wire tmp1047;
  wire tmp1048;
  wire tmp1049;
  wire tmp1050;
  wire tmp1051;
  wire tmp1052;
  wire tmp1053;
  wire tmp1054;
  wire tmp1055;
  wire tmp1056;
  wire tmp1057;
  wire tmp1058;
  wire tmp1059;
  wire tmp1060;
  wire tmp1061;
  wire tmp1062;
  wire tmp1063;
  wire tmp1064;
  wire tmp1065;
  wire tmp1066;
  wire tmp1067;
  wire tmp1068;
  wire tmp1069;
  wire tmp1070;
  wire tmp1071;
  wire tmp1072;
  wire tmp1073;
  wire tmp1074;
  wire tmp1075;
  wire tmp1076;
  wire tmp1077;
  wire tmp1078;
  wire tmp1079;
  wire tmp1080;
  wire tmp1081;
  wire tmp1082;
  wire tmp1083;
  wire tmp1084;
  wire tmp1085;
  wire tmp1086;
  wire tmp1087;
  wire tmp1088;
  wire tmp1089;
  wire tmp1090;
  wire tmp1091;
  wire tmp1092;
  wire tmp1093;
  wire tmp1094;
  wire tmp1095;
  wire tmp1096;
  wire tmp1097;
  wire tmp1098;
  wire tmp1099;
  wire tmp1100;
  wire tmp1101;
  wire tmp1102;
  wire tmp1103;
  wire tmp1104;
  wire tmp1105;
  wire tmp1106;
  wire tmp1107;
  wire tmp1108;
  wire tmp1109;
  wire tmp1110;
  wire tmp1111;
  wire tmp1112;
  wire tmp1113;
  wire tmp1114;
  wire tmp1115;
  wire tmp1116;
  wire tmp1117;
  wire tmp1118;
  wire tmp1119;
  wire tmp1120;
  wire tmp1121;
  wire tmp1122;
  wire tmp1123;
  wire tmp1124;
  wire tmp1125;
  wire tmp1126;
  wire tmp1127;
  wire tmp1128;
  wire tmp1129;
  wire tmp1130;
  wire tmp1131;
  wire tmp1132;
  wire tmp1133;
  wire tmp1134;
  wire tmp1135;
  wire tmp1136;
  wire tmp1137;
  wire tmp1138;
  wire tmp1139;
  wire tmp1140;
  wire tmp1141;
  wire tmp1142;
  wire tmp1143;
  wire tmp1144;
  wire tmp1145;
  wire tmp1146;
  wire tmp1147;
  wire tmp1148;
  wire tmp1149;
  wire tmp1150;
  wire tmp1151;
  wire tmp1152;
  wire tmp1153;
  wire tmp1154;
  wire tmp1155;
  wire tmp1156;
  wire tmp1157;
  wire tmp1158;
  wire tmp1159;
  wire tmp1160;
  wire tmp1161;
  wire tmp1162;
  wire tmp1163;
  wire tmp1164;
  wire tmp1165;
  wire tmp1166;
  wire tmp1167;
  wire tmp1168;
  wire tmp1169;
  wire tmp1170;
  wire tmp1171;
  wire tmp1172;
  wire tmp1173;
  wire tmp1174;
  wire tmp1175;
  wire tmp1176;
  wire tmp1177;
  wire tmp1178;
  wire tmp1179;
  wire tmp1180;
  wire tmp1181;
  wire tmp1182;
  wire tmp1183;
  wire tmp1184;
  wire tmp1185;
  wire tmp1186;
  wire tmp1187;
  wire tmp1188;
  wire tmp1189;
  wire tmp1190;
  wire tmp1191;
  wire tmp1192;
  wire tmp1193;
  wire tmp1194;
  wire tmp1195;
  wire tmp1196;
  wire tmp1197;
  wire tmp1198;
  wire tmp1199;
  wire tmp1200;
  wire tmp1201;
  wire tmp1202;
  wire tmp1203;
  wire tmp1204;
  wire tmp1205;
  wire tmp1206;
  wire tmp1207;
  wire tmp1208;
  wire tmp1209;
  wire tmp1210;
  wire tmp1211;
  wire tmp1212;
  wire tmp1213;
  wire tmp1214;
  wire tmp1215;
  wire tmp1216;
  wire tmp1217;
  wire tmp1218;
  wire tmp1219;
  wire tmp1220;
  wire tmp1221;
  wire tmp1222;
  wire tmp1223;
  wire tmp1224;
  wire tmp1225;
  wire tmp1226;
  wire tmp1227;
  wire tmp1228;
  wire tmp1229;
  wire tmp1230;
  wire tmp1231;
  wire tmp1232;
  wire tmp1233;
  wire tmp1234;
  wire tmp1235;
  wire tmp1236;
  wire tmp1237;
  wire tmp1238;
  wire tmp1239;
  wire tmp1240;
  wire tmp1241;
  wire tmp1242;
  wire tmp1243;
  wire tmp1244;
  wire tmp1245;
  wire tmp1246;
  wire tmp1247;
  wire tmp1248;
  wire tmp1249;
  wire tmp1250;
  wire tmp1251;
  wire tmp1252;
  wire tmp1253;
  wire tmp1254;
  wire tmp1255;
  wire tmp1256;
  wire tmp1257;
  wire tmp1258;
  wire tmp1259;
  wire tmp1260;
  wire tmp1261;
  wire tmp1262;
  wire tmp1263;
  wire tmp1264;
  wire tmp1265;
  wire tmp1266;
  wire tmp1267;
  wire tmp1268;
  wire tmp1269;
  wire tmp1270;
  wire tmp1271;
  wire tmp1272;
  wire tmp1273;
  wire tmp1274;
  wire tmp1275;
  wire tmp1276;
  wire tmp1277;
  wire tmp1278;
  wire tmp1279;
  wire tmp1280;
  wire tmp1281;
  wire tmp1282;
  wire tmp1283;
  wire tmp1284;
  wire tmp1285;
  wire tmp1286;
  wire tmp1287;
  wire tmp1288;
  wire tmp1289;
  wire tmp1290;
  wire tmp1291;
  wire tmp1292;
  wire tmp1293;
  wire tmp1294;
  wire tmp1295;
  wire tmp1296;
  wire tmp1297;
  wire tmp1298;
  wire tmp1299;
  wire tmp1300;
  wire tmp1301;
  wire tmp1302;
  wire tmp1303;
  wire tmp1304;
  wire tmp1305;
  wire tmp1306;
  wire tmp1307;
  wire tmp1308;
  wire tmp1309;
  wire tmp1310;
  wire tmp1311;
  wire tmp1312;
  wire tmp1313;
  wire tmp1314;
  wire tmp1315;
  wire tmp1316;
  wire tmp1317;
  wire tmp1318;
  wire tmp1319;
  wire tmp1320;
  wire tmp1321;
  wire tmp1322;
  wire tmp1323;
  wire tmp1324;
  wire tmp1325;
  wire tmp1326;
  wire tmp1327;
  wire tmp1328;
  wire tmp1329;
  wire tmp1330;
  wire tmp1331;
  wire tmp1332;
  wire tmp1333;
  wire tmp1334;
  wire tmp1335;
  wire tmp1336;
  wire tmp1337;
  wire tmp1338;
  wire tmp1339;
  wire tmp1340;
  wire tmp1341;
  wire tmp1342;
  wire tmp1343;
  wire tmp1344;
  wire tmp1345;
  wire tmp1346;
  wire tmp1347;
  wire tmp1348;
  wire tmp1349;
  wire tmp1350;
  wire tmp1351;
  wire tmp1352;
  wire tmp1353;
  wire tmp1354;
  wire tmp1355;
  wire tmp1356;
  wire tmp1357;
  wire tmp1358;
  wire tmp1359;
  wire tmp1360;
  wire tmp1361;
  wire tmp1362;
  wire tmp1363;
  wire tmp1364;
  wire tmp1365;
  wire tmp1366;
  wire tmp1367;
  wire tmp1368;
  wire tmp1369;
  wire tmp1370;
  wire tmp1371;
  wire tmp1372;
  wire tmp1373;
  wire tmp1374;
  wire tmp1375;
  wire tmp1376;
  wire tmp1377;
  wire tmp1378;
  wire tmp1379;
  wire tmp1380;
  wire tmp1381;
  wire tmp1382;
  wire tmp1383;
  wire tmp1384;
  wire tmp1385;
  wire tmp1386;
  wire tmp1387;
  wire tmp1388;
  wire tmp1389;
  wire tmp1390;
  wire tmp1391;
  wire tmp1392;
  wire tmp1393;
  wire tmp1394;
  wire tmp1395;
  wire tmp1396;
  wire tmp1397;
  wire tmp1398;
  wire tmp1399;
  wire tmp1400;
  wire tmp1401;
  wire tmp1402;
  wire tmp1403;
  wire tmp1404;
  wire tmp1405;
  wire tmp1406;
  wire tmp1407;
  wire tmp1408;
  wire tmp1409;
  wire tmp1410;
  wire tmp1411;
  wire tmp1412;
  wire tmp1413;
  wire tmp1414;
  wire tmp1415;
  wire tmp1416;
  wire tmp1417;
  wire tmp1418;
  wire tmp1419;
  wire tmp1420;
  wire tmp1421;
  wire tmp1422;
  wire tmp1423;
  wire tmp1424;
  wire tmp1425;
  wire tmp1426;
  wire tmp1427;
  wire tmp1428;
  wire tmp1429;
  wire tmp1430;
  wire tmp1431;
  wire tmp1432;
  wire tmp1433;
  wire tmp1434;
  wire tmp1435;
  wire tmp1436;
  wire tmp1437;
  wire tmp1438;
  wire tmp1439;
  wire tmp1440;
  wire tmp1441;
  wire tmp1442;
  wire tmp1443;
  wire tmp1444;
  wire tmp1445;
  wire tmp1446;
  wire tmp1447;
  wire tmp1448;
  wire tmp1449;
  wire tmp1450;
  wire tmp1451;
  wire tmp1452;
  wire tmp1453;
  wire tmp1454;
  wire tmp1455;
  wire tmp1456;
  wire tmp1457;
  wire tmp1458;
  wire tmp1459;
  wire tmp1460;
  wire tmp1461;
  wire tmp1462;
  wire tmp1463;
  wire tmp1464;
  wire tmp1465;
  wire tmp1466;
  wire tmp1467;
  wire tmp1468;
  wire tmp1469;
  wire tmp1470;
  wire tmp1471;
  wire tmp1472;
  wire tmp1473;
  wire tmp1474;
  wire tmp1475;
  wire tmp1476;
  wire tmp1477;
  wire tmp1478;
  wire tmp1479;
  wire tmp1480;
  wire tmp1481;
  wire tmp1482;
  wire tmp1483;
  wire tmp1484;
  wire tmp1485;
  wire tmp1486;
  wire tmp1487;
  wire tmp1488;
  wire tmp1489;
  wire tmp1490;
  wire tmp1491;
  wire tmp1492;
  wire tmp1493;
  wire tmp1494;
  wire tmp1495;
  wire tmp1496;
  wire tmp1497;
  wire tmp1498;
  wire tmp1499;
  wire tmp1500;
  wire tmp1501;
  wire tmp1502;
  wire tmp1503;
  wire tmp1504;
  wire tmp1505;
  wire tmp1506;
  wire tmp1507;
  wire tmp1508;
  wire tmp1509;
  wire tmp1510;
  wire tmp1511;
  wire tmp1512;
  wire tmp1513;
  wire tmp1514;
  wire tmp1515;
  wire tmp1516;
  wire tmp1517;
  wire tmp1518;
  wire tmp1519;
  wire tmp1520;
  wire tmp1521;
  wire tmp1522;
  wire tmp1523;
  wire tmp1524;
  wire tmp1525;
  wire tmp1526;
  wire tmp1527;
  wire tmp1528;
  wire tmp1529;
  wire tmp1530;
  wire tmp1531;
  wire tmp1532;
  wire tmp1533;
  wire tmp1534;
  wire tmp1535;
  wire tmp1536;
  wire tmp1537;
  wire tmp1538;
  wire tmp1539;
  wire tmp1540;
  wire tmp1541;
  wire tmp1542;
  wire tmp1543;
  wire tmp1544;
  wire tmp1545;
  wire tmp1546;
  wire tmp1547;
  wire tmp1548;
  wire tmp1549;
  wire tmp1550;
  wire tmp1551;
  wire tmp1552;
  wire tmp1553;
  wire tmp1554;
  wire tmp1555;
  wire tmp1556;
  wire tmp1557;
  wire tmp1558;
  wire tmp1559;
  wire tmp1560;
  wire tmp1561;
  wire tmp1562;
  wire tmp1563;
  wire tmp1564;
  wire tmp1565;
  wire tmp1566;
  wire tmp1567;
  wire tmp1568;
  wire tmp1569;
  wire tmp1570;
  wire tmp1571;
  wire tmp1572;
  wire tmp1573;
  wire tmp1574;
  wire tmp1575;
  wire tmp1576;
  wire tmp1577;
  wire tmp1578;
  wire tmp1579;
  wire tmp1580;
  wire tmp1581;
  wire tmp1582;
  wire tmp1583;
  wire tmp1584;
  wire tmp1585;
  wire tmp1586;
  wire tmp1587;
  wire tmp1588;
  wire tmp1589;
  wire tmp1590;
  wire tmp1591;
  wire tmp1592;
  wire tmp1593;
  wire tmp1594;
  wire tmp1595;
  wire tmp1596;
  wire tmp1597;
  wire tmp1598;
  wire tmp1599;
  wire tmp1600;
  wire tmp1601;
  wire tmp1602;
  wire tmp1603;
  wire tmp1604;
  wire tmp1605;
  wire tmp1606;
  wire tmp1607;
  wire tmp1608;
  wire tmp1609;
  wire tmp1610;
  wire tmp1611;
  wire tmp1612;
  wire tmp1613;
  wire tmp1614;
  wire tmp1615;
  wire tmp1616;
  wire tmp1617;
  wire tmp1618;
  wire tmp1619;
  wire tmp1620;
  wire tmp1621;
  wire tmp1622;
  wire tmp1623;
  wire tmp1624;
  wire tmp1625;
  wire tmp1626;
  wire tmp1627;
  wire tmp1628;
  wire tmp1629;
  wire tmp1630;
  wire tmp1631;
  wire tmp1632;
  wire tmp1633;
  wire tmp1634;
  wire tmp1635;
  wire tmp1636;
  wire tmp1637;
  wire tmp1638;
  wire tmp1639;
  wire tmp1640;
  wire tmp1641;
  wire tmp1642;
  wire tmp1643;
  wire tmp1644;
  wire tmp1645;
  wire tmp1646;
  wire tmp1647;
  wire tmp1648;
  wire tmp1649;
  wire tmp1650;
  wire tmp1651;
  wire tmp1652;
  wire tmp1653;
  wire tmp1654;
  wire tmp1655;
  wire tmp1656;
  wire tmp1657;
  wire tmp1658;
  wire tmp1659;
  wire tmp1660;
  wire tmp1661;
  wire tmp1662;
  wire tmp1663;
  wire tmp1664;
  wire tmp1665;
  wire tmp1666;
  wire tmp1667;
  wire tmp1668;
  wire tmp1669;
  wire tmp1670;
  wire tmp1671;
  wire tmp1672;
  wire tmp1673;
  wire tmp1674;
  wire tmp1675;
  wire tmp1676;
  wire tmp1677;
  wire tmp1678;
  wire tmp1679;
  wire tmp1680;
  wire tmp1681;
  wire tmp1682;
  wire tmp1683;
  wire tmp1684;
  wire tmp1685;
  wire tmp1686;
  wire tmp1687;
  wire tmp1688;
  wire tmp1689;
  wire tmp1690;
  wire tmp1691;
  wire tmp1692;
  wire tmp1693;
  wire tmp1694;
  wire tmp1695;
  wire tmp1696;
  wire tmp1697;
  wire tmp1698;
  wire tmp1699;
  wire tmp1700;
  wire tmp1701;
  wire tmp1702;
  wire tmp1703;
  wire tmp1704;
  wire tmp1705;
  wire tmp1706;
  wire tmp1707;
  wire tmp1708;
  wire tmp1709;
  wire tmp1710;
  wire tmp1711;
  wire tmp1712;
  wire tmp1713;
  wire tmp1714;
  wire tmp1715;
  wire tmp1716;
  wire tmp1717;
  wire tmp1718;
  wire tmp1719;
  wire tmp1720;
  wire tmp1721;
  wire tmp1722;
  wire tmp1723;
  wire tmp1724;
  wire tmp1725;
  wire tmp1726;
  wire tmp1727;
  wire tmp1728;
  wire tmp1729;
  wire tmp1730;
  wire tmp1731;
  wire tmp1732;
  wire tmp1733;
  wire tmp1734;
  wire tmp1735;
  wire tmp1736;
  wire tmp1737;
  wire tmp1738;
  wire tmp1739;
  wire tmp1740;
  wire tmp1741;
  wire tmp1742;
  wire tmp1743;
  wire tmp1744;
  wire tmp1745;
  wire tmp1746;
  wire tmp1747;
  wire tmp1748;
  wire tmp1749;
  wire tmp1750;
  wire tmp1751;
  wire tmp1752;
  wire tmp1753;
  wire tmp1754;
  wire tmp1755;
  wire tmp1756;
  wire tmp1757;
  wire tmp1758;
  wire tmp1759;
  wire tmp1760;
  wire tmp1761;
  wire tmp1762;
  wire tmp1763;
  wire tmp1764;
  wire tmp1765;
  wire tmp1766;
  wire tmp1767;
  wire tmp1768;
  wire tmp1769;
  wire tmp1770;
  wire tmp1771;
  wire tmp1772;
  wire tmp1773;
  wire tmp1774;
  wire tmp1775;
  wire tmp1776;
  wire tmp1777;
  wire tmp1778;
  wire tmp1779;
  wire tmp1780;
  wire tmp1781;
  wire tmp1782;
  wire tmp1783;
  wire tmp1784;
  wire tmp1785;
  wire tmp1786;
  wire tmp1787;
  wire tmp1788;
  wire tmp1789;
  wire tmp1790;
  wire tmp1791;
  wire tmp1792;
  wire tmp1793;
  wire tmp1794;
  wire tmp1795;
  wire tmp1796;
  wire tmp1797;
  wire tmp1798;
  wire tmp1799;
  wire tmp1800;
  wire tmp1801;
  wire tmp1802;
  wire tmp1803;
  wire tmp1804;
  wire tmp1805;
  wire tmp1806;
  wire tmp1807;
  wire tmp1808;
  wire tmp1809;
  wire tmp1810;
  wire tmp1811;
  wire tmp1812;
  wire tmp1813;
  wire tmp1814;
  wire tmp1815;
  wire tmp1816;
  wire tmp1817;
  wire tmp1818;
  wire tmp1819;
  wire tmp1820;
  wire tmp1821;
  wire tmp1822;
  wire tmp1823;
  wire tmp1824;
  wire tmp1825;
  wire tmp1826;
  wire tmp1827;
  wire tmp1828;
  wire tmp1829;
  wire tmp1830;
  wire tmp1831;
  wire tmp1832;
  wire tmp1833;
  wire tmp1834;
  wire tmp1835;
  wire tmp1836;
  wire tmp1837;
  wire tmp1838;
  wire tmp1839;
  wire tmp1840;
  wire tmp1841;
  wire tmp1842;
  wire tmp1843;
  wire tmp1844;
  wire tmp1845;
  wire tmp1846;
  wire tmp1847;
  wire tmp1848;
  wire tmp1849;
  wire tmp1850;
  wire tmp1851;
  wire tmp1852;
  wire tmp1853;
  wire tmp1854;
  wire tmp1855;
  wire tmp1856;
  wire tmp1857;
  wire tmp1858;
  wire tmp1859;
  wire tmp1860;
  wire tmp1861;
  wire tmp1862;
  wire tmp1863;
  wire tmp1864;
  wire tmp1865;
  wire tmp1866;
  wire tmp1867;
  wire tmp1868;
  wire tmp1869;
  wire tmp1870;
  wire tmp1871;
  wire tmp1872;
  wire tmp1873;
  wire tmp1874;
  wire tmp1875;
  wire tmp1876;
  wire tmp1877;
  wire tmp1878;
  wire tmp1879;
  wire tmp1880;
  wire tmp1881;
  wire tmp1882;
  wire tmp1883;
  wire tmp1884;
  wire tmp1885;
  wire tmp1886;
  wire tmp1887;
  wire tmp1888;
  wire tmp1889;
  wire tmp1890;
  wire tmp1891;
  wire tmp1892;
  wire tmp1893;
  wire tmp1894;
  wire tmp1895;
  wire tmp1896;
  wire tmp1897;
  wire tmp1898;
  wire tmp1899;
  wire tmp1900;
  wire tmp1901;
  wire tmp1902;
  wire tmp1903;
  wire tmp1904;
  wire tmp1905;
  wire tmp1906;
  wire tmp1907;
  wire tmp1908;
  wire tmp1909;
  wire tmp1910;
  wire tmp1911;
  wire tmp1912;
  wire tmp1913;
  wire tmp1914;
  wire tmp1915;
  wire tmp1916;
  wire tmp1917;
  wire tmp1918;
  wire tmp1919;
  wire tmp1920;
  wire tmp1921;
  wire tmp1922;
  wire tmp1923;
  wire tmp1924;
  wire tmp1925;
  wire tmp1926;
  wire tmp1927;
  wire tmp1928;
  wire tmp1929;
  wire tmp1930;
  wire tmp1931;
  wire tmp1932;
  wire tmp1933;
  wire tmp1934;
  wire tmp1935;
  wire tmp1936;
  wire tmp1937;
  wire tmp1938;
  wire tmp1939;
  wire tmp1940;
  wire tmp1941;
  wire tmp1942;
  wire tmp1943;
  wire tmp1944;
  wire tmp1945;
  wire tmp1946;
  wire tmp1947;
  wire tmp1948;
  wire tmp1949;
  wire tmp1950;
  wire tmp1951;
  wire tmp1952;
  wire tmp1953;
  wire tmp1954;
  wire tmp1955;
  wire tmp1956;
  wire tmp1957;
  wire tmp1958;
  wire tmp1959;
  wire tmp1960;
  wire tmp1961;
  wire tmp1962;
  wire tmp1963;
  wire tmp1964;
  wire tmp1965;
  wire tmp1966;
  wire tmp1967;
  wire tmp1968;
  wire tmp1969;
  wire tmp1970;
  wire tmp1971;
  wire tmp1972;
  wire tmp1973;
  wire tmp1974;
  wire tmp1975;
  wire tmp1976;
  wire tmp1977;
  wire tmp1978;
  wire tmp1979;
  wire tmp1980;
  wire tmp1981;
  wire tmp1982;
  wire tmp1983;
  wire tmp1984;
  wire tmp1985;
  wire tmp1986;
  wire tmp1987;
  wire tmp1988;
  wire tmp1989;
  wire tmp1990;
  wire tmp1991;
  wire tmp1992;
  wire tmp1993;
  wire tmp1994;
  wire tmp1995;
  wire tmp1996;
  wire tmp1997;
  wire tmp1998;
  wire tmp1999;
  wire tmp2000;
  wire tmp2001;
  wire tmp2002;
  wire tmp2003;
  wire tmp2004;
  wire tmp2005;
  wire tmp2006;
  wire tmp2007;
  wire tmp2008;
  wire tmp2009;
  wire tmp2010;
  wire tmp2011;
  wire tmp2012;
  wire tmp2013;
  wire tmp2014;
  wire tmp2015;
  wire tmp2016;
  wire tmp2017;
  wire tmp2018;
  wire tmp2019;
  wire tmp2020;
  wire tmp2021;
  wire tmp2022;
  wire tmp2023;
  wire tmp2024;
  wire tmp2025;
  wire tmp2026;
  wire tmp2027;
  wire tmp2028;
  wire tmp2029;
  wire tmp2030;
  wire tmp2031;
  wire tmp2032;
  wire tmp2033;
  wire tmp2034;
  wire tmp2035;
  wire tmp2036;
  wire tmp2037;
  wire tmp2038;
  wire tmp2039;
  wire tmp2040;
  wire tmp2041;
  wire tmp2042;
  wire tmp2043;
  wire tmp2044;
  wire tmp2045;
  wire tmp2046;
  wire tmp2047;
  wire tmp2048;
  wire tmp2049;
  wire tmp2050;
  wire tmp2051;
  wire tmp2052;
  wire tmp2053;
  wire tmp2054;
  wire tmp2055;
  wire tmp2056;
  wire tmp2057;
  wire tmp2058;
  wire tmp2059;
  wire tmp2060;
  wire tmp2061;
  wire tmp2062;
  wire tmp2063;
  wire tmp2064;
  wire tmp2065;
  wire tmp2066;
  wire tmp2067;
  wire tmp2068;
  wire tmp2069;
  wire tmp2070;
  wire tmp2071;
  wire tmp2072;
  wire tmp2073;
  wire tmp2074;
  wire tmp2075;
  wire tmp2076;
  wire tmp2077;
  wire tmp2078;
  wire tmp2079;
  wire tmp2080;
  wire tmp2081;
  wire tmp2082;
  wire tmp2083;
  wire tmp2084;
  wire tmp2085;
  wire tmp2086;
  wire tmp2087;
  wire tmp2088;
  wire tmp2089;
  wire tmp2090;
  wire tmp2091;
  wire tmp2092;
  wire tmp2093;
  wire tmp2094;
  wire tmp2095;
  wire tmp2096;
  wire tmp2097;
  wire tmp2098;
  wire tmp2099;
  wire tmp2100;
  wire tmp2101;
  wire tmp2102;
  wire tmp2103;
  wire tmp2104;
  wire tmp2105;
  wire tmp2106;
  wire tmp2107;
  wire tmp2108;
  wire tmp2109;
  wire tmp2110;
  wire tmp2111;
  wire tmp2112;
  wire tmp2113;
  wire tmp2114;
  wire tmp2115;
  wire tmp2116;
  wire tmp2117;
  wire tmp2118;
  wire tmp2119;
  wire tmp2120;
  wire tmp2121;
  wire tmp2122;
  wire tmp2123;
  wire tmp2124;
  wire tmp2125;
  wire tmp2126;
  wire tmp2127;
  wire tmp2128;
  wire tmp2129;
  wire tmp2130;
  wire tmp2131;
  wire tmp2132;
  wire tmp2133;
  wire tmp2134;
  wire tmp2135;
  wire tmp2136;
  wire tmp2137;
  wire tmp2138;
  wire tmp2139;
  wire tmp2140;
  wire tmp2141;
  wire tmp2142;
  wire tmp2143;
  wire tmp2144;
  wire tmp2145;
  wire tmp2146;
  wire tmp2147;
  wire tmp2148;
  wire tmp2149;
  wire tmp2150;
  wire tmp2151;
  wire tmp2152;
  wire tmp2153;
  wire tmp2154;
  wire tmp2155;
  wire tmp2156;
  wire tmp2157;
  wire tmp2158;
  wire tmp2159;
  wire tmp2160;
  wire tmp2161;
  wire tmp2162;
  wire tmp2163;
  wire tmp2164;
  wire tmp2165;
  wire tmp2166;
  wire tmp2167;
  wire tmp2168;
  wire tmp2169;
  wire tmp2170;
  wire tmp2171;
  wire tmp2172;
  wire tmp2173;
  wire tmp2174;
  wire tmp2175;
  wire tmp2176;
  wire tmp2177;
  wire tmp2178;
  wire tmp2179;
  wire tmp2180;
  wire tmp2181;
  wire tmp2182;
  wire tmp2183;
  wire tmp2184;
  wire tmp2185;
  wire tmp2186;
  wire tmp2187;
  wire tmp2188;
  wire tmp2189;
  wire tmp2190;
  wire tmp2191;
  wire tmp2192;
  wire tmp2193;
  wire tmp2194;
  wire tmp2195;
  wire tmp2196;
  wire tmp2197;
  wire tmp2198;
  wire tmp2199;
  wire tmp2200;
  wire tmp2201;
  wire tmp2202;
  wire tmp2203;
  wire tmp2204;
  wire tmp2205;
  wire tmp2206;
  wire tmp2207;
  wire tmp2208;
  wire tmp2209;
  wire tmp2210;
  wire tmp2211;
  wire tmp2212;
  wire tmp2213;
  wire tmp2214;
  wire tmp2215;
  wire tmp2216;
  wire tmp2217;
  wire tmp2218;
  wire tmp2219;
  wire tmp2220;
  wire tmp2221;
  wire tmp2222;
  wire tmp2223;
  wire tmp2224;
  wire tmp2225;
  wire tmp2226;
  wire tmp2227;
  wire tmp2228;
  wire tmp2229;
  wire tmp2230;
  wire tmp2231;
  wire tmp2232;
  wire tmp2233;
  wire tmp2234;
  wire tmp2235;
  wire tmp2236;
  wire tmp2237;
  wire tmp2238;
  wire tmp2239;
  wire tmp2240;
  wire tmp2241;
  wire tmp2242;
  wire tmp2243;
  wire tmp2244;
  wire tmp2245;
  wire tmp2246;
  wire tmp2247;
  wire tmp2248;
  wire tmp2249;
  wire tmp2250;
  wire tmp2251;
  wire tmp2252;
  wire tmp2253;
  wire tmp2254;
  wire tmp2255;
  wire tmp2256;
  wire tmp2257;
  wire tmp2258;
  wire tmp2259;
  wire tmp2260;
  wire tmp2261;
  wire tmp2262;
  wire tmp2263;
  wire tmp2264;
  wire tmp2265;
  wire tmp2266;
  wire tmp2267;
  wire tmp2268;
  wire tmp2269;
  wire tmp2270;
  wire tmp2271;
  wire tmp2272;
  wire tmp2273;
  wire tmp2274;
  wire tmp2275;
  wire tmp2276;
  wire tmp2277;
  wire tmp2278;
  wire tmp2279;
  wire tmp2280;
  wire tmp2281;
  wire tmp2282;
  wire tmp2283;
  wire tmp2284;
  wire tmp2285;
  wire tmp2286;
  wire tmp2287;
  wire tmp2288;
  wire tmp2289;
  wire tmp2290;
  wire tmp2291;
  wire tmp2292;
  wire tmp2293;
  wire tmp2294;
  wire tmp2295;
  wire tmp2296;
  wire tmp2297;
  wire tmp2298;
  wire tmp2299;
  wire tmp2300;
  wire tmp2301;
  wire tmp2302;
  wire tmp2303;
  wire tmp2304;
  wire tmp2305;
  wire tmp2306;
  wire tmp2307;
  wire tmp2308;
  wire tmp2309;
  wire tmp2310;
  wire tmp2311;
  wire tmp2312;
  wire tmp2313;
  wire tmp2314;
  wire tmp2315;
  wire tmp2316;
  wire tmp2317;
  wire tmp2318;
  wire tmp2319;
  wire tmp2320;
  wire tmp2321;
  wire tmp2322;
  wire tmp2323;
  wire tmp2324;
  wire tmp2325;
  wire tmp2326;
  wire tmp2327;
  wire tmp2328;
  wire tmp2329;
  wire tmp2330;
  wire tmp2331;
  wire tmp2332;
  wire tmp2333;
  wire tmp2334;
  wire tmp2335;
  wire tmp2336;
  wire tmp2337;
  wire tmp2338;
  wire tmp2339;
  wire tmp2340;
  wire tmp2341;
  wire tmp2342;
  wire tmp2343;
  wire tmp2344;
  wire tmp2345;
  wire tmp2346;
  wire tmp2347;
  wire tmp2348;
  wire tmp2349;
  wire tmp2350;
  wire tmp2351;
  wire tmp2352;
  wire tmp2353;
  wire tmp2354;
  wire tmp2355;
  wire tmp2356;
  wire tmp2357;
  wire tmp2358;
  wire tmp2359;
  wire tmp2360;
  wire tmp2361;
  wire tmp2362;
  wire tmp2363;
  wire tmp2364;
  wire tmp2365;
  wire tmp2366;
  wire tmp2367;
  wire tmp2368;
  wire tmp2369;
  wire tmp2370;
  wire tmp2371;
  wire tmp2372;
  wire tmp2373;
  wire tmp2374;
  wire tmp2375;
  wire tmp2376;
  wire tmp2377;
  wire tmp2378;
  wire tmp2379;
  wire tmp2380;
  wire tmp2381;
  wire tmp2382;
  wire tmp2383;
  wire tmp2384;
  wire tmp2385;
  wire tmp2386;
  wire tmp2387;
  wire tmp2388;
  wire tmp2389;
  wire tmp2390;
  wire tmp2391;
  wire tmp2392;
  wire tmp2393;
  wire tmp2394;
  wire tmp2395;
  wire tmp2396;
  wire tmp2397;
  wire tmp2398;
  wire tmp2399;
  wire tmp2400;
  wire tmp2401;
  wire tmp2402;
  wire tmp2403;
  wire tmp2404;
  wire tmp2405;
  wire tmp2406;
  wire tmp2407;
  wire tmp2408;
  wire tmp2409;
  wire tmp2410;
  wire tmp2411;
  wire tmp2412;
  wire tmp2413;
  wire tmp2414;
  wire tmp2415;
  wire tmp2416;
  wire tmp2417;
  wire tmp2418;
  wire tmp2419;
  wire tmp2420;
  wire tmp2421;
  wire tmp2422;
  wire tmp2423;
  wire tmp2424;
  wire tmp2425;
  wire tmp2426;
  wire tmp2427;
  wire tmp2428;
  wire tmp2429;
  wire tmp2430;
  wire tmp2431;
  wire tmp2432;
  wire tmp2433;
  wire tmp2434;
  wire tmp2435;
  wire tmp2436;
  wire tmp2437;
  wire tmp2438;
  wire tmp2439;
  wire tmp2440;
  wire tmp2441;
  wire tmp2442;
  wire tmp2443;
  wire tmp2444;
  wire tmp2445;
  wire tmp2446;
  wire tmp2447;
  wire tmp2448;
  wire tmp2449;
  wire tmp2450;
  wire tmp2451;
  wire tmp2452;
  wire tmp2453;
  wire tmp2454;
  wire tmp2455;
  wire tmp2456;
  wire tmp2457;
  wire tmp2458;
  wire tmp2459;
  wire tmp2460;
  wire tmp2461;
  wire tmp2462;
  wire tmp2463;
  wire tmp2464;
  wire tmp2465;
  wire tmp2466;
  wire tmp2467;
  wire tmp2468;
  wire tmp2469;
  wire tmp2470;
  wire tmp2471;
  wire tmp2472;
  wire tmp2473;
  wire tmp2474;
  wire tmp2475;
  wire tmp2476;
  wire tmp2477;
  wire tmp2478;
  wire tmp2479;
  wire tmp2480;
  wire tmp2481;
  wire tmp2482;
  wire tmp2483;
  wire tmp2484;
  wire tmp2485;
  wire tmp2486;
  wire tmp2487;
  wire tmp2488;
  wire tmp2489;
  wire tmp2490;
  wire tmp2491;
  wire tmp2492;
  wire tmp2493;
  wire tmp2494;
  wire tmp2495;
  wire tmp2496;
  wire tmp2497;
  wire tmp2498;
  wire tmp2499;
  wire tmp2500;
  wire tmp2501;
  wire tmp2502;
  wire tmp2503;
  wire tmp2504;
  wire tmp2505;
  wire tmp2506;
  wire tmp2507;
  wire tmp2508;
  wire tmp2509;
  wire tmp2510;
  wire tmp2511;
  wire tmp2512;
  wire tmp2513;
  wire tmp2514;
  wire tmp2515;
  wire tmp2516;
  wire tmp2517;
  wire tmp2518;
  wire tmp2519;
  wire tmp2520;
  wire tmp2521;
  wire tmp2522;
  wire tmp2523;
  wire tmp2524;
  wire tmp2525;
  wire tmp2526;
  wire tmp2527;
  wire tmp2528;
  wire tmp2529;
  wire tmp2530;
  wire tmp2531;
  wire tmp2532;
  wire tmp2533;
  wire tmp2534;
  wire tmp2535;
  wire tmp2536;
  wire tmp2537;
  wire tmp2538;
  wire tmp2539;
  wire tmp2540;
  wire tmp2541;
  wire tmp2542;
  wire tmp2543;
  wire tmp2544;
  wire tmp2545;
  wire tmp2546;
  wire tmp2547;
  wire tmp2548;
  wire tmp2549;
  wire tmp2550;
  wire tmp2551;
  wire tmp2552;
  wire tmp2553;
  wire tmp2554;
  wire tmp2555;
  wire tmp2556;
  wire tmp2557;
  wire tmp2558;
  wire tmp2559;
  wire tmp2560;
  wire tmp2561;
  wire tmp2562;
  wire tmp2563;
  wire tmp2564;
  wire tmp2565;
  wire tmp2566;
  wire tmp2567;
  wire tmp2568;
  wire tmp2569;
  wire tmp2570;
  wire tmp2571;
  wire tmp2572;
  wire tmp2573;
  wire tmp2574;
  wire tmp2575;
  wire tmp2576;
  wire tmp2577;
  wire tmp2578;
  wire tmp2579;
  wire tmp2580;
  wire tmp2581;
  wire tmp2582;
  wire tmp2583;
  wire tmp2584;
  wire tmp2585;
  wire tmp2586;
  wire tmp2587;
  wire tmp2588;
  wire tmp2589;
  wire tmp2590;
  wire tmp2591;
  wire tmp2592;
  wire tmp2593;
  wire tmp2594;
  wire tmp2595;
  wire tmp2596;
  wire tmp2597;
  wire tmp2598;
  wire tmp2599;
  wire tmp2600;
  wire tmp2601;
  wire tmp2602;
  wire tmp2603;
  wire tmp2604;
  wire tmp2605;
  wire tmp2606;
  wire tmp2607;
  wire tmp2608;
  wire tmp2609;
  wire tmp2610;
  wire tmp2611;
  wire tmp2612;
  wire tmp2613;
  wire tmp2614;
  wire tmp2615;
  wire tmp2616;
  wire tmp2617;
  wire tmp2618;
  wire tmp2619;
  wire tmp2620;
  wire tmp2621;
  wire tmp2622;
  wire tmp2623;
  wire tmp2624;
  wire tmp2625;
  wire tmp2626;
  wire tmp2627;
  wire tmp2628;
  wire tmp2629;
  wire tmp2630;
  wire tmp2631;
  wire tmp2632;
  wire tmp2633;
  wire tmp2634;
  wire tmp2635;
  wire tmp2636;
  wire tmp2637;
  wire tmp2638;
  wire tmp2639;
  wire tmp2640;
  wire tmp2641;
  wire tmp2642;
  wire tmp2643;
  wire tmp2644;
  wire tmp2645;
  wire tmp2646;
  wire tmp2647;
  wire tmp2648;
  wire tmp2649;
  wire tmp2650;
  wire tmp2651;
  wire tmp2652;
  wire tmp2653;
  wire tmp2654;
  wire tmp2655;
  wire tmp2656;
  wire tmp2657;
  wire tmp2658;
  wire tmp2659;
  wire tmp2660;
  wire tmp2661;
  wire tmp2662;
  wire tmp2663;
  wire tmp2664;
  wire tmp2665;
  wire tmp2666;
  wire tmp2667;
  wire tmp2668;
  wire tmp2669;
  wire tmp2670;
  wire tmp2671;
  wire tmp2672;
  wire tmp2673;
  wire tmp2674;
  wire tmp2675;
  wire tmp2676;
  wire tmp2677;
  wire tmp2678;
  wire tmp2679;
  wire tmp2680;
  wire tmp2681;
  wire tmp2682;
  wire tmp2683;
  wire tmp2684;
  wire tmp2685;
  wire tmp2686;
  wire tmp2687;
  wire tmp2688;
  wire tmp2689;
  wire tmp2690;
  wire tmp2691;
  wire tmp2692;
  wire tmp2693;
  wire tmp2694;
  wire tmp2695;
  wire tmp2696;
  wire tmp2697;
  wire tmp2698;
  wire tmp2699;
  wire tmp2700;
  wire tmp2701;
  wire tmp2702;
  wire tmp2703;
  wire tmp2704;
  wire tmp2705;
  wire tmp2706;
  wire tmp2707;
  wire tmp2708;
  wire tmp2709;
  wire tmp2710;
  wire tmp2711;
  wire tmp2712;
  wire tmp2713;
  wire tmp2714;
  wire tmp2715;
  wire tmp2716;
  wire tmp2717;
  wire tmp2718;
  wire tmp2719;
  wire tmp2720;
  wire tmp2721;
  wire tmp2722;
  wire tmp2723;
  wire tmp2724;
  wire tmp2725;
  wire tmp2726;
  wire tmp2727;
  wire tmp2728;
  wire tmp2729;
  wire tmp2730;
  wire tmp2731;
  wire tmp2732;
  wire tmp2733;
  wire tmp2734;
  wire tmp2735;
  wire tmp2736;
  wire tmp2737;
  wire tmp2738;
  wire tmp2739;
  wire tmp2740;
  wire tmp2741;
  wire tmp2742;
  wire tmp2743;
  wire tmp2744;
  wire tmp2745;
  wire tmp2746;
  wire tmp2747;
  wire tmp2748;
  wire tmp2749;
  wire tmp2750;
  wire tmp2751;
  wire tmp2752;
  wire tmp2753;
  wire tmp2754;
  wire tmp2755;
  wire tmp2756;
  wire tmp2757;
  wire tmp2758;
  wire tmp2759;
  wire tmp2760;
  wire tmp2761;
  wire tmp2762;
  wire tmp2763;
  wire tmp2764;
  wire tmp2765;
  wire tmp2766;
  wire tmp2767;
  wire tmp2768;
  wire tmp2769;
  wire tmp2770;
  wire tmp2771;
  wire tmp2772;
  wire tmp2773;
  wire tmp2774;
  wire tmp2775;
  wire tmp2776;
  wire tmp2777;
  wire tmp2778;
  wire tmp2779;
  wire tmp2780;
  wire tmp2781;
  wire tmp2782;
  wire tmp2783;
  wire tmp2784;
  wire tmp2785;
  wire tmp2786;
  wire tmp2787;
  wire tmp2788;
  wire tmp2789;
  wire tmp2790;
  wire tmp2791;
  wire tmp2792;
  wire tmp2793;
  wire tmp2794;
  wire tmp2795;
  wire tmp2796;
  wire tmp2797;
  wire tmp2798;
  wire tmp2799;
  wire tmp2800;
  wire tmp2801;
  wire tmp2802;
  wire tmp2803;
  wire tmp2804;
  wire tmp2805;
  wire tmp2806;
  wire tmp2807;
  wire tmp2808;
  wire tmp2809;
  wire tmp2810;
  wire tmp2811;
  wire tmp2812;
  wire tmp2813;
  wire tmp2814;
  wire tmp2815;
  wire tmp2816;
  wire tmp2817;
  wire tmp2818;
  wire tmp2819;
  wire tmp2820;
  wire tmp2821;
  wire tmp2822;
  wire tmp2823;
  wire tmp2824;
  wire tmp2825;
  wire tmp2826;
  wire tmp2827;
  wire tmp2828;
  wire tmp2829;
  wire tmp2830;
  wire tmp2831;
  wire tmp2832;
  wire tmp2833;
  wire tmp2834;
  wire tmp2835;
  wire tmp2836;
  wire tmp2837;
  wire tmp2838;
  wire tmp2839;
  wire tmp2840;
  wire tmp2841;
  wire tmp2842;
  wire tmp2843;
  wire tmp2844;
  wire tmp2845;
  wire tmp2846;
  wire tmp2847;
  wire tmp2848;
  wire tmp2849;
  wire tmp2850;
  wire tmp2851;
  wire tmp2852;
  wire tmp2853;
  wire tmp2854;
  wire tmp2855;
  wire tmp2856;
  wire tmp2857;
  wire tmp2858;
  wire tmp2859;
  wire tmp2860;
  wire tmp2861;
  wire tmp2862;
  wire tmp2863;
  wire tmp2864;
  wire tmp2865;
  wire tmp2866;
  wire tmp2867;
  wire tmp2868;
  wire tmp2869;
  wire tmp2870;
  wire tmp2871;
  wire tmp2872;
  wire tmp2873;
  wire tmp2874;
  wire tmp2875;
  wire tmp2876;
  wire tmp2877;
  wire tmp2878;
  wire tmp2879;
  wire tmp2880;
  wire tmp2881;
  wire tmp2882;
  wire tmp2883;
  wire tmp2884;
  wire tmp2885;
  wire tmp2886;
  wire tmp2887;
  wire tmp2888;
  wire tmp2889;
  wire tmp2890;
  wire tmp2891;
  wire tmp2892;
  wire tmp2893;
  wire tmp2894;
  wire tmp2895;
  wire tmp2896;
  wire tmp2897;
  wire tmp2898;
  wire tmp2899;
  wire tmp2900;
  wire tmp2901;
  wire tmp2902;
  wire tmp2903;
  wire tmp2904;
  wire tmp2905;
  wire tmp2906;
  wire tmp2907;
  wire tmp2908;
  wire tmp2909;
  wire tmp2910;
  wire tmp2911;
  wire tmp2912;
  wire tmp2913;
  wire tmp2914;
  wire tmp2915;
  wire tmp2916;
  wire tmp2917;
  wire tmp2918;
  wire tmp2919;
  wire tmp2920;
  wire tmp2921;
  wire tmp2922;
  wire tmp2923;
  wire tmp2924;
  wire tmp2925;
  wire tmp2926;
  wire tmp2927;
  wire tmp2928;
  wire tmp2929;
  wire tmp2930;
  wire tmp2931;
  wire tmp2932;
  wire tmp2933;
  wire tmp2934;
  wire tmp2935;
  wire tmp2936;
  wire tmp2937;
  wire tmp2938;
  wire tmp2939;
  wire tmp2940;
  wire tmp2941;
  wire tmp2942;
  wire tmp2943;
  wire tmp2944;
  wire tmp2945;
  wire tmp2946;
  wire tmp2947;
  wire tmp2948;
  wire tmp2949;
  wire tmp2950;
  wire tmp2951;
  wire tmp2952;
  wire tmp2953;
  wire tmp2954;
  wire tmp2955;
  wire tmp2956;
  wire tmp2957;
  wire tmp2958;
  wire tmp2959;
  wire tmp2960;
  wire tmp2961;
  wire tmp2962;
  wire tmp2963;
  wire tmp2964;
  wire tmp2965;
  wire tmp2966;
  wire tmp2967;
  wire tmp2968;
  wire tmp2969;
  wire tmp2970;
  wire tmp2971;
  wire tmp2972;
  wire tmp2973;
  wire tmp2974;
  wire tmp2975;
  wire tmp2976;
  wire tmp2977;
  wire tmp2978;
  wire tmp2979;
  wire tmp2980;
  wire tmp2981;
  wire tmp2982;
  wire tmp2983;
  wire tmp2984;
  wire tmp2985;
  wire tmp2986;
  wire tmp2987;
  wire tmp2988;
  wire tmp2989;
  wire tmp2990;
  wire tmp2991;
  wire tmp2992;
  wire tmp2993;
  wire tmp2994;
  wire tmp2995;
  wire tmp2996;
  wire tmp2997;
  wire tmp2998;
  wire tmp2999;
  wire tmp3000;
  wire tmp3001;
  wire tmp3002;
  wire tmp3003;
  wire tmp3004;
  wire tmp3005;
  wire tmp3006;
  wire tmp3007;
  wire tmp3008;
  wire tmp3009;
  wire tmp3010;
  wire tmp3011;
  wire tmp3012;
  wire tmp3013;
  wire tmp3014;
  wire tmp3015;
  wire tmp3016;
  wire tmp3017;
  wire tmp3018;
  wire tmp3019;
  wire tmp3020;
  wire tmp3021;
  wire tmp3022;
  wire tmp3023;
  wire tmp3024;
  wire tmp3025;
  wire tmp3026;
  wire tmp3027;
  wire tmp3028;
  wire tmp3029;
  wire tmp3030;
  wire tmp3031;
  wire tmp3032;
  wire tmp3033;
  wire tmp3034;
  wire tmp3035;
  wire tmp3036;
  wire tmp3037;
  wire tmp3038;
  wire tmp3039;
  wire tmp3040;
  wire tmp3041;
  wire tmp3042;
  wire tmp3043;
  wire tmp3044;
  wire tmp3045;
  wire tmp3046;
  wire tmp3047;
  wire tmp3048;
  wire tmp3049;
  wire tmp3050;
  wire tmp3051;
  wire tmp3052;
  wire tmp3053;
  wire tmp3054;
  wire tmp3055;
  wire tmp3056;
  wire tmp3057;
  wire tmp3058;
  wire tmp3059;
  wire tmp3060;
  wire tmp3061;
  wire tmp3062;
  wire tmp3063;
  wire tmp3064;
  wire tmp3065;
  wire tmp3066;
  wire tmp3067;
  wire tmp3068;
  wire tmp3069;
  wire tmp3070;
  wire tmp3071;
  wire tmp3072;
  wire tmp3073;
  wire tmp3074;
  wire tmp3075;
  wire tmp3076;
  wire tmp3077;
  wire tmp3078;
  wire tmp3079;
  wire tmp3080;
  wire tmp3081;
  wire tmp3082;
  wire tmp3083;
  wire tmp3084;
  wire tmp3085;
  wire tmp3086;
  wire tmp3087;
  wire tmp3088;
  wire tmp3089;
  wire tmp3090;
  wire tmp3091;
  wire tmp3092;
  wire tmp3093;
  wire tmp3094;
  wire tmp3095;
  wire tmp3096;
  wire tmp3097;
  wire tmp3098;
  wire tmp3099;
  wire tmp3100;
  wire tmp3101;
  wire tmp3102;
  wire tmp3103;
  wire tmp3104;
  wire tmp3105;
  wire tmp3106;
  wire tmp3107;
  wire tmp3108;
  wire tmp3109;
  wire tmp3110;
  wire tmp3111;
  wire tmp3112;
  wire tmp3113;
  wire tmp3114;
  wire tmp3115;
  wire tmp3116;
  wire tmp3117;
  wire tmp3118;
  wire tmp3119;
  wire tmp3120;
  wire tmp3121;
  wire tmp3122;
  wire tmp3123;
  wire tmp3124;
  wire tmp3125;
  wire tmp3126;
  wire tmp3127;
  wire tmp3128;
  wire tmp3129;
  wire tmp3130;
  wire tmp3131;
  wire tmp3132;
  wire tmp3133;
  wire tmp3134;
  wire tmp3135;
  wire tmp3136;
  wire tmp3137;
  wire tmp3138;
  wire tmp3139;
  wire tmp3140;
  wire tmp3141;
  wire tmp3142;
  wire tmp3143;
  wire tmp3144;
  wire tmp3145;
  wire tmp3146;
  wire tmp3147;
  wire tmp3148;
  wire tmp3149;
  wire tmp3150;
  wire tmp3151;
  wire tmp3152;
  wire tmp3153;
  wire tmp3154;
  wire tmp3155;
  wire tmp3156;
  wire tmp3157;
  wire tmp3158;
  wire tmp3159;
  wire tmp3160;
  wire tmp3161;
  wire tmp3162;
  wire tmp3163;
  wire tmp3164;
  wire tmp3165;
  wire tmp3166;
  wire tmp3167;
  wire tmp3168;
  wire tmp3169;
  wire tmp3170;
  wire tmp3171;
  wire tmp3172;
  wire tmp3173;
  wire tmp3174;
  wire tmp3175;
  wire tmp3176;
  wire tmp3177;
  wire tmp3178;
  wire tmp3179;
  wire tmp3180;
  wire tmp3181;
  wire tmp3182;
  wire tmp3183;
  wire tmp3184;
  wire tmp3185;
  wire tmp3186;
  wire tmp3187;
  wire tmp3188;
  wire tmp3189;
  wire tmp3190;
  wire tmp3191;
  wire tmp3192;
  wire tmp3193;
  wire tmp3194;
  wire tmp3195;
  wire tmp3196;
  wire tmp3197;
  wire tmp3198;
  wire tmp3199;
  wire tmp3200;
  wire tmp3201;
  wire tmp3202;
  wire tmp3203;
  wire tmp3204;
  wire tmp3205;
  wire tmp3206;
  wire tmp3207;
  wire tmp3208;
  wire tmp3209;
  wire tmp3210;
  wire tmp3211;
  wire tmp3212;
  wire tmp3213;
  wire tmp3214;
  wire tmp3215;
  wire tmp3216;
  wire tmp3217;
  wire tmp3218;
  wire tmp3219;
  wire tmp3220;
  wire tmp3221;
  wire tmp3222;
  wire tmp3223;
  wire tmp3224;
  wire tmp3225;
  wire tmp3226;
  wire tmp3227;
  wire tmp3228;
  wire tmp3229;
  wire tmp3230;
  wire tmp3231;
  wire tmp3232;
  wire tmp3233;
  wire tmp3234;
  wire tmp3235;
  wire tmp3236;
  wire tmp3237;
  wire tmp3238;
  wire tmp3239;
  wire tmp3240;
  wire tmp3241;
  wire tmp3242;
  wire tmp3243;
  wire tmp3244;
  wire tmp3245;
  wire tmp3246;
  wire tmp3247;
  wire tmp3248;
  wire tmp3249;
  wire tmp3250;
  wire tmp3251;
  wire tmp3252;
  wire tmp3253;
  wire tmp3254;
  wire tmp3255;
  wire tmp3256;
  wire tmp3257;
  wire tmp3258;
  wire tmp3259;
  wire tmp3260;
  wire tmp3261;
  wire tmp3262;
  wire tmp3263;
  wire tmp3264;
  wire tmp3265;
  wire tmp3266;
  wire tmp3267;
  wire tmp3268;
  wire tmp3269;
  wire tmp3270;
  wire tmp3271;
  wire tmp3272;
  wire tmp3273;
  wire tmp3274;
  wire tmp3275;
  wire tmp3276;
  wire tmp3277;
  wire tmp3278;
  wire tmp3279;
  wire tmp3280;
  wire tmp3281;
  wire tmp3282;
  wire tmp3283;
  wire tmp3284;
  wire tmp3285;
  wire tmp3286;
  wire tmp3287;
  wire tmp3288;
  wire tmp3289;
  wire tmp3290;
  wire tmp3291;
  wire tmp3292;
  wire tmp3293;
  wire tmp3294;
  wire tmp3295;
  wire tmp3296;
  wire tmp3297;
  wire tmp3298;
  wire tmp3299;
  wire tmp3300;
  wire tmp3301;
  wire tmp3302;
  wire tmp3303;
  wire tmp3304;
  wire tmp3305;
  wire tmp3306;
  wire tmp3307;
  wire tmp3308;
  wire tmp3309;
  wire tmp3310;
  wire tmp3311;
  wire tmp3312;
  wire tmp3313;
  wire tmp3314;
  wire tmp3315;
  wire tmp3316;
  wire tmp3317;
  wire tmp3318;
  wire tmp3319;
  wire tmp3320;
  wire tmp3321;
  wire tmp3322;
  wire tmp3323;
  wire tmp3324;
  wire tmp3325;
  wire tmp3326;
  wire tmp3327;
  wire tmp3328;
  wire tmp3329;
  wire tmp3330;
  wire tmp3331;
  wire tmp3332;
  wire tmp3333;
  wire tmp3334;
  wire tmp3335;
  wire tmp3336;
  wire tmp3337;
  wire tmp3338;
  wire tmp3339;
  wire tmp3340;
  wire tmp3341;
  wire tmp3342;
  wire tmp3343;
  wire tmp3344;
  wire tmp3345;
  wire tmp3346;
  wire tmp3347;
  wire tmp3348;
  wire tmp3349;
  wire tmp3350;
  wire tmp3351;
  wire tmp3352;
  wire tmp3353;
  wire tmp3354;
  wire tmp3355;
  wire tmp3356;
  wire tmp3357;
  wire tmp3358;
  wire tmp3359;
  wire tmp3360;
  wire tmp3361;
  wire tmp3362;
  wire tmp3363;
  wire tmp3364;
  wire tmp3365;
  wire tmp3366;
  wire tmp3367;
  wire tmp3368;
  wire tmp3369;
  wire tmp3370;
  wire tmp3371;
  wire tmp3372;
  wire tmp3373;
  wire tmp3374;
  wire tmp3375;
  wire tmp3376;
  wire tmp3377;
  wire tmp3378;
  wire tmp3379;
  wire tmp3380;
  wire tmp3381;
  wire tmp3382;
  wire tmp3383;
  wire tmp3384;
  wire tmp3385;
  wire tmp3386;
  wire tmp3387;
  wire tmp3388;
  wire tmp3389;
  wire tmp3390;
  wire tmp3391;
  wire tmp3392;
  wire tmp3393;
  wire tmp3394;
  wire tmp3395;
  wire tmp3396;
  wire tmp3397;
  wire tmp3398;
  wire tmp3399;
  wire tmp3400;
  wire tmp3401;
  wire tmp3402;
  wire tmp3403;
  wire tmp3404;
  wire tmp3405;
  wire tmp3406;
  wire tmp3407;
  wire tmp3408;
  wire tmp3409;
  wire tmp3410;
  wire tmp3411;
  wire tmp3412;
  wire tmp3413;
  wire tmp3414;
  wire tmp3415;
  wire tmp3416;
  wire tmp3417;
  wire tmp3418;
  wire tmp3419;
  wire tmp3420;
  wire tmp3421;
  wire tmp3422;
  wire tmp3423;
  wire tmp3424;
  wire tmp3425;
  wire tmp3426;
  wire tmp3427;
  wire tmp3428;
  wire tmp3429;
  wire tmp3430;
  wire tmp3431;
  wire tmp3432;
  wire tmp3433;
  wire tmp3434;
  wire tmp3435;
  wire tmp3436;
  wire tmp3437;
  wire tmp3438;
  wire tmp3439;
  wire tmp3440;
  wire tmp3441;
  wire tmp3442;
  wire tmp3443;
  wire tmp3444;
  wire tmp3445;
  wire tmp3446;
  wire tmp3447;
  wire tmp3448;
  wire tmp3449;
  wire tmp3450;
  wire tmp3451;
  wire tmp3452;
  wire tmp3453;
  wire tmp3454;
  wire tmp3455;
  wire tmp3456;
  wire tmp3457;
  wire tmp3458;
  wire tmp3459;
  wire tmp3460;
  wire tmp3461;
  wire tmp3462;
  wire tmp3463;
  wire tmp3464;
  wire tmp3465;
  wire tmp3466;
  wire tmp3467;
  wire tmp3468;
  wire tmp3469;
  wire tmp3470;
  wire tmp3471;
  wire tmp3472;
  wire tmp3473;
  wire tmp3474;
  wire tmp3475;
  wire tmp3476;
  wire tmp3477;
  wire tmp3478;
  wire tmp3479;
  wire tmp3480;
  wire tmp3481;
  wire tmp3482;
  wire tmp3483;
  wire tmp3484;
  wire tmp3485;
  wire tmp3486;
  wire tmp3487;
  wire tmp3488;
  wire tmp3489;
  wire tmp3490;
  wire tmp3491;
  wire tmp3492;
  wire tmp3493;
  wire tmp3494;
  wire tmp3495;
  wire tmp3496;
  wire tmp3497;
  wire tmp3498;
  wire tmp3499;
  wire tmp3500;
  wire tmp3501;
  wire tmp3502;
  wire tmp3503;
  wire tmp3504;
  wire tmp3505;
  wire tmp3506;
  wire tmp3507;
  wire tmp3508;
  wire tmp3509;
  wire tmp3510;
  wire tmp3511;
  wire tmp3512;
  wire tmp3513;
  wire tmp3514;
  wire tmp3515;
  wire tmp3516;
  wire tmp3517;
  wire tmp3518;
  wire tmp3519;
  wire tmp3520;
  wire tmp3521;
  wire tmp3522;
  wire tmp3523;
  wire tmp3524;
  wire tmp3525;
  wire tmp3526;
  wire tmp3527;
  wire tmp3528;
  wire tmp3529;
  wire tmp3530;
  wire tmp3531;
  wire tmp3532;
  wire tmp3533;
  wire tmp3534;
  wire tmp3535;
  wire tmp3536;
  wire tmp3537;
  wire tmp3538;
  wire tmp3539;
  wire tmp3540;
  wire tmp3541;
  wire tmp3542;
  wire tmp3543;
  wire tmp3544;
  wire tmp3545;
  wire tmp3546;
  wire tmp3547;
  wire tmp3548;
  wire tmp3549;
  wire tmp3550;
  wire tmp3551;
  wire tmp3552;
  wire tmp3553;
  wire tmp3554;
  wire tmp3555;
  wire tmp3556;
  wire tmp3557;
  wire tmp3558;
  wire tmp3559;
  wire tmp3560;
  wire tmp3561;
  wire tmp3562;
  wire tmp3563;
  wire tmp3564;
  wire tmp3565;
  wire tmp3566;
  wire tmp3567;
  wire tmp3568;
  wire tmp3569;
  wire tmp3570;
  wire tmp3571;
  wire tmp3572;
  wire tmp3573;
  wire tmp3574;
  wire tmp3575;
  wire tmp3576;
  wire tmp3577;
  wire tmp3578;
  wire tmp3579;
  wire tmp3580;
  wire tmp3581;
  wire tmp3582;
  wire tmp3583;
  wire tmp3584;
  wire tmp3585;
  wire tmp3586;
  wire tmp3587;
  wire tmp3588;
  wire tmp3589;
  wire tmp3590;
  wire tmp3591;
  wire tmp3592;
  wire tmp3593;
  wire tmp3594;
  wire tmp3595;
  wire tmp3596;
  wire tmp3597;
  wire tmp3598;
  wire tmp3599;
  wire tmp3600;
  wire tmp3601;
  wire tmp3602;
  wire tmp3603;
  wire tmp3604;
  wire tmp3605;
  wire tmp3606;
  wire tmp3607;
  wire tmp3608;
  wire tmp3609;
  wire tmp3610;
  wire tmp3611;
  wire tmp3612;
  wire tmp3613;
  wire tmp3614;
  wire tmp3615;
  wire tmp3616;
  wire tmp3617;
  wire tmp3618;
  wire tmp3619;
  wire tmp3620;
  wire tmp3621;
  wire tmp3622;
  wire tmp3623;
  wire tmp3624;
  wire tmp3625;
  wire tmp3626;
  wire tmp3627;
  wire tmp3628;
  wire tmp3629;
  wire tmp3630;
  wire tmp3631;
  wire tmp3632;
  wire tmp3633;
  wire tmp3634;
  wire tmp3635;
  wire tmp3636;
  wire tmp3637;
  wire tmp3638;
  wire tmp3639;
  wire tmp3640;
  wire tmp3641;
  wire tmp3642;
  wire tmp3643;
  wire tmp3644;
  wire tmp3645;
  wire tmp3646;
  wire tmp3647;
  wire tmp3648;
  wire tmp3649;
  wire tmp3650;
  wire tmp3651;
  wire tmp3652;
  wire tmp3653;
  wire tmp3654;
  wire tmp3655;
  wire tmp3656;
  wire tmp3657;
  wire tmp3658;
  wire tmp3659;
  wire tmp3660;
  wire tmp3661;
  wire tmp3662;
  wire tmp3663;
  wire tmp3664;
  wire tmp3665;
  wire tmp3666;
  wire tmp3667;
  wire tmp3668;
  wire tmp3669;
  wire tmp3670;
  wire tmp3671;
  wire tmp3672;
  wire tmp3673;
  wire tmp3674;
  wire tmp3675;
  wire tmp3676;
  wire tmp3677;
  wire tmp3678;
  wire tmp3679;
  wire tmp3680;
  wire tmp3681;
  wire tmp3682;
  wire tmp3683;
  wire tmp3684;
  wire tmp3685;
  wire tmp3686;
  wire tmp3687;
  wire tmp3688;
  wire tmp3689;
  wire tmp3690;
  wire tmp3691;
  wire tmp3692;
  wire tmp3693;
  wire tmp3694;
  wire tmp3695;
  wire tmp3696;
  wire tmp3697;
  wire tmp3698;
  wire tmp3699;
  wire tmp3700;
  wire tmp3701;
  wire tmp3702;
  wire tmp3703;
  wire tmp3704;
  wire tmp3705;
  wire tmp3706;
  wire tmp3707;
  wire tmp3708;
  wire tmp3709;
  wire tmp3710;
  wire tmp3711;
  wire tmp3712;
  wire tmp3713;
  wire tmp3714;
  wire tmp3715;
  wire tmp3716;
  wire tmp3717;
  wire tmp3718;
  wire tmp3719;
  wire tmp3720;
  wire tmp3721;
  wire tmp3722;
  wire tmp3723;
  wire tmp3724;
  wire tmp3725;
  wire tmp3726;
  wire tmp3727;
  wire tmp3728;
  wire tmp3729;
  wire tmp3730;
  wire tmp3731;
  wire tmp3732;
  wire tmp3733;
  wire tmp3734;
  wire tmp3735;
  wire tmp3736;
  wire tmp3737;
  wire tmp3738;
  wire tmp3739;
  wire tmp3740;
  wire tmp3741;
  wire tmp3742;
  wire tmp3743;
  wire tmp3744;
  wire tmp3745;
  wire tmp3746;
  wire tmp3747;
  wire tmp3748;
  wire tmp3749;
  wire tmp3750;
  wire tmp3751;
  wire tmp3752;
  wire tmp3753;
  wire tmp3754;
  wire tmp3755;
  wire tmp3756;
  wire tmp3757;
  wire tmp3758;
  wire tmp3759;
  wire tmp3760;
  wire tmp3761;
  wire tmp3762;
  wire tmp3763;
  wire tmp3764;
  wire tmp3765;
  wire tmp3766;
  wire tmp3767;
  wire tmp3768;
  wire tmp3769;
  wire tmp3770;
  wire tmp3771;
  wire tmp3772;
  wire tmp3773;
  wire tmp3774;
  wire tmp3775;
  wire tmp3776;
  wire tmp3777;
  wire tmp3778;
  wire tmp3779;
  wire tmp3780;
  wire tmp3781;
  wire tmp3782;
  wire tmp3783;
  wire tmp3784;
  wire tmp3785;
  wire tmp3786;
  wire tmp3787;
  wire tmp3788;
  wire tmp3789;
  wire tmp3790;
  wire tmp3791;
  wire tmp3792;
  wire tmp3793;
  wire tmp3794;
  wire tmp3795;
  wire tmp3796;
  wire tmp3797;
  wire tmp3798;
  wire tmp3799;
  wire tmp3800;
  wire tmp3801;
  wire tmp3802;
  wire tmp3803;
  wire tmp3804;
  wire tmp3805;
  wire tmp3806;
  wire tmp3807;
  wire tmp3808;
  wire tmp3809;
  wire tmp3810;
  wire tmp3811;
  wire tmp3812;
  wire tmp3813;
  wire tmp3814;
  wire tmp3815;
  wire tmp3816;
  wire tmp3817;
  wire tmp3818;
  wire tmp3819;
  wire tmp3820;
  wire tmp3821;
  wire tmp3822;
  wire tmp3823;
  wire tmp3824;
  wire tmp3825;
  wire tmp3826;
  wire tmp3827;
  wire tmp3828;
  wire tmp3829;
  wire tmp3830;
  wire tmp3831;
  wire tmp3832;
  wire tmp3833;
  wire tmp3834;
  wire tmp3835;
  wire tmp3836;
  wire tmp3837;
  wire tmp3838;
  wire tmp3839;
  wire tmp3840;
  wire tmp3841;
  wire tmp3842;
  wire tmp3843;
  wire tmp3844;
  wire tmp3845;
  wire tmp3846;
  wire tmp3847;
  wire tmp3848;
  wire tmp3849;
  wire tmp3850;
  wire tmp3851;
  wire tmp3852;
  wire tmp3853;
  wire tmp3854;
  wire tmp3855;
  wire tmp3856;
  wire tmp3857;
  wire tmp3858;
  wire tmp3859;
  wire tmp3860;
  wire tmp3861;
  wire tmp3862;
  wire tmp3863;
  wire tmp3864;
  wire tmp3865;
  wire tmp3866;
  wire tmp3867;
  wire tmp3868;
  wire tmp3869;
  wire tmp3870;
  wire tmp3871;
  wire tmp3872;
  wire tmp3873;
  wire tmp3874;
  wire tmp3875;
  wire tmp3876;
  wire tmp3877;
  wire tmp3878;
  wire tmp3879;
  wire tmp3880;
  wire tmp3881;
  wire tmp3882;
  wire tmp3883;
  wire tmp3884;
  wire tmp3885;
  wire tmp3886;
  wire tmp3887;
  wire tmp3888;
  wire tmp3889;
  wire tmp3890;
  wire tmp3891;
  wire tmp3892;
  wire tmp3893;
  wire tmp3894;
  wire tmp3895;
  wire tmp3896;
  wire tmp3897;
  wire tmp3898;
  wire tmp3899;
  wire tmp3900;
  wire tmp3901;
  wire tmp3902;
  wire tmp3903;
  wire tmp3904;
  wire tmp3905;
  wire tmp3906;
  wire tmp3907;
  wire tmp3908;
  wire tmp3909;
  wire tmp3910;
  wire tmp3911;
  wire tmp3912;
  wire tmp3913;
  wire tmp3914;
  wire tmp3915;
  wire tmp3916;
  wire tmp3917;
  wire tmp3918;
  wire tmp3919;
  wire tmp3920;
  wire tmp3921;
  wire tmp3922;
  wire tmp3923;
  wire tmp3924;
  wire tmp3925;
  wire tmp3926;
  wire tmp3927;
  wire tmp3928;
  wire tmp3929;
  wire tmp3930;
  wire tmp3931;
  wire tmp3932;
  wire tmp3933;
  wire tmp3934;
  wire tmp3935;
  wire tmp3936;
  wire tmp3937;
  wire tmp3938;
  wire tmp3939;
  wire tmp3940;
  wire tmp3941;
  wire tmp3942;
  wire tmp3943;
  wire tmp3944;
  wire tmp3945;
  wire tmp3946;
  wire tmp3947;
  wire tmp3948;
  wire tmp3949;
  wire tmp3950;
  wire tmp3951;
  wire tmp3952;
  wire tmp3953;
  wire tmp3954;
  wire tmp3955;
  wire tmp3956;
  wire tmp3957;
  wire tmp3958;
  wire tmp3959;
  wire tmp3960;
  wire tmp3961;
  wire tmp3962;
  wire tmp3963;
  wire tmp3964;
  wire tmp3965;
  wire tmp3966;
  wire tmp3967;
  wire tmp3968;
  wire tmp3969;
  wire tmp3970;
  wire tmp3971;
  wire tmp3972;
  wire tmp3973;
  wire tmp3974;
  wire tmp3975;
  wire tmp3976;
  wire tmp3977;
  wire tmp3978;
  wire tmp3979;
  wire tmp3980;
  wire tmp3981;
  wire tmp3982;
  wire tmp3983;
  wire tmp3984;
  wire tmp3985;
  wire tmp3986;
  wire tmp3987;
  wire tmp3988;
  wire tmp3989;
  wire tmp3990;
  wire tmp3991;
  wire tmp3992;
  wire tmp3993;
  wire tmp3994;
  wire tmp3995;
  wire tmp3996;
  wire tmp3997;
  wire tmp3998;
  wire tmp3999;
  wire tmp4000;
  wire tmp4001;
  wire tmp4002;
  wire tmp4003;
  wire tmp4004;
  wire tmp4005;
  wire tmp4006;
  wire tmp4007;
  wire tmp4008;
  wire tmp4009;
  wire tmp4010;
  wire tmp4011;
  wire tmp4012;
  wire tmp4013;
  wire tmp4014;
  wire tmp4015;
  wire tmp4016;
  wire tmp4017;
  wire tmp4018;
  wire tmp4019;
  wire tmp4020;
  wire tmp4021;
  wire tmp4022;
  wire tmp4023;
  wire tmp4024;
  wire tmp4025;
  wire tmp4026;
  wire tmp4027;
  wire tmp4028;
  wire tmp4029;
  wire tmp4030;
  wire tmp4031;
  wire tmp4032;
  wire tmp4033;
  wire tmp4034;
  wire tmp4035;
  wire tmp4036;
  wire tmp4037;
  wire tmp4038;
  wire tmp4039;
  wire tmp4040;
  wire tmp4041;
  wire tmp4042;
  wire tmp4043;
  wire tmp4044;
  wire tmp4045;
  wire tmp4046;
  wire tmp4047;
  wire tmp4048;
  wire tmp4049;
  wire tmp4050;
  wire tmp4051;
  wire tmp4052;
  wire tmp4053;
  wire tmp4054;
  wire tmp4055;
  wire tmp4056;
  wire tmp4057;
  wire tmp4058;
  wire tmp4059;
  wire tmp4060;
  wire tmp4061;
  wire tmp4062;
  wire tmp4063;
  wire tmp4064;
  wire tmp4065;
  wire tmp4066;
  wire tmp4067;
  wire tmp4068;
  wire tmp4069;
  wire tmp4070;
  wire tmp4071;
  wire tmp4072;
  wire tmp4073;
  wire tmp4074;
  wire tmp4075;
  wire tmp4076;
  wire tmp4077;
  wire tmp4078;
  wire tmp4079;
  wire tmp4080;
  wire tmp4081;
  wire tmp4082;
  wire tmp4083;
  wire tmp4084;
  wire tmp4085;
  wire tmp4086;
  wire tmp4087;
  wire tmp4088;
  wire tmp4089;
  wire tmp4090;
  wire tmp4091;
  wire tmp4092;
  wire tmp4093;
  wire tmp4094;
  wire tmp4095;
  wire tmp4096;
  wire tmp4097;
  wire tmp4098;
  wire tmp4099;
  wire tmp4100;
  wire tmp4101;
  wire tmp4102;
  wire tmp4103;
  wire tmp4104;
  wire tmp4105;
  wire tmp4106;
  wire tmp4107;
  wire tmp4108;
  wire tmp4109;
  wire tmp4110;
  wire tmp4111;
  wire tmp4112;
  wire tmp4113;
  wire tmp4114;
  wire tmp4115;
  wire tmp4116;
  wire tmp4117;
  wire tmp4118;
  wire tmp4119;
  wire tmp4120;
  wire tmp4121;
  wire tmp4122;
  wire tmp4123;
  wire tmp4124;
  wire tmp4125;
  wire tmp4126;
  wire tmp4127;
  wire tmp4128;
  wire tmp4129;
  wire tmp4130;
  wire tmp4131;
  wire tmp4132;
  wire tmp4133;
  wire tmp4134;
  wire tmp4135;
  wire tmp4136;
  wire tmp4137;
  wire tmp4138;
  wire tmp4139;
  wire tmp4140;
  wire tmp4141;
  wire tmp4142;
  wire tmp4143;
  wire tmp4144;
  wire tmp4145;
  wire tmp4146;
  wire tmp4147;
  wire tmp4148;
  wire tmp4149;
  wire tmp4150;
  wire tmp4151;
  wire tmp4152;
  wire tmp4153;
  wire tmp4154;
  wire tmp4155;
  wire tmp4156;
  wire tmp4157;
  wire tmp4158;
  wire tmp4159;
  wire tmp4160;
  wire tmp4161;
  wire tmp4162;
  wire tmp4163;
  wire tmp4164;
  wire tmp4165;
  wire tmp4166;
  wire tmp4167;
  wire tmp4168;
  wire tmp4169;
  wire tmp4170;
  wire tmp4171;
  wire tmp4172;
  wire tmp4173;
  wire tmp4174;
  wire tmp4175;
  wire tmp4176;
  wire tmp4177;
  wire tmp4178;
  wire tmp4179;
  wire tmp4180;
  wire tmp4181;
  wire tmp4182;
  wire tmp4183;
  wire tmp4184;
  wire tmp4185;
  wire tmp4186;
  wire tmp4187;
  wire tmp4188;
  wire tmp4189;
  wire tmp4190;
  wire tmp4191;
  wire tmp4192;
  wire tmp4193;
  wire tmp4194;
  wire tmp4195;
  wire tmp4196;
  wire tmp4197;
  wire tmp4198;
  wire tmp4199;
  wire tmp4200;
  wire tmp4201;
  wire tmp4202;
  wire tmp4203;
  wire tmp4204;
  wire tmp4205;
  wire tmp4206;
  wire tmp4207;
  wire tmp4208;
  wire tmp4209;
  wire tmp4210;
  wire tmp4211;
  wire tmp4212;
  wire tmp4213;
  wire tmp4214;
  wire tmp4215;
  wire tmp4216;
  wire tmp4217;
  wire tmp4218;
  wire tmp4219;
  wire tmp4220;
  wire tmp4221;
  wire tmp4222;
  wire tmp4223;
  wire tmp4224;
  wire tmp4225;
  wire tmp4226;
  wire tmp4227;
  wire tmp4228;
  wire tmp4229;
  wire tmp4230;
  wire tmp4231;
  wire tmp4232;
  wire tmp4233;
  wire tmp4234;
  wire tmp4235;
  wire tmp4236;
  wire tmp4237;
  wire tmp4238;
  wire tmp4239;
  wire tmp4240;
  wire tmp4241;
  wire tmp4242;
  wire tmp4243;
  wire tmp4244;
  wire tmp4245;
  wire tmp4246;
  wire tmp4247;
  wire tmp4248;
  wire tmp4249;
  wire tmp4250;
  wire tmp4251;
  wire tmp4252;
  wire tmp4253;
  wire tmp4254;
  wire tmp4255;
  wire tmp4256;
  wire tmp4257;
  wire tmp4258;
  wire tmp4259;
  wire tmp4260;
  wire tmp4261;
  wire tmp4262;
  wire tmp4263;
  wire tmp4264;
  wire tmp4265;
  wire tmp4266;
  wire tmp4267;
  wire tmp4268;
  wire tmp4269;
  wire tmp4270;
  wire tmp4271;
  wire tmp4272;
  wire tmp4273;
  wire tmp4274;
  wire tmp4275;
  wire tmp4276;
  wire tmp4277;
  wire tmp4278;
  wire tmp4279;
  wire tmp4280;
  wire tmp4281;
  wire tmp4282;
  wire tmp4283;
  wire tmp4284;
  wire tmp4285;
  wire tmp4286;
  wire tmp4287;
  wire tmp4288;
  wire tmp4289;
  wire tmp4290;
  wire tmp4291;
  wire tmp4292;
  wire tmp4293;
  wire tmp4294;
  wire tmp4295;
  wire tmp4296;
  wire tmp4297;
  wire tmp4298;
  wire tmp4299;
  wire tmp4300;
  wire tmp4301;
  wire tmp4302;
  wire tmp4303;
  wire tmp4304;
  wire tmp4305;
  wire tmp4306;
  wire tmp4307;
  wire tmp4308;
  wire tmp4309;
  wire tmp4310;
  wire tmp4311;
  wire tmp4312;
  wire tmp4313;
  wire tmp4314;
  wire tmp4315;
  wire tmp4316;
  wire tmp4317;
  wire tmp4318;
  wire tmp4319;
  wire tmp4320;
  wire tmp4321;
  wire tmp4322;
  wire tmp4323;
  wire tmp4324;
  wire tmp4325;
  wire tmp4326;
  wire tmp4327;
  wire tmp4328;
  wire tmp4329;
  wire tmp4330;
  wire tmp4331;
  wire tmp4332;
  wire tmp4333;
  wire tmp4334;
  wire tmp4335;
  wire tmp4336;
  wire tmp4337;
  wire tmp4338;
  wire tmp4339;
  wire tmp4340;
  wire tmp4341;
  wire tmp4342;
  wire tmp4343;
  wire tmp4344;
  wire tmp4345;
  wire tmp4346;
  wire tmp4347;
  wire tmp4348;
  wire tmp4349;
  wire tmp4350;
  wire tmp4351;
  wire tmp4352;
  wire tmp4353;
  wire tmp4354;
  wire tmp4355;
  wire tmp4356;
  wire tmp4357;
  wire tmp4358;
  wire tmp4359;
  wire tmp4360;
  wire tmp4361;
  wire tmp4362;
  wire tmp4363;
  wire tmp4364;
  wire tmp4365;
  wire tmp4366;
  wire tmp4367;
  wire tmp4368;
  wire tmp4369;
  wire tmp4370;
  wire tmp4371;
  wire tmp4372;
  wire tmp4373;
  wire tmp4374;
  wire tmp4375;
  wire tmp4376;
  wire tmp4377;
  wire tmp4378;
  wire tmp4379;
  wire tmp4380;
  wire tmp4381;
  wire tmp4382;
  wire tmp4383;
  wire tmp4384;
  wire tmp4385;
  wire tmp4386;
  wire tmp4387;
  wire tmp4388;
  wire tmp4389;
  wire tmp4390;
  wire tmp4391;
  wire tmp4392;
  wire tmp4393;
  wire tmp4394;
  wire tmp4395;
  wire tmp4396;
  wire tmp4397;
  wire tmp4398;
  wire tmp4399;
  wire tmp4400;
  wire tmp4401;
  wire tmp4402;
  wire tmp4403;
  wire tmp4404;
  wire tmp4405;
  wire tmp4406;
  wire tmp4407;
  wire tmp4408;
  wire tmp4409;
  wire tmp4410;
  wire tmp4411;
  wire tmp4412;
  wire tmp4413;
  wire tmp4414;
  wire tmp4415;
  wire tmp4416;
  wire tmp4417;
  wire tmp4418;
  wire tmp4419;
  wire tmp4420;
  wire tmp4421;
  wire tmp4422;
  wire tmp4423;
  wire tmp4424;
  wire tmp4425;
  wire tmp4426;
  wire tmp4427;
  wire tmp4428;
  wire tmp4429;
  wire tmp4430;
  wire tmp4431;
  wire tmp4432;
  wire tmp4433;
  wire tmp4434;
  wire tmp4435;
  wire tmp4436;
  wire tmp4437;
  wire tmp4438;
  wire tmp4439;
  wire tmp4440;
  wire tmp4441;
  wire tmp4442;
  wire tmp4443;
  wire tmp4444;
  wire tmp4445;
  wire tmp4446;
  wire tmp4447;
  wire tmp4448;
  wire tmp4449;
  wire tmp4450;
  wire tmp4451;
  wire tmp4452;
  wire tmp4453;
  wire tmp4454;
  wire tmp4455;
  wire tmp4456;
  wire tmp4457;
  wire tmp4458;
  wire tmp4459;
  wire tmp4460;
  wire tmp4461;
  wire tmp4462;
  wire tmp4463;
  wire tmp4464;
  wire tmp4465;
  wire tmp4466;
  wire tmp4467;
  wire tmp4468;
  wire tmp4469;
  wire tmp4470;
  wire tmp4471;
  wire tmp4472;
  wire tmp4473;
  wire tmp4474;
  wire tmp4475;
  wire tmp4476;
  wire tmp4477;
  wire tmp4478;
  wire tmp4479;
  wire tmp4480;
  wire tmp4481;
  wire tmp4482;
  wire tmp4483;
  wire tmp4484;
  wire tmp4485;
  wire tmp4486;
  wire tmp4487;
  wire tmp4488;
  wire tmp4489;
  wire tmp4490;
  wire tmp4491;
  wire tmp4492;
  wire tmp4493;
  wire tmp4494;
  wire tmp4495;
  wire tmp4496;
  wire tmp4497;
  wire tmp4498;
  wire tmp4499;
  wire tmp4500;
  wire tmp4501;
  wire tmp4502;
  wire tmp4503;
  wire tmp4504;
  wire tmp4505;
  wire tmp4506;
  wire tmp4507;
  wire tmp4508;
  wire tmp4509;
  wire tmp4510;
  wire tmp4511;
  wire tmp4512;
  wire tmp4513;
  wire tmp4514;
  wire tmp4515;
  wire tmp4516;
  wire tmp4517;
  wire tmp4518;
  wire tmp4519;
  wire tmp4520;
  wire tmp4521;
  wire tmp4522;
  wire tmp4523;
  wire tmp4524;
  wire tmp4525;
  wire tmp4526;
  wire tmp4527;
  wire tmp4528;
  wire tmp4529;
  wire tmp4530;
  wire tmp4531;
  wire tmp4532;
  wire tmp4533;
  wire tmp4534;
  wire tmp4535;
  wire tmp4536;
  wire tmp4537;
  wire tmp4538;
  wire tmp4539;
  wire tmp4540;
  wire tmp4541;
  wire tmp4542;
  wire tmp4543;
  wire tmp4544;
  wire tmp4545;
  wire tmp4546;
  wire tmp4547;
  wire tmp4548;
  wire tmp4549;
  wire tmp4550;
  wire tmp4551;
  wire tmp4552;
  wire tmp4553;
  wire tmp4554;
  wire tmp4555;
  wire tmp4556;
  wire tmp4557;
  wire tmp4558;
  wire tmp4559;
  wire tmp4560;
  wire tmp4561;
  wire tmp4562;
  wire tmp4563;
  wire tmp4564;
  wire tmp4565;
  wire tmp4566;
  wire tmp4567;
  wire tmp4568;
  wire tmp4569;
  wire tmp4570;
  wire tmp4571;
  wire tmp4572;
  wire tmp4573;
  wire tmp4574;
  wire tmp4575;
  wire tmp4576;
  wire tmp4577;
  wire tmp4578;
  wire tmp4579;
  wire tmp4580;
  wire tmp4581;
  wire tmp4582;
  wire tmp4583;
  wire tmp4584;
  wire tmp4585;
  wire tmp4586;
  wire tmp4587;
  wire tmp4588;
  wire tmp4589;
  wire tmp4590;
  wire tmp4591;
  wire tmp4592;
  wire tmp4593;
  wire tmp4594;
  wire tmp4595;
  wire tmp4596;
  wire tmp4597;
  wire tmp4598;
  wire tmp4599;
  wire tmp4600;
  wire tmp4601;
  wire tmp4602;
  wire tmp4603;
  wire tmp4604;
  wire tmp4605;
  wire tmp4606;
  wire tmp4607;
  wire tmp4608;
  wire tmp4609;
  wire tmp4610;
  wire tmp4611;
  wire tmp4612;
  wire tmp4613;
  wire tmp4614;
  wire tmp4615;
  wire tmp4616;
  wire tmp4617;
  wire tmp4618;
  wire tmp4619;
  wire tmp4620;
  wire tmp4621;
  wire tmp4622;
  wire tmp4623;
  wire tmp4624;
  wire tmp4625;
  wire tmp4626;
  wire tmp4627;
  wire tmp4628;
  wire tmp4629;
  wire tmp4630;
  wire tmp4631;
  wire tmp4632;
  wire tmp4633;
  wire tmp4634;
  wire tmp4635;
  wire tmp4636;
  wire tmp4637;
  wire tmp4638;
  wire tmp4639;
  wire tmp4640;
  wire tmp4641;
  wire tmp4642;
  wire tmp4643;
  wire tmp4644;
  wire tmp4645;
  wire tmp4646;
  wire tmp4647;
  wire tmp4648;
  wire tmp4649;
  wire tmp4650;
  wire tmp4651;
  wire tmp4652;
  wire tmp4653;
  wire tmp4654;
  wire tmp4655;
  wire tmp4656;
  wire tmp4657;
  wire tmp4658;
  wire tmp4659;
  wire tmp4660;
  wire tmp4661;
  wire tmp4662;
  wire tmp4663;
  wire tmp4664;
  wire tmp4665;
  wire tmp4666;
  wire tmp4667;
  wire tmp4668;
  wire tmp4669;
  wire tmp4670;
  wire tmp4671;
  wire tmp4672;
  wire tmp4673;
  wire tmp4674;
  wire tmp4675;
  wire tmp4676;
  wire tmp4677;
  wire tmp4678;
  wire tmp4679;
  wire tmp4680;
  wire tmp4681;
  wire tmp4682;
  wire tmp4683;
  wire tmp4684;
  wire tmp4685;
  wire tmp4686;
  wire tmp4687;
  wire tmp4688;
  wire tmp4689;
  wire tmp4690;
  wire tmp4691;
  wire tmp4692;
  wire tmp4693;
  wire tmp4694;
  wire tmp4695;
  wire tmp4696;
  wire tmp4697;
  wire tmp4698;
  wire tmp4699;
  wire tmp4700;
  wire tmp4701;
  wire tmp4702;
  wire tmp4703;
  wire tmp4704;
  wire tmp4705;
  wire tmp4706;
  wire tmp4707;
  wire tmp4708;
  wire tmp4709;
  wire tmp4710;
  wire tmp4711;
  wire tmp4712;
  wire tmp4713;
  wire tmp4714;
  wire tmp4715;
  wire tmp4716;
  wire tmp4717;
  wire tmp4718;
  wire tmp4719;
  wire tmp4720;
  wire tmp4721;
  wire tmp4722;
  wire tmp4723;
  wire tmp4724;
  wire tmp4725;
  wire tmp4726;
  wire tmp4727;
  wire tmp4728;
  wire tmp4729;
  wire tmp4730;
  wire tmp4731;
  wire tmp4732;
  wire tmp4733;
  wire tmp4734;
  wire tmp4735;
  wire tmp4736;
  wire tmp4737;
  wire tmp4738;
  wire tmp4739;
  wire tmp4740;
  wire tmp4741;
  wire tmp4742;
  wire tmp4743;
  wire tmp4744;
  wire tmp4745;
  wire tmp4746;
  wire tmp4747;
  wire tmp4748;
  wire tmp4749;
  wire tmp4750;
  wire tmp4751;
  wire tmp4752;
  wire tmp4753;
  wire tmp4754;
  wire tmp4755;
  wire tmp4756;
  wire tmp4757;
  wire tmp4758;
  wire tmp4759;
  wire tmp4760;
  wire tmp4761;
  wire tmp4762;
  wire tmp4763;
  wire tmp4764;
  wire tmp4765;
  wire tmp4766;
  wire tmp4767;
  wire tmp4768;
  wire tmp4769;
  wire tmp4770;
  wire tmp4771;
  wire tmp4772;
  wire tmp4773;
  wire tmp4774;
  wire tmp4775;
  wire tmp4776;
  wire tmp4777;
  wire tmp4778;
  wire tmp4779;
  wire tmp4780;
  wire tmp4781;
  wire tmp4782;
  wire tmp4783;
  wire tmp4784;
  wire tmp4785;
  wire tmp4786;
  wire tmp4787;
  wire tmp4788;
  wire tmp4789;
  wire tmp4790;
  wire tmp4791;
  wire tmp4792;
  wire tmp4793;
  wire tmp4794;
  wire tmp4795;
  wire tmp4796;
  wire tmp4797;
  wire tmp4798;
  wire tmp4799;
  wire tmp4800;
  wire tmp4801;
  wire tmp4802;
  wire tmp4803;
  wire tmp4804;
  wire tmp4805;
  wire tmp4806;
  wire tmp4807;
  wire tmp4808;
  wire tmp4809;
  wire tmp4810;
  wire tmp4811;
  wire tmp4812;
  wire tmp4813;
  wire tmp4814;
  wire tmp4815;
  wire tmp4816;
  wire tmp4817;
  wire tmp4818;
  wire tmp4819;
  wire tmp4820;
  wire tmp4821;
  wire tmp4822;
  wire tmp4823;
  wire tmp4824;
  wire tmp4825;
  wire tmp4826;
  wire tmp4827;
  wire tmp4828;
  wire tmp4829;
  wire tmp4830;
  wire tmp4831;
  wire tmp4832;
  wire tmp4833;
  wire tmp4834;
  wire tmp4835;
  wire tmp4836;
  wire tmp4837;
  wire tmp4838;
  wire tmp4839;
  wire tmp4840;
  wire tmp4841;
  wire tmp4842;
  wire tmp4843;
  wire tmp4844;
  wire tmp4845;
  wire tmp4846;
  wire tmp4847;
  wire tmp4848;
  wire tmp4849;
  wire tmp4850;
  wire tmp4851;
  wire tmp4852;
  wire tmp4853;
  wire tmp4854;
  wire tmp4855;
  wire tmp4856;
  wire tmp4857;
  wire tmp4858;
  wire tmp4859;
  wire tmp4860;
  wire tmp4861;
  wire tmp4862;
  wire tmp4863;
  wire tmp4864;
  wire tmp4865;
  wire tmp4866;
  wire tmp4867;
  wire tmp4868;
  wire tmp4869;
  wire tmp4870;
  wire tmp4871;
  wire tmp4872;
  wire tmp4873;
  wire tmp4874;
  wire tmp4875;
  wire tmp4876;
  wire tmp4877;
  wire tmp4878;
  wire tmp4879;
  wire tmp4880;
  wire tmp4881;
  wire tmp4882;
  wire tmp4883;
  wire tmp4884;
  wire tmp4885;
  wire tmp4886;
  wire tmp4887;
  wire tmp4888;
  wire tmp4889;
  wire tmp4890;
  wire tmp4891;
  wire tmp4892;
  wire tmp4893;
  wire tmp4894;
  wire tmp4895;
  wire tmp4896;
  wire tmp4897;
  wire tmp4898;
  wire tmp4899;
  wire tmp4900;
  wire tmp4901;
  wire tmp4902;
  wire tmp4903;
  wire tmp4904;
  wire tmp4905;
  wire tmp4906;
  wire tmp4907;
  wire tmp4908;
  wire tmp4909;
  wire tmp4910;
  wire tmp4911;
  wire tmp4912;
  wire tmp4913;
  wire tmp4914;
  wire tmp4915;
  wire tmp4916;
  wire tmp4917;
  wire tmp4918;
  wire tmp4919;
  wire tmp4920;
  wire tmp4921;
  wire tmp4922;
  wire tmp4923;
  wire tmp4924;
  wire tmp4925;
  wire tmp4926;
  wire tmp4927;
  wire tmp4928;
  wire tmp4929;
  wire tmp4930;
  wire tmp4931;
  wire tmp4932;
  wire tmp4933;
  wire tmp4934;
  wire tmp4935;
  wire tmp4936;
  wire tmp4937;
  wire tmp4938;
  wire tmp4939;
  wire tmp4940;
  wire tmp4941;
  wire tmp4942;
  wire tmp4943;
  wire tmp4944;
  wire tmp4945;
  wire tmp4946;
  wire tmp4947;
  wire tmp4948;
  wire tmp4949;
  wire tmp4950;
  wire tmp4951;
  wire tmp4952;
  wire tmp4953;
  wire tmp4954;
  wire tmp4955;
  wire tmp4956;
  wire tmp4957;
  wire tmp4958;
  wire tmp4959;
  wire tmp4960;
  wire tmp4961;
  wire tmp4962;
  wire tmp4963;
  wire tmp4964;
  wire tmp4965;
  wire tmp4966;
  wire tmp4967;
  wire tmp4968;
  wire tmp4969;
  wire tmp4970;
  wire tmp4971;
  wire tmp4972;
  wire tmp4973;
  wire tmp4974;
  wire tmp4975;
  wire tmp4976;
  wire tmp4977;
  wire tmp4978;
  wire tmp4979;
  wire tmp4980;
  wire tmp4981;
  wire tmp4982;
  wire tmp4983;
  wire tmp4984;
  wire tmp4985;
  wire tmp4986;
  wire tmp4987;
  wire tmp4988;
  wire tmp4989;
  wire tmp4990;
  wire tmp4991;
  wire tmp4992;
  wire tmp4993;
  wire tmp4994;
  wire tmp4995;
  wire tmp4996;
  wire tmp4997;
  wire tmp4998;
  wire tmp4999;
  wire tmp5000;
  wire tmp5001;
  wire tmp5002;
  wire tmp5003;
  wire tmp5004;
  wire tmp5005;
  wire tmp5006;
  wire tmp5007;
  wire tmp5008;
  wire tmp5009;
  wire tmp5010;
  wire tmp5011;
  wire tmp5012;
  wire tmp5013;
  wire tmp5014;
  wire tmp5015;
  wire tmp5016;
  wire tmp5017;
  wire tmp5018;
  wire tmp5019;
  wire tmp5020;
  wire tmp5021;
  wire tmp5022;
  wire tmp5023;
  wire tmp5024;
  wire tmp5025;
  wire tmp5026;
  wire tmp5027;
  wire tmp5028;
  wire tmp5029;
  wire tmp5030;
  wire tmp5031;
  wire tmp5032;
  wire tmp5033;
  wire tmp5034;
  wire tmp5035;
  wire tmp5036;
  wire tmp5037;
  wire tmp5038;
  wire tmp5039;
  wire tmp5040;
  wire tmp5041;
  wire tmp5042;
  wire tmp5043;
  wire tmp5044;
  wire tmp5045;
  wire tmp5046;
  wire tmp5047;
  wire tmp5048;
  wire tmp5049;
  wire tmp5050;
  wire tmp5051;
  wire tmp5052;
  wire tmp5053;
  wire tmp5054;
  wire tmp5055;
  wire tmp5056;
  wire tmp5057;
  wire tmp5058;
  wire tmp5059;
  wire tmp5060;
  wire tmp5061;
  wire tmp5062;
  wire tmp5063;
  wire tmp5064;
  wire tmp5065;
  wire tmp5066;
  wire tmp5067;
  wire tmp5068;
  wire tmp5069;
  wire tmp5070;
  wire tmp5071;
  wire tmp5072;
  wire tmp5073;
  wire tmp5074;
  wire tmp5075;
  wire tmp5076;
  wire tmp5077;
  wire tmp5078;
  wire tmp5079;
  wire tmp5080;
  wire tmp5081;
  wire tmp5082;
  wire tmp5083;
  wire tmp5084;
  wire tmp5085;
  wire tmp5086;
  wire tmp5087;
  wire tmp5088;
  wire tmp5089;
  wire tmp5090;
  wire tmp5091;
  wire tmp5092;
  wire tmp5093;
  wire tmp5094;
  wire tmp5095;
  wire tmp5096;
  wire tmp5097;
  wire tmp5098;
  wire tmp5099;
  wire tmp5100;
  wire tmp5101;
  wire tmp5102;
  wire tmp5103;
  wire tmp5104;
  wire tmp5105;
  wire tmp5106;
  wire tmp5107;
  wire tmp5108;
  wire tmp5109;
  wire tmp5110;
  wire tmp5111;
  wire tmp5112;
  wire tmp5113;
  wire tmp5114;
  wire tmp5115;
  wire tmp5116;
  wire tmp5117;
  wire tmp5118;
  wire tmp5119;
  wire tmp5120;
  wire tmp5121;
  wire tmp5122;
  wire tmp5123;
  wire tmp5124;
  wire tmp5125;
  wire tmp5126;
  wire tmp5127;
  wire tmp5128;
  wire tmp5129;
  wire tmp5130;
  wire tmp5131;
  wire tmp5132;
  wire tmp5133;
  wire tmp5134;
  wire tmp5135;
  wire tmp5136;
  wire tmp5137;
  wire tmp5138;
  wire tmp5139;
  wire tmp5140;
  wire tmp5141;
  wire tmp5142;
  wire tmp5143;
  wire tmp5144;
  wire tmp5145;
  wire tmp5146;
  wire tmp5147;
  wire tmp5148;
  wire tmp5149;
  wire tmp5150;
  wire tmp5151;
  wire tmp5152;
  wire tmp5153;
  wire tmp5154;
  wire tmp5155;
  wire tmp5156;
  wire tmp5157;
  wire tmp5158;
  wire tmp5159;
  wire tmp5160;
  wire tmp5161;
  wire tmp5162;
  wire tmp5163;
  wire tmp5164;
  wire tmp5165;
  wire tmp5166;
  wire tmp5167;
  wire tmp5168;
  wire tmp5169;
  wire tmp5170;
  wire tmp5171;
  wire tmp5172;
  wire tmp5173;
  wire tmp5174;
  wire tmp5175;
  wire tmp5176;
  wire tmp5177;
  wire tmp5178;
  wire tmp5179;
  wire tmp5180;
  wire tmp5181;
  wire tmp5182;
  wire tmp5183;
  wire tmp5184;
  wire tmp5185;
  wire tmp5186;
  wire tmp5187;
  wire tmp5188;
  wire tmp5189;
  wire tmp5190;
  wire tmp5191;
  wire tmp5192;
  wire tmp5193;
  wire tmp5194;
  wire tmp5195;
  wire tmp5196;
  wire tmp5197;
  wire tmp5198;
  wire tmp5199;
  wire tmp5200;
  wire tmp5201;
  wire tmp5202;
  wire tmp5203;
  wire tmp5204;
  wire tmp5205;
  wire tmp5206;
  wire tmp5207;
  wire tmp5208;
  wire tmp5209;
  wire tmp5210;
  wire tmp5211;
  wire tmp5212;
  wire tmp5213;
  wire tmp5214;
  wire tmp5215;
  wire tmp5216;
  wire tmp5217;
  wire tmp5218;
  wire tmp5219;
  wire tmp5220;
  wire tmp5221;
  wire tmp5222;
  wire tmp5223;
  wire tmp5224;
  wire tmp5225;
  wire tmp5226;
  wire tmp5227;
  wire tmp5228;
  wire tmp5229;
  wire tmp5230;
  wire tmp5231;
  wire tmp5232;
  wire tmp5233;
  wire tmp5234;
  wire tmp5235;
  wire tmp5236;
  wire tmp5237;
  wire tmp5238;
  wire tmp5239;
  wire tmp5240;
  wire tmp5241;
  wire tmp5242;
  wire tmp5243;
  wire tmp5244;
  wire tmp5245;
  wire tmp5246;
  wire tmp5247;
  wire tmp5248;
  wire tmp5249;
  wire tmp5250;
  wire tmp5251;
  wire tmp5252;
  wire tmp5253;
  wire tmp5254;
  wire tmp5255;
  wire tmp5256;
  wire tmp5257;
  wire tmp5258;
  wire tmp5259;
  wire tmp5260;
  wire tmp5261;
  wire tmp5262;
  wire tmp5263;
  wire tmp5264;
  wire tmp5265;
  wire tmp5266;
  wire tmp5267;
  wire tmp5268;
  wire tmp5269;
  wire tmp5270;
  wire tmp5271;
  wire tmp5272;
  wire tmp5273;
  wire tmp5274;
  wire tmp5275;
  wire tmp5276;
  wire tmp5277;
  wire tmp5278;
  wire tmp5279;
  wire tmp5280;
  wire tmp5281;
  wire tmp5282;
  wire tmp5283;
  wire tmp5284;
  wire tmp5285;
  wire tmp5286;
  wire tmp5287;
  wire tmp5288;
  wire tmp5289;
  wire tmp5290;
  wire tmp5291;
  wire tmp5292;
  wire tmp5293;
  wire tmp5294;
  wire tmp5295;
  wire tmp5296;
  wire tmp5297;
  wire tmp5298;
  wire tmp5299;
  wire tmp5300;
  wire tmp5301;
  wire tmp5302;
  wire tmp5303;
  wire tmp5304;
  wire tmp5305;
  wire tmp5306;
  wire tmp5307;
  wire tmp5308;
  wire tmp5309;
  wire tmp5310;
  wire tmp5311;
  wire tmp5312;
  wire tmp5313;
  wire tmp5314;
  wire tmp5315;
  wire tmp5316;
  wire tmp5317;
  wire tmp5318;
  wire tmp5319;
  wire tmp5320;
  wire tmp5321;
  wire tmp5322;
  wire tmp5323;
  wire tmp5324;
  wire tmp5325;
  wire tmp5326;
  wire tmp5327;
  wire tmp5328;
  wire tmp5329;
  wire tmp5330;
  wire tmp5331;
  wire tmp5332;
  wire tmp5333;
  wire tmp5334;
  wire tmp5335;
  wire tmp5336;
  wire tmp5337;
  wire tmp5338;
  wire tmp5339;
  wire tmp5340;
  wire tmp5341;
  wire tmp5342;
  wire tmp5343;
  wire tmp5344;
  wire tmp5345;
  wire tmp5346;
  wire tmp5347;
  wire tmp5348;
  wire tmp5349;
  wire tmp5350;
  wire tmp5351;
  wire tmp5352;
  wire tmp5353;
  wire tmp5354;
  wire tmp5355;
  wire tmp5356;
  wire tmp5357;
  wire tmp5358;
  wire tmp5359;
  wire tmp5360;
  wire tmp5361;
  wire tmp5362;
  wire tmp5363;
  wire tmp5364;
  wire tmp5365;
  wire tmp5366;
  wire tmp5367;
  wire tmp5368;
  wire tmp5369;
  wire tmp5370;
  wire tmp5371;
  wire tmp5372;
  wire tmp5373;
  wire tmp5374;
  wire tmp5375;
  wire tmp5376;
  wire tmp5377;
  wire tmp5378;
  wire tmp5379;
  wire tmp5380;
  wire tmp5381;
  wire tmp5382;
  wire tmp5383;
  wire tmp5384;
  wire tmp5385;
  wire tmp5386;
  wire tmp5387;
  wire tmp5388;
  wire tmp5389;
  wire tmp5390;
  wire tmp5391;
  wire tmp5392;
  wire tmp5393;
  wire tmp5394;
  wire tmp5395;
  wire tmp5396;
  wire tmp5397;
  wire tmp5398;
  wire tmp5399;
  wire tmp5400;
  wire tmp5401;
  wire tmp5402;
  wire tmp5403;
  wire tmp5404;
  wire tmp5405;
  wire tmp5406;
  wire tmp5407;
  wire tmp5408;
  wire tmp5409;
  wire tmp5410;
  wire tmp5411;
  wire tmp5412;
  wire tmp5413;
  wire tmp5414;
  wire tmp5415;
  wire tmp5416;
  wire tmp5417;
  wire tmp5418;
  wire tmp5419;
  wire tmp5420;
  wire tmp5421;
  wire tmp5422;
  wire tmp5423;
  wire tmp5424;
  wire tmp5425;
  wire tmp5426;
  wire tmp5427;
  wire tmp5428;
  wire tmp5429;
  wire tmp5430;
  wire tmp5431;
  wire tmp5432;
  wire tmp5433;
  wire tmp5434;
  wire tmp5435;
  wire tmp5436;
  wire tmp5437;
  wire tmp5438;
  wire tmp5439;
  wire tmp5440;
  wire tmp5441;
  wire tmp5442;
  wire tmp5443;
  wire tmp5444;
  wire tmp5445;
  wire tmp5446;
  wire tmp5447;
  wire tmp5448;
  wire tmp5449;
  wire tmp5450;
  wire tmp5451;
  wire tmp5452;
  wire tmp5453;
  wire tmp5454;
  wire tmp5455;
  wire tmp5456;
  wire tmp5457;
  wire tmp5458;
  wire tmp5459;
  wire tmp5460;
  wire tmp5461;
  wire tmp5462;
  wire tmp5463;
  wire tmp5464;
  wire tmp5465;
  wire tmp5466;
  wire tmp5467;
  wire tmp5468;
  wire tmp5469;
  wire tmp5470;
  wire tmp5471;
  wire tmp5472;
  wire tmp5473;
  wire tmp5474;
  wire tmp5475;
  wire tmp5476;
  wire tmp5477;
  wire tmp5478;
  wire tmp5479;
  wire tmp5480;
  wire tmp5481;
  wire tmp5482;
  wire tmp5483;
  wire tmp5484;
  wire tmp5485;
  wire tmp5486;
  wire tmp5487;
  wire tmp5488;
  wire tmp5489;
  wire tmp5490;
  wire tmp5491;
  wire tmp5492;
  wire tmp5493;
  wire tmp5494;
  wire tmp5495;
  wire tmp5496;
  wire tmp5497;
  wire tmp5498;
  wire tmp5499;
  wire tmp5500;
  wire tmp5501;
  wire tmp5502;
  wire tmp5503;
  wire tmp5504;
  wire tmp5505;
  wire tmp5506;
  wire tmp5507;
  wire tmp5508;
  wire tmp5509;
  wire tmp5510;
  wire tmp5511;
  wire tmp5512;
  wire tmp5513;
  wire tmp5514;
  wire tmp5515;
  wire tmp5516;
  wire tmp5517;
  wire tmp5518;
  wire tmp5519;
  wire tmp5520;
  wire tmp5521;
  wire tmp5522;
  wire tmp5523;
  wire tmp5524;
  wire tmp5525;
  wire tmp5526;
  wire tmp5527;
  wire tmp5528;
  wire tmp5529;
  wire tmp5530;
  wire tmp5531;
  wire tmp5532;
  wire tmp5533;
  wire tmp5534;
  wire tmp5535;
  wire tmp5536;
  wire tmp5537;
  wire tmp5538;
  wire tmp5539;
  wire tmp5540;
  wire tmp5541;
  wire tmp5542;
  wire tmp5543;
  wire tmp5544;
  wire tmp5545;
  wire tmp5546;
  wire tmp5547;
  wire tmp5548;
  wire tmp5549;
  wire tmp5550;
  wire tmp5551;
  wire tmp5552;
  wire tmp5553;
  wire tmp5554;
  wire tmp5555;
  wire tmp5556;
  wire tmp5557;
  wire tmp5558;
  wire tmp5559;
  wire tmp5560;
  wire tmp5561;
  wire tmp5562;
  wire tmp5563;
  wire tmp5564;
  wire tmp5565;
  wire tmp5566;
  wire tmp5567;
  wire tmp5568;
  wire tmp5569;
  wire tmp5570;
  wire tmp5571;
  wire tmp5572;
  wire tmp5573;
  wire tmp5574;
  wire tmp5575;
  wire tmp5576;
  wire tmp5577;
  wire tmp5578;
  wire tmp5579;
  wire tmp5580;
  wire tmp5581;
  wire tmp5582;
  wire tmp5583;
  wire tmp5584;
  wire tmp5585;
  wire tmp5586;
  wire tmp5587;
  wire tmp5588;
  wire tmp5589;
  wire tmp5590;
  wire tmp5591;
  wire tmp5592;
  wire tmp5593;
  wire tmp5594;
  wire tmp5595;
  wire tmp5596;
  wire tmp5597;
  wire tmp5598;
  wire tmp5599;
  wire tmp5600;
  wire tmp5601;
  wire tmp5602;
  wire tmp5603;
  wire tmp5604;
  wire tmp5605;
  wire tmp5606;
  wire tmp5607;
  wire tmp5608;
  wire tmp5609;
  wire tmp5610;
  wire tmp5611;
  wire tmp5612;
  wire tmp5613;
  wire tmp5614;
  wire tmp5615;
  wire tmp5616;
  wire tmp5617;
  wire tmp5618;
  wire tmp5619;
  wire tmp5620;
  wire tmp5621;
  wire tmp5622;
  wire tmp5623;
  wire tmp5624;
  wire tmp5625;
  wire tmp5626;
  wire tmp5627;
  wire tmp5628;
  wire tmp5629;
  wire tmp5630;
  wire tmp5631;
  wire tmp5632;
  wire tmp5633;
  wire tmp5634;
  wire tmp5635;
  wire tmp5636;
  wire tmp5637;
  wire tmp5638;
  wire tmp5639;
  wire tmp5640;
  wire tmp5641;
  wire tmp5642;
  wire tmp5643;
  wire tmp5644;
  wire tmp5645;
  wire tmp5646;
  wire tmp5647;
  wire tmp5648;
  wire tmp5649;
  wire tmp5650;
  wire tmp5651;
  wire tmp5652;
  wire tmp5653;
  wire tmp5654;
  wire tmp5655;
  wire tmp5656;
  wire tmp5657;
  wire tmp5658;
  wire tmp5659;
  wire tmp5660;
  wire tmp5661;
  wire tmp5662;
  wire tmp5663;
  wire tmp5664;
  wire tmp5665;
  wire tmp5666;
  wire tmp5667;
  wire tmp5668;
  wire tmp5669;
  wire tmp5670;
  wire tmp5671;
  wire tmp5672;
  wire tmp5673;
  wire tmp5674;
  wire tmp5675;
  wire tmp5676;
  wire tmp5677;
  wire tmp5678;
  wire tmp5679;
  wire tmp5680;
  wire tmp5681;
  wire tmp5682;
  wire tmp5683;
  wire tmp5684;
  wire tmp5685;
  wire tmp5686;
  wire tmp5687;
  wire tmp5688;
  wire tmp5689;
  wire tmp5690;
  wire tmp5691;
  wire tmp5692;
  wire tmp5693;
  wire tmp5694;
  wire tmp5695;
  wire tmp5696;
  wire tmp5697;
  wire tmp5698;
  wire tmp5699;
  wire tmp5700;
  wire tmp5701;
  wire tmp5702;
  wire tmp5703;
  wire tmp5704;
  wire tmp5705;
  wire tmp5706;
  wire tmp5707;
  wire tmp5708;
  wire tmp5709;
  wire tmp5710;
  wire tmp5711;
  wire tmp5712;
  wire tmp5713;
  wire tmp5714;
  wire tmp5715;
  wire tmp5716;
  wire tmp5717;
  wire tmp5718;
  wire tmp5719;
  wire tmp5720;
  wire tmp5721;
  wire tmp5722;
  wire tmp5723;
  wire tmp5724;
  wire tmp5725;
  wire tmp5726;
  wire tmp5727;
  wire tmp5728;
  wire tmp5729;
  wire tmp5730;
  wire tmp5731;
  wire tmp5732;
  wire tmp5733;
  wire tmp5734;
  wire tmp5735;
  wire tmp5736;
  wire tmp5737;
  wire tmp5738;
  wire tmp5739;
  wire tmp5740;
  wire tmp5741;
  wire tmp5742;
  wire tmp5743;
  wire tmp5744;
  wire tmp5745;
  wire tmp5746;
  wire tmp5747;
  wire tmp5748;
  wire tmp5749;
  wire tmp5750;
  wire tmp5751;
  wire tmp5752;
  wire tmp5753;
  wire tmp5754;
  wire tmp5755;
  wire tmp5756;
  wire tmp5757;
  wire tmp5758;
  wire tmp5759;
  wire tmp5760;
  wire tmp5761;
  wire tmp5762;
  wire tmp5763;
  wire tmp5764;
  wire tmp5765;
  wire tmp5766;
  wire tmp5767;
  wire tmp5768;
  wire tmp5769;
  wire tmp5770;
  wire tmp5771;
  wire tmp5772;
  wire tmp5773;
  wire tmp5774;
  wire tmp5775;
  wire tmp5776;
  wire tmp5777;
  wire tmp5778;
  wire tmp5779;
  wire tmp5780;
  wire tmp5781;
  wire tmp5782;
  wire tmp5783;
  wire tmp5784;
  wire tmp5785;
  wire tmp5786;
  wire tmp5787;
  wire tmp5788;
  wire tmp5789;
  wire tmp5790;
  wire tmp5791;
  wire tmp5792;
  wire tmp5793;
  wire tmp5794;
  wire tmp5795;
  wire tmp5796;
  wire tmp5797;
  wire tmp5798;
  wire tmp5799;
  wire tmp5800;
  wire tmp5801;
  wire tmp5802;
  wire tmp5803;
  wire tmp5804;
  wire tmp5805;
  wire tmp5806;
  wire tmp5807;
  wire tmp5808;
  wire tmp5809;
  wire tmp5810;
  wire tmp5811;
  wire tmp5812;
  wire tmp5813;
  wire tmp5814;
  wire tmp5815;
  wire tmp5816;
  wire tmp5817;
  wire tmp5818;
  wire tmp5819;
  wire tmp5820;
  wire tmp5821;
  wire tmp5822;
  wire tmp5823;
  wire tmp5824;
  wire tmp5825;
  wire tmp5826;
  wire tmp5827;
  wire tmp5828;
  wire tmp5829;
  wire tmp5830;
  wire tmp5831;
  wire tmp5832;
  wire tmp5833;
  wire tmp5834;
  wire tmp5835;
  wire tmp5836;
  wire tmp5837;
  wire tmp5838;
  wire tmp5839;
  wire tmp5840;
  wire tmp5841;
  wire tmp5842;
  wire tmp5843;
  wire tmp5844;
  wire tmp5845;
  wire tmp5846;
  wire tmp5847;
  wire tmp5848;
  wire tmp5849;
  wire tmp5850;
  wire tmp5851;
  wire tmp5852;
  wire tmp5853;
  wire tmp5854;
  wire tmp5855;
  wire tmp5856;
  wire tmp5857;
  wire tmp5858;
  wire tmp5859;
  wire tmp5860;
  wire tmp5861;
  wire tmp5862;
  wire tmp5863;
  wire tmp5864;
  wire tmp5865;
  wire tmp5866;
  wire tmp5867;
  wire tmp5868;
  wire tmp5869;
  wire tmp5870;
  wire tmp5871;
  wire tmp5872;
  wire tmp5873;
  wire tmp5874;
  wire tmp5875;
  wire tmp5876;
  wire tmp5877;
  wire tmp5878;
  wire tmp5879;
  wire tmp5880;
  wire tmp5881;
  wire tmp5882;
  wire tmp5883;
  wire tmp5884;
  wire tmp5885;
  wire tmp5886;
  wire tmp5887;
  wire tmp5888;
  wire tmp5889;
  wire tmp5890;
  wire tmp5891;
  wire tmp5892;
  wire tmp5893;
  wire tmp5894;
  wire tmp5895;
  wire tmp5896;
  wire tmp5897;
  wire tmp5898;
  wire tmp5899;
  wire tmp5900;
  wire tmp5901;
  wire tmp5902;
  wire tmp5903;
  wire tmp5904;
  wire tmp5905;
  wire tmp5906;
  wire tmp5907;
  wire tmp5908;
  wire tmp5909;
  wire tmp5910;
  wire tmp5911;
  wire tmp5912;
  wire tmp5913;
  wire tmp5914;
  wire tmp5915;
  wire tmp5916;
  wire tmp5917;
  wire tmp5918;
  wire tmp5919;
  wire tmp5920;
  wire tmp5921;
  wire tmp5922;
  wire tmp5923;
  wire tmp5924;
  wire tmp5925;
  wire tmp5926;
  wire tmp5927;
  wire tmp5928;
  wire tmp5929;
  wire tmp5930;
  wire tmp5931;
  wire tmp5932;
  wire tmp5933;
  wire tmp5934;
  wire tmp5935;
  wire tmp5936;
  wire tmp5937;
  wire tmp5938;
  wire tmp5939;
  wire tmp5940;
  wire tmp5941;
  wire tmp5942;
  wire tmp5943;
  wire tmp5944;
  wire tmp5945;
  wire tmp5946;
  wire tmp5947;
  wire tmp5948;
  wire tmp5949;
  wire tmp5950;
  wire tmp5951;
  wire tmp5952;
  wire tmp5953;
  wire tmp5954;
  wire tmp5955;
  wire tmp5956;
  wire tmp5957;
  wire tmp5958;
  wire tmp5959;
  wire tmp5960;
  wire tmp5961;
  wire tmp5962;
  wire tmp5963;
  wire tmp5964;
  wire tmp5965;
  wire tmp5966;
  wire tmp5967;
  wire tmp5968;
  wire tmp5969;
  wire tmp5970;
  wire tmp5971;
  wire tmp5972;
  wire tmp5973;
  wire tmp5974;
  wire tmp5975;
  wire tmp5976;
  wire tmp5977;
  wire tmp5978;
  wire tmp5979;
  wire tmp5980;
  wire tmp5981;
  wire tmp5982;
  wire tmp5983;
  wire tmp5984;
  wire tmp5985;
  wire tmp5986;
  wire tmp5987;
  wire tmp5988;
  wire tmp5989;
  wire tmp5990;
  wire tmp5991;
  wire tmp5992;
  wire tmp5993;
  wire tmp5994;
  wire tmp5995;
  wire tmp5996;
  wire tmp5997;
  wire tmp5998;
  wire tmp5999;
  wire tmp6000;
  wire tmp6001;
  wire tmp6002;
  wire tmp6003;
  wire tmp6004;
  wire tmp6005;
  wire tmp6006;
  wire tmp6007;
  wire tmp6008;
  wire tmp6009;
  wire tmp6010;
  wire tmp6011;
  wire tmp6012;
  wire tmp6013;
  wire tmp6014;
  wire tmp6015;
  wire tmp6016;
  wire tmp6017;
  wire tmp6018;
  wire tmp6019;
  wire tmp6020;
  wire tmp6021;
  wire tmp6022;
  wire tmp6023;
  wire tmp6024;
  wire tmp6025;
  wire tmp6026;
  wire tmp6027;
  wire tmp6028;
  wire tmp6029;
  wire tmp6030;
  wire tmp6031;
  wire tmp6032;
  wire tmp6033;
  wire tmp6034;
  wire tmp6035;
  wire tmp6036;
  wire tmp6037;
  wire tmp6038;
  wire tmp6039;
  wire tmp6040;
  wire tmp6041;
  wire tmp6042;
  wire tmp6043;
  wire tmp6044;
  wire tmp6045;
  wire tmp6046;
  wire tmp6047;
  wire tmp6048;
  wire tmp6049;
  wire tmp6050;
  wire tmp6051;
  wire tmp6052;
  wire tmp6053;
  wire tmp6054;
  wire tmp6055;
  wire tmp6056;
  wire tmp6057;
  wire tmp6058;
  wire tmp6059;
  wire tmp6060;
  wire tmp6061;
  wire tmp6062;
  wire tmp6063;
  wire tmp6064;
  wire tmp6065;
  wire tmp6066;
  wire tmp6067;
  wire tmp6068;
  wire tmp6069;
  wire tmp6070;
  wire tmp6071;
  wire tmp6072;
  wire tmp6073;
  wire tmp6074;
  wire tmp6075;
  wire tmp6076;
  wire tmp6077;
  wire tmp6078;
  wire tmp6079;
  wire tmp6080;
  wire tmp6081;
  wire tmp6082;
  wire tmp6083;
  wire tmp6084;
  wire tmp6085;
  wire tmp6086;
  wire tmp6087;
  wire tmp6088;
  wire tmp6089;
  wire tmp6090;
  wire tmp6091;
  wire tmp6092;
  wire tmp6093;
  wire tmp6094;
  wire tmp6095;
  wire tmp6096;
  wire tmp6097;
  wire tmp6098;
  wire tmp6099;
  wire tmp6100;
  wire tmp6101;
  wire tmp6102;
  wire tmp6103;
  wire tmp6104;
  wire tmp6105;
  wire tmp6106;
  wire tmp6107;
  wire tmp6108;
  wire tmp6109;
  wire tmp6110;
  wire tmp6111;
  wire tmp6112;
  wire tmp6113;
  wire tmp6114;
  wire tmp6115;
  wire tmp6116;
  wire tmp6117;
  wire tmp6118;
  wire tmp6119;
  wire tmp6120;
  wire tmp6121;
  wire tmp6122;
  wire tmp6123;
  wire tmp6124;
  wire tmp6125;
  wire tmp6126;
  wire tmp6127;
  wire tmp6128;
  wire tmp6129;
  wire tmp6130;
  wire tmp6131;
  wire tmp6132;
  wire tmp6133;
  wire tmp6134;
  wire tmp6135;
  wire tmp6136;
  wire tmp6137;
  wire tmp6138;
  wire tmp6139;
  wire tmp6140;
  wire tmp6141;
  wire tmp6142;
  wire tmp6143;
  wire tmp6144;
  wire tmp6145;
  wire tmp6146;
  wire tmp6147;
  wire tmp6148;
  wire tmp6149;
  wire tmp6150;
  wire tmp6151;
  wire tmp6152;
  wire tmp6153;
  wire tmp6154;
  wire tmp6155;
  wire tmp6156;
  wire tmp6157;
  wire tmp6158;
  wire tmp6159;
  wire tmp6160;
  wire tmp6161;
  wire tmp6162;
  wire tmp6163;
  wire tmp6164;
  wire tmp6165;
  wire tmp6166;
  wire tmp6167;
  wire tmp6168;
  wire tmp6169;
  wire tmp6170;
  wire tmp6171;
  wire tmp6172;
  wire tmp6173;
  wire tmp6174;
  wire tmp6175;
  wire tmp6176;
  wire tmp6177;
  wire tmp6178;
  wire tmp6179;
  wire tmp6180;
  wire tmp6181;
  wire tmp6182;
  wire tmp6183;
  wire tmp6184;
  wire tmp6185;
  wire tmp6186;
  wire tmp6187;
  wire tmp6188;
  wire tmp6189;
  wire tmp6190;
  wire tmp6191;
  wire tmp6192;
  wire tmp6193;
  wire tmp6194;
  wire tmp6195;
  wire tmp6196;
  wire tmp6197;
  wire tmp6198;
  wire tmp6199;
  wire tmp6200;
  wire tmp6201;
  wire tmp6202;
  wire tmp6203;
  wire tmp6204;
  wire tmp6205;
  wire tmp6206;
  wire tmp6207;
  wire tmp6208;
  wire tmp6209;
  wire tmp6210;
  wire tmp6211;
  wire tmp6212;
  wire tmp6213;
  wire tmp6214;
  wire tmp6215;
  wire tmp6216;
  wire tmp6217;
  wire tmp6218;
  wire tmp6219;
  wire tmp6220;
  wire tmp6221;
  wire tmp6222;
  wire tmp6223;
  wire tmp6224;
  wire tmp6225;
  wire tmp6226;
  wire tmp6227;
  wire tmp6228;
  wire tmp6229;
  wire tmp6230;
  wire tmp6231;
  wire tmp6232;
  wire tmp6233;
  wire tmp6234;
  wire tmp6235;
  wire tmp6236;
  wire tmp6237;
  wire tmp6238;
  wire tmp6239;
  wire tmp6240;
  wire tmp6241;
  wire tmp6242;
  wire tmp6243;
  wire tmp6244;
  wire tmp6245;
  wire tmp6246;
  wire tmp6247;
  wire tmp6248;
  wire tmp6249;
  wire tmp6250;
  wire tmp6251;
  wire tmp6252;
  wire tmp6253;
  wire tmp6254;
  wire tmp6255;
  wire tmp6256;
  wire tmp6257;
  wire tmp6258;
  wire tmp6259;
  wire tmp6260;
  wire tmp6261;
  wire tmp6262;
  wire tmp6263;
  wire tmp6264;
  wire tmp6265;
  wire tmp6266;
  wire tmp6267;
  wire tmp6268;
  wire tmp6269;
  wire tmp6270;
  wire tmp6271;
  wire tmp6272;
  wire tmp6273;
  wire tmp6274;
  wire tmp6275;
  wire tmp6276;
  wire tmp6277;
  wire tmp6278;
  wire tmp6279;
  wire tmp6280;
  wire tmp6281;
  wire tmp6282;
  wire tmp6283;
  wire tmp6284;
  wire tmp6285;
  wire tmp6286;
  wire tmp6287;
  wire tmp6288;
  wire tmp6289;
  wire tmp6290;
  wire tmp6291;
  wire tmp6292;
  wire tmp6293;
  wire tmp6294;
  wire tmp6295;
  wire tmp6296;
  wire tmp6297;
  wire tmp6298;
  wire tmp6299;
  wire tmp6300;
  wire tmp6301;
  wire tmp6302;
  wire tmp6303;
  wire tmp6304;
  wire tmp6305;
  wire tmp6306;
  wire tmp6307;
  wire tmp6308;
  wire tmp6309;
  wire tmp6310;
  wire tmp6311;
  wire tmp6312;
  wire tmp6313;
  wire tmp6314;
  wire tmp6315;
  wire tmp6316;
  wire tmp6317;
  wire tmp6318;
  wire tmp6319;
  wire tmp6320;
  wire tmp6321;
  wire tmp6322;
  wire tmp6323;
  wire tmp6324;
  wire tmp6325;
  wire tmp6326;
  wire tmp6327;
  wire tmp6328;
  wire tmp6329;
  wire tmp6330;
  wire tmp6331;
  wire tmp6332;
  wire tmp6333;
  wire tmp6334;
  wire tmp6335;
  wire tmp6336;
  wire tmp6337;
  wire tmp6338;
  wire tmp6339;
  wire tmp6340;
  wire tmp6341;
  wire tmp6342;
  wire tmp6343;
  wire tmp6344;
  wire tmp6345;
  wire tmp6346;
  wire tmp6347;
  wire tmp6348;
  wire tmp6349;
  wire tmp6350;
  wire tmp6351;
  wire tmp6352;
  wire tmp6353;
  wire tmp6354;
  wire tmp6355;
  wire tmp6356;
  wire tmp6357;
  wire tmp6358;
  wire tmp6359;
  wire tmp6360;
  wire tmp6361;
  wire tmp6362;
  wire tmp6363;
  wire tmp6364;
  wire tmp6365;
  wire tmp6366;
  wire tmp6367;
  wire tmp6368;
  wire tmp6369;
  wire tmp6370;
  wire tmp6371;
  wire tmp6372;
  wire tmp6373;
  wire tmp6374;
  wire tmp6375;
  wire tmp6376;
  wire tmp6377;
  wire tmp6378;
  wire tmp6379;
  wire tmp6380;
  wire tmp6381;
  wire tmp6382;
  wire tmp6383;
  wire tmp6384;
  wire tmp6385;
  wire tmp6386;
  wire tmp6387;
  wire tmp6388;
  wire tmp6389;
  wire tmp6390;
  wire tmp6391;
  wire tmp6392;
  wire tmp6393;
  wire tmp6394;
  wire tmp6395;
  wire tmp6396;
  wire tmp6397;
  wire tmp6398;
  wire tmp6399;
  wire tmp6400;
  wire tmp6401;
  wire tmp6402;
  wire tmp6403;
  wire tmp6404;
  wire tmp6405;
  wire tmp6406;
  wire tmp6407;
  wire tmp6408;
  wire tmp6409;
  wire tmp6410;
  wire tmp6411;
  wire tmp6412;
  wire tmp6413;
  wire tmp6414;
  wire tmp6415;
  wire tmp6416;
  wire tmp6417;
  wire tmp6418;
  wire tmp6419;
  wire tmp6420;
  wire tmp6421;
  wire tmp6422;
  wire tmp6423;
  wire tmp6424;
  wire tmp6425;
  wire tmp6426;
  wire tmp6427;
  wire tmp6428;
  wire tmp6429;
  wire tmp6430;
  wire tmp6431;
  wire tmp6432;
  wire tmp6433;
  wire tmp6434;
  wire tmp6435;
  wire tmp6436;
  wire tmp6437;
  wire tmp6438;
  wire tmp6439;
  wire tmp6440;
  wire tmp6441;
  wire tmp6442;
  wire tmp6443;
  wire tmp6444;
  wire tmp6445;
  wire tmp6446;
  wire tmp6447;
  wire tmp6448;
  wire tmp6449;
  wire tmp6450;
  wire tmp6451;
  wire tmp6452;
  wire tmp6453;
  wire tmp6454;
  wire tmp6455;
  wire tmp6456;
  wire tmp6457;
  wire tmp6458;
  wire tmp6459;
  wire tmp6460;
  wire tmp6461;
  wire tmp6462;
  wire tmp6463;
  wire tmp6464;
  wire tmp6465;
  wire tmp6466;
  wire tmp6467;
  wire tmp6468;
  wire tmp6469;
  wire tmp6470;
  wire tmp6471;
  wire tmp6472;
  wire tmp6473;
  wire tmp6474;
  wire tmp6475;
  wire tmp6476;
  wire tmp6477;
  wire tmp6478;
  wire tmp6479;
  wire tmp6480;
  wire tmp6481;
  wire tmp6482;
  wire tmp6483;
  wire tmp6484;
  wire tmp6485;
  wire tmp6486;
  wire tmp6487;
  wire tmp6488;
  wire tmp6489;
  wire tmp6490;
  wire tmp6491;
  wire tmp6492;
  wire tmp6493;
  wire tmp6494;
  wire tmp6495;
  wire tmp6496;
  wire tmp6497;
  wire tmp6498;
  wire tmp6499;
  wire tmp6500;
  wire tmp6501;
  wire tmp6502;
  wire tmp6503;
  wire tmp6504;
  wire tmp6505;
  wire tmp6506;
  wire tmp6507;
  wire tmp6508;
  wire tmp6509;
  wire tmp6510;
  wire tmp6511;
  wire tmp6512;
  wire tmp6513;
  wire tmp6514;
  wire tmp6515;
  wire tmp6516;
  wire tmp6517;
  wire tmp6518;
  wire tmp6519;
  wire tmp6520;
  wire tmp6521;
  wire tmp6522;
  wire tmp6523;
  wire tmp6524;
  wire tmp6525;
  wire tmp6526;
  wire tmp6527;
  wire tmp6528;
  wire tmp6529;
  wire tmp6530;
  wire tmp6531;
  wire tmp6532;
  wire tmp6533;
  wire tmp6534;
  wire tmp6535;
  wire tmp6536;
  wire tmp6537;
  wire tmp6538;
  wire tmp6539;
  wire tmp6540;
  wire tmp6541;
  wire tmp6542;
  wire tmp6543;
  wire tmp6544;
  wire tmp6545;
  wire tmp6546;
  wire tmp6547;
  wire tmp6548;
  wire tmp6549;
  wire tmp6550;
  wire tmp6551;
  wire tmp6552;
  wire tmp6553;
  wire tmp6554;
  wire tmp6555;
  wire tmp6556;
  wire tmp6557;
  wire tmp6558;
  wire tmp6559;
  wire tmp6560;
  wire tmp6561;
  wire tmp6562;
  wire tmp6563;
  wire tmp6564;
  wire tmp6565;
  wire tmp6566;
  wire tmp6567;
  wire tmp6568;
  wire tmp6569;
  wire tmp6570;
  wire tmp6571;
  wire tmp6572;
  wire tmp6573;
  wire tmp6574;
  wire tmp6575;
  wire tmp6576;
  wire tmp6577;
  wire tmp6578;
  wire tmp6579;
  wire tmp6580;
  wire tmp6581;
  wire tmp6582;
  wire tmp6583;
  wire tmp6584;
  wire tmp6585;
  wire tmp6586;
  wire tmp6587;
  wire tmp6588;
  wire tmp6589;
  wire tmp6590;
  wire tmp6591;
  wire tmp6592;
  wire tmp6593;
  wire tmp6594;
  wire tmp6595;
  wire tmp6596;
  wire tmp6597;
  wire tmp6598;
  wire tmp6599;
  wire tmp6600;
  wire tmp6601;
  wire tmp6602;
  wire tmp6603;
  wire tmp6604;
  wire tmp6605;
  wire tmp6606;
  wire tmp6607;
  wire tmp6608;
  wire tmp6609;
  wire tmp6610;
  wire tmp6611;
  wire tmp6612;
  wire tmp6613;
  wire tmp6614;
  wire tmp6615;
  wire tmp6616;
  wire tmp6617;
  wire tmp6618;
  wire tmp6619;
  wire tmp6620;
  wire tmp6621;
  wire tmp6622;
  wire tmp6623;
  wire tmp6624;
  wire tmp6625;
  wire tmp6626;
  wire tmp6627;
  wire tmp6628;
  wire tmp6629;
  wire tmp6630;
  wire tmp6631;
  wire tmp6632;
  wire tmp6633;
  wire tmp6634;
  wire tmp6635;
  wire tmp6636;
  wire tmp6637;
  wire tmp6638;
  wire tmp6639;
  wire tmp6640;
  wire tmp6641;
  wire tmp6642;
  wire tmp6643;
  wire tmp6644;
  wire tmp6645;
  wire tmp6646;
  wire tmp6647;
  wire tmp6648;
  wire tmp6649;
  wire tmp6650;
  wire tmp6651;
  wire tmp6652;
  wire tmp6653;
  wire tmp6654;
  wire tmp6655;
  wire tmp6656;
  wire tmp6657;
  wire tmp6658;
  wire tmp6659;
  wire tmp6660;
  wire tmp6661;
  wire tmp6662;
  wire tmp6663;
  wire tmp6664;
  wire tmp6665;
  wire tmp6666;
  wire tmp6667;
  wire tmp6668;
  wire tmp6669;
  wire tmp6670;
  wire tmp6671;
  wire tmp6672;
  wire tmp6673;
  wire tmp6674;
  wire tmp6675;
  wire tmp6676;
  wire tmp6677;
  wire tmp6678;
  wire tmp6679;
  wire tmp6680;
  wire tmp6681;
  wire tmp6682;
  wire tmp6683;
  wire tmp6684;
  wire tmp6685;
  wire tmp6686;
  wire tmp6687;
  wire tmp6688;
  wire tmp6689;
  wire tmp6690;
  wire tmp6691;
  wire tmp6692;
  wire tmp6693;
  wire tmp6694;
  wire tmp6695;
  wire tmp6696;
  wire tmp6697;
  wire tmp6698;
  wire tmp6699;
  wire tmp6700;
  wire tmp6701;
  wire tmp6702;
  wire tmp6703;
  wire tmp6704;
  wire tmp6705;
  wire tmp6706;
  wire tmp6707;
  wire tmp6708;
  wire tmp6709;
  wire tmp6710;
  wire tmp6711;
  wire tmp6712;
  wire tmp6713;
  wire tmp6714;
  wire tmp6715;
  wire tmp6716;
  wire tmp6717;
  wire tmp6718;
  wire tmp6719;
  wire tmp6720;
  wire tmp6721;
  wire tmp6722;
  wire tmp6723;
  wire tmp6724;
  wire tmp6725;
  wire tmp6726;
  wire tmp6727;
  wire tmp6728;
  wire tmp6729;
  wire tmp6730;
  wire tmp6731;
  wire tmp6732;
  wire tmp6733;
  wire tmp6734;
  wire tmp6735;
  wire tmp6736;
  wire tmp6737;
  wire tmp6738;
  wire tmp6739;
  wire tmp6740;
  wire tmp6741;
  wire tmp6742;
  wire tmp6743;
  wire tmp6744;
  wire tmp6745;
  wire tmp6746;
  wire tmp6747;
  wire tmp6748;
  wire tmp6749;
  wire tmp6750;
  wire tmp6751;
  wire tmp6752;
  wire tmp6753;
  wire tmp6754;
  wire tmp6755;
  wire tmp6756;
  wire tmp6757;
  wire tmp6758;
  wire tmp6759;
  wire tmp6760;
  wire tmp6761;
  wire tmp6762;
  wire tmp6763;
  wire tmp6764;
  wire tmp6765;
  wire tmp6766;
  wire tmp6767;
  wire tmp6768;
  wire tmp6769;
  wire tmp6770;
  wire tmp6771;
  wire tmp6772;
  wire tmp6773;
  wire tmp6774;
  wire tmp6775;
  wire tmp6776;
  wire tmp6777;
  wire tmp6778;
  wire tmp6779;
  wire tmp6780;
  wire tmp6781;
  wire tmp6782;
  wire tmp6783;
  wire tmp6784;
  wire tmp6785;
  wire tmp6786;
  wire tmp6787;
  wire tmp6788;
  wire tmp6789;
  wire tmp6790;
  wire tmp6791;
  wire tmp6792;
  wire tmp6793;
  wire tmp6794;
  wire tmp6795;
  wire tmp6796;
  wire tmp6797;
  wire tmp6798;
  wire tmp6799;
  wire tmp6800;
  wire tmp6801;
  wire tmp6802;
  wire tmp6803;
  wire tmp6804;
  wire tmp6805;
  wire tmp6806;
  wire tmp6807;
  wire tmp6808;
  wire tmp6809;
  wire tmp6810;
  wire tmp6811;
  wire tmp6812;
  wire tmp6813;
  wire tmp6814;
  wire tmp6815;
  wire tmp6816;
  wire tmp6817;
  wire tmp6818;
  wire tmp6819;
  wire tmp6820;
  wire tmp6821;
  wire tmp6822;
  wire tmp6823;
  wire tmp6824;
  wire tmp6825;
  wire tmp6826;
  wire tmp6827;
  wire tmp6828;
  wire tmp6829;
  wire tmp6830;
  wire tmp6831;
  wire tmp6832;
  wire tmp6833;
  wire tmp6834;
  wire tmp6835;
  wire tmp6836;
  wire tmp6837;
  wire tmp6838;
  wire tmp6839;
  wire tmp6840;
  wire tmp6841;
  wire tmp6842;
  wire tmp6843;
  wire tmp6844;
  wire tmp6845;
  wire tmp6846;
  wire tmp6847;
  wire tmp6848;
  wire tmp6849;
  wire tmp6850;
  wire tmp6851;
  wire tmp6852;
  wire tmp6853;
  wire tmp6854;
  wire tmp6855;
  wire tmp6856;
  wire tmp6857;
  wire tmp6858;
  wire tmp6859;
  wire tmp6860;
  wire tmp6861;
  wire tmp6862;
  wire tmp6863;
  wire tmp6864;
  wire tmp6865;
  wire tmp6866;
  wire tmp6867;
  wire tmp6868;
  wire tmp6869;
  wire tmp6870;
  wire tmp6871;
  wire tmp6872;
  wire tmp6873;
  wire tmp6874;
  wire tmp6875;
  wire tmp6876;
  wire tmp6877;
  wire tmp6878;
  wire tmp6879;
  wire tmp6880;
  wire tmp6881;
  wire tmp6882;
  wire tmp6883;
  wire tmp6884;
  wire tmp6885;
  wire tmp6886;
  wire tmp6887;
  wire tmp6888;
  wire tmp6889;
  wire tmp6890;
  wire tmp6891;
  wire tmp6892;
  wire tmp6893;
  wire tmp6894;
  wire tmp6895;
  wire tmp6896;
  wire tmp6897;
  wire tmp6898;
  wire tmp6899;
  wire tmp6900;
  wire tmp6901;
  wire tmp6902;
  wire tmp6903;
  wire tmp6904;
  wire tmp6905;
  wire tmp6906;
  wire tmp6907;
  wire tmp6908;
  wire tmp6909;
  wire tmp6910;
  wire tmp6911;
  wire tmp6912;
  wire tmp6913;
  wire tmp6914;
  wire tmp6915;
  wire tmp6916;
  wire tmp6917;
  wire tmp6918;
  wire tmp6919;
  wire tmp6920;
  wire tmp6921;
  wire tmp6922;
  wire tmp6923;
  wire tmp6924;
  wire tmp6925;
  wire tmp6926;
  wire tmp6927;
  wire tmp6928;
  wire tmp6929;
  wire tmp6930;
  wire tmp6931;
  wire tmp6932;
  wire tmp6933;
  wire tmp6934;
  wire tmp6935;
  wire tmp6936;
  wire tmp6937;
  wire tmp6938;
  wire tmp6939;
  wire tmp6940;
  wire tmp6941;
  wire tmp6942;
  wire tmp6943;
  wire tmp6944;
  wire tmp6945;
  wire tmp6946;
  wire tmp6947;
  wire tmp6948;
  wire tmp6949;
  wire tmp6950;
  wire tmp6951;
  wire tmp6952;
  wire tmp6953;
  wire tmp6954;
  wire tmp6955;
  wire tmp6956;
  wire tmp6957;
  wire tmp6958;
  wire tmp6959;
  wire tmp6960;
  wire tmp6961;
  wire tmp6962;
  wire tmp6963;
  wire tmp6964;
  wire tmp6965;
  wire tmp6966;
  wire tmp6967;
  wire tmp6968;
  wire tmp6969;
  wire tmp6970;
  wire tmp6971;
  wire tmp6972;
  wire tmp6973;
  wire tmp6974;
  wire tmp6975;
  wire tmp6976;
  wire tmp6977;
  wire tmp6978;
  wire tmp6979;
  wire tmp6980;
  wire tmp6981;
  wire tmp6982;
  wire tmp6983;
  wire tmp6984;
  wire tmp6985;
  wire tmp6986;
  wire tmp6987;
  wire tmp6988;
  wire tmp6989;
  wire tmp6990;
  wire tmp6991;
  wire tmp6992;
  wire tmp6993;
  wire tmp6994;
  wire tmp6995;
  wire tmp6996;
  wire tmp6997;
  wire tmp6998;
  wire tmp6999;
  wire tmp7000;
  wire tmp7001;
  wire tmp7002;
  wire tmp7003;
  wire tmp7004;
  wire tmp7005;
  wire tmp7006;
  wire tmp7007;
  wire tmp7008;
  wire tmp7009;
  wire tmp7010;
  wire tmp7011;
  wire tmp7012;
  wire tmp7013;
  wire tmp7014;
  wire tmp7015;
  wire tmp7016;
  wire tmp7017;
  wire tmp7018;
  wire tmp7019;
  wire tmp7020;
  wire tmp7021;
  wire tmp7022;
  wire tmp7023;
  wire tmp7024;
  wire tmp7025;
  wire tmp7026;
  wire tmp7027;
  wire tmp7028;
  wire tmp7029;
  wire tmp7030;
  wire tmp7031;
  wire tmp7032;
  wire tmp7033;
  wire tmp7034;
  wire tmp7035;
  wire tmp7036;
  wire tmp7037;
  wire tmp7038;
  wire tmp7039;
  wire tmp7040;
  wire tmp7041;
  wire tmp7042;
  wire tmp7043;
  wire tmp7044;
  wire tmp7045;
  wire tmp7046;
  wire tmp7047;
  wire tmp7048;
  wire tmp7049;
  wire tmp7050;
  wire tmp7051;
  wire tmp7052;
  wire tmp7053;
  wire tmp7054;
  wire tmp7055;
  wire tmp7056;
  wire tmp7057;
  wire tmp7058;
  wire tmp7059;
  wire tmp7060;
  wire tmp7061;
  wire tmp7062;
  wire tmp7063;
  wire tmp7064;
  wire tmp7065;
  wire tmp7066;
  wire tmp7067;
  wire tmp7068;
  wire tmp7069;
  wire tmp7070;
  wire tmp7071;
  wire tmp7072;
  wire tmp7073;
  wire tmp7074;
  wire tmp7075;
  wire tmp7076;
  wire tmp7077;
  wire tmp7078;
  wire tmp7079;
  wire tmp7080;
  wire tmp7081;
  wire tmp7082;
  wire tmp7083;
  wire tmp7084;
  wire tmp7085;
  wire tmp7086;
  wire tmp7087;
  wire tmp7088;
  wire tmp7089;
  wire tmp7090;
  wire tmp7091;
  wire tmp7092;
  wire tmp7093;
  wire tmp7094;
  wire tmp7095;
  wire tmp7096;
  wire tmp7097;
  wire tmp7098;
  wire tmp7099;
  wire tmp7100;
  wire tmp7101;
  wire tmp7102;
  wire tmp7103;
  wire tmp7104;
  wire tmp7105;
  wire tmp7106;
  wire tmp7107;
  wire tmp7108;
  wire tmp7109;
  wire tmp7110;
  wire tmp7111;
  wire tmp7112;
  wire tmp7113;
  wire tmp7114;
  wire tmp7115;
  wire tmp7116;
  wire tmp7117;
  wire tmp7118;
  wire tmp7119;
  wire tmp7120;
  wire tmp7121;
  wire tmp7122;
  wire tmp7123;
  wire tmp7124;
  wire tmp7125;
  wire tmp7126;
  wire tmp7127;
  wire tmp7128;
  wire tmp7129;
  wire tmp7130;
  wire tmp7131;
  wire tmp7132;
  wire tmp7133;
  wire tmp7134;
  wire tmp7135;
  wire tmp7136;
  wire tmp7137;
  wire tmp7138;
  wire tmp7139;
  wire tmp7140;
  wire tmp7141;
  wire tmp7142;
  wire tmp7143;
  wire tmp7144;
  wire tmp7145;
  wire tmp7146;
  wire tmp7147;
  wire tmp7148;
  wire tmp7149;
  wire tmp7150;
  wire tmp7151;
  wire tmp7152;
  wire tmp7153;
  wire tmp7154;
  wire tmp7155;
  wire tmp7156;
  wire tmp7157;
  wire tmp7158;
  wire tmp7159;
  wire tmp7160;
  wire tmp7161;
  wire tmp7162;
  wire tmp7163;
  wire tmp7164;
  wire tmp7165;
  wire tmp7166;
  wire tmp7167;
  wire tmp7168;
  wire tmp7169;
  wire tmp7170;
  wire tmp7171;
  wire tmp7172;
  wire tmp7173;
  wire tmp7174;
  wire tmp7175;
  wire tmp7176;
  wire tmp7177;
  wire tmp7178;
  wire tmp7179;
  wire tmp7180;
  wire tmp7181;
  wire tmp7182;
  wire tmp7183;
  wire tmp7184;
  wire tmp7185;
  wire tmp7186;
  wire tmp7187;
  wire tmp7188;
  wire tmp7189;
  wire tmp7190;
  wire tmp7191;
  wire tmp7192;
  wire tmp7193;
  wire tmp7194;
  wire tmp7195;
  wire tmp7196;
  wire tmp7197;
  wire tmp7198;
  wire tmp7199;
  wire tmp7200;
  wire tmp7201;
  wire tmp7202;
  wire tmp7203;
  wire tmp7204;
  wire tmp7205;
  wire tmp7206;
  wire tmp7207;
  wire tmp7208;
  wire tmp7209;
  wire tmp7210;
  wire tmp7211;
  wire tmp7212;
  wire tmp7213;
  wire tmp7214;
  wire tmp7215;
  wire tmp7216;
  wire tmp7217;
  wire tmp7218;
  wire tmp7219;
  wire tmp7220;
  wire tmp7221;
  wire tmp7222;
  wire tmp7223;
  wire tmp7224;
  wire tmp7225;
  wire tmp7226;
  wire tmp7227;
  wire tmp7228;
  wire tmp7229;
  wire tmp7230;
  wire tmp7231;
  wire tmp7232;
  wire tmp7233;
  wire tmp7234;
  wire tmp7235;
  wire tmp7236;
  wire tmp7237;
  wire tmp7238;
  wire tmp7239;
  wire tmp7240;
  wire tmp7241;
  wire tmp7242;
  wire tmp7243;
  wire tmp7244;
  wire tmp7245;
  wire tmp7246;
  wire tmp7247;
  wire tmp7248;
  wire tmp7249;
  wire tmp7250;
  wire tmp7251;
  wire tmp7252;
  wire tmp7253;
  wire tmp7254;
  wire tmp7255;
  wire tmp7256;
  wire tmp7257;
  wire tmp7258;
  wire tmp7259;
  wire tmp7260;
  wire tmp7261;
  wire tmp7262;
  wire tmp7263;
  wire tmp7264;
  wire tmp7265;
  wire tmp7266;
  wire tmp7267;
  wire tmp7268;
  wire tmp7269;
  wire tmp7270;
  wire tmp7271;
  wire tmp7272;
  wire tmp7273;
  wire tmp7274;
  wire tmp7275;
  wire tmp7276;
  wire tmp7277;
  wire tmp7278;
  wire tmp7279;
  wire tmp7280;
  wire tmp7281;
  wire tmp7282;
  wire tmp7283;
  wire tmp7284;
  wire tmp7285;
  wire tmp7286;
  wire tmp7287;
  wire tmp7288;
  wire tmp7289;
  wire tmp7290;
  wire tmp7291;
  wire tmp7292;
  wire tmp7293;
  wire tmp7294;
  wire tmp7295;
  wire tmp7296;
  wire tmp7297;
  wire tmp7298;
  wire tmp7299;
  wire tmp7300;
  wire tmp7301;
  wire tmp7302;
  wire tmp7303;
  wire tmp7304;
  wire tmp7305;
  wire tmp7306;
  wire tmp7307;
  wire tmp7308;
  wire tmp7309;
  wire tmp7310;
  wire tmp7311;
  wire tmp7312;
  wire tmp7313;
  wire tmp7314;
  wire tmp7315;
  wire tmp7316;
  wire tmp7317;
  wire tmp7318;
  wire tmp7319;
  wire tmp7320;
  wire tmp7321;
  wire tmp7322;
  wire tmp7323;
  wire tmp7324;
  wire tmp7325;
  wire tmp7326;
  wire tmp7327;
  wire tmp7328;
  wire tmp7329;
  wire tmp7330;
  wire tmp7331;
  wire tmp7332;
  wire tmp7333;
  wire tmp7334;
  wire tmp7335;
  wire tmp7336;
  wire tmp7337;
  wire tmp7338;
  wire tmp7339;
  wire tmp7340;
  wire tmp7341;
  wire tmp7342;
  wire tmp7343;
  wire tmp7344;
  wire tmp7345;
  wire tmp7346;
  wire tmp7347;
  wire tmp7348;
  wire tmp7349;
  wire tmp7350;
  wire tmp7351;
  wire tmp7352;
  wire tmp7353;
  wire tmp7354;
  wire tmp7355;
  wire tmp7356;
  wire tmp7357;
  wire tmp7358;
  wire tmp7359;
  wire tmp7360;
  wire tmp7361;
  wire tmp7362;
  wire tmp7363;
  wire tmp7364;
  wire tmp7365;
  wire tmp7366;
  wire tmp7367;
  wire tmp7368;
  wire tmp7369;
  wire tmp7370;
  wire tmp7371;
  wire tmp7372;
  wire tmp7373;
  wire tmp7374;
  wire tmp7375;
  wire tmp7376;
  wire tmp7377;
  wire tmp7378;
  wire tmp7379;
  wire tmp7380;
  wire tmp7381;
  wire tmp7382;
  wire tmp7383;
  wire tmp7384;
  wire tmp7385;
  wire tmp7386;
  wire tmp7387;
  wire tmp7388;
  wire tmp7389;
  wire tmp7390;
  wire tmp7391;
  wire tmp7392;
  wire tmp7393;
  wire tmp7394;
  wire tmp7395;
  wire tmp7396;
  wire tmp7397;
  wire tmp7398;
  wire tmp7399;
  wire tmp7400;
  wire tmp7401;
  wire tmp7402;
  wire tmp7403;
  wire tmp7404;
  wire tmp7405;
  wire tmp7406;
  wire tmp7407;
  wire tmp7408;
  wire tmp7409;
  wire tmp7410;
  wire tmp7411;
  wire tmp7412;
  wire tmp7413;
  wire tmp7414;
  wire tmp7415;
  wire tmp7416;
  wire tmp7417;
  wire tmp7418;
  wire tmp7419;
  wire tmp7420;
  wire tmp7421;
  wire tmp7422;
  wire tmp7423;
  wire tmp7424;
  wire tmp7425;
  wire tmp7426;
  wire tmp7427;
  wire tmp7428;
  wire tmp7429;
  wire tmp7430;
  wire tmp7431;
  wire tmp7432;
  wire tmp7433;
  wire tmp7434;
  wire tmp7435;
  wire tmp7436;
  wire tmp7437;
  wire tmp7438;
  wire tmp7439;
  wire tmp7440;
  wire tmp7441;
  wire tmp7442;
  wire tmp7443;
  wire tmp7444;
  wire tmp7445;
  wire tmp7446;
  wire tmp7447;
  wire tmp7448;
  wire tmp7449;
  wire tmp7450;
  wire tmp7451;
  wire tmp7452;
  wire tmp7453;
  wire tmp7454;
  wire tmp7455;
  wire tmp7456;
  wire tmp7457;
  wire tmp7458;
  wire tmp7459;
  wire tmp7460;
  wire tmp7461;
  wire tmp7462;
  wire tmp7463;
  wire tmp7464;
  wire tmp7465;
  wire tmp7466;
  wire tmp7467;
  wire tmp7468;
  wire tmp7469;
  wire tmp7470;
  wire tmp7471;
  wire tmp7472;
  wire tmp7473;
  wire tmp7474;
  wire tmp7475;
  wire tmp7476;
  wire tmp7477;
  wire tmp7478;
  wire tmp7479;
  wire tmp7480;
  wire tmp7481;
  wire tmp7482;
  wire tmp7483;
  wire tmp7484;
  wire tmp7485;
  wire tmp7486;
  wire tmp7487;
  wire tmp7488;
  wire tmp7489;
  wire tmp7490;
  wire tmp7491;
  wire tmp7492;
  wire tmp7493;
  wire tmp7494;
  wire tmp7495;
  wire tmp7496;
  wire tmp7497;
  wire tmp7498;
  wire tmp7499;
  wire tmp7500;
  wire tmp7501;
  wire tmp7502;
  wire tmp7503;
  wire tmp7504;
  wire tmp7505;
  wire tmp7506;
  wire tmp7507;
  wire tmp7508;
  wire tmp7509;
  wire tmp7510;
  wire tmp7511;
  wire tmp7512;
  wire tmp7513;
  wire tmp7514;
  wire tmp7515;
  wire tmp7516;
  wire tmp7517;
  wire tmp7518;
  wire tmp7519;
  wire tmp7520;
  wire tmp7521;
  wire tmp7522;
  wire tmp7523;
  wire tmp7524;
  wire tmp7525;
  wire tmp7526;
  wire tmp7527;
  wire tmp7528;
  wire tmp7529;
  wire tmp7530;
  wire tmp7531;
  wire tmp7532;
  wire tmp7533;
  wire tmp7534;
  wire tmp7535;
  wire tmp7536;
  wire tmp7537;
  wire tmp7538;
  wire tmp7539;
  wire tmp7540;
  wire tmp7541;
  wire tmp7542;
  wire tmp7543;
  wire tmp7544;
  wire tmp7545;
  wire tmp7546;
  wire tmp7547;
  wire tmp7548;
  wire tmp7549;
  wire tmp7550;
  wire tmp7551;
  wire tmp7552;
  wire tmp7553;
  wire tmp7554;
  wire tmp7555;
  wire tmp7556;
  wire tmp7557;
  wire tmp7558;
  wire tmp7559;
  wire tmp7560;
  wire tmp7561;
  wire tmp7562;
  wire tmp7563;
  wire tmp7564;
  wire tmp7565;
  wire tmp7566;
  wire tmp7567;
  wire tmp7568;
  wire tmp7569;
  wire tmp7570;
  wire tmp7571;
  wire tmp7572;
  wire tmp7573;
  wire tmp7574;
  wire tmp7575;
  wire tmp7576;
  wire tmp7577;
  wire tmp7578;
  wire tmp7579;
  wire tmp7580;
  wire tmp7581;
  wire tmp7582;
  wire tmp7583;
  wire tmp7584;
  wire tmp7585;
  wire tmp7586;
  wire tmp7587;
  wire tmp7588;
  wire tmp7589;
  wire tmp7590;
  wire tmp7591;
  wire tmp7592;
  wire tmp7593;
  wire tmp7594;
  wire tmp7595;
  wire tmp7596;
  wire tmp7597;
  wire tmp7598;
  wire tmp7599;
  wire tmp7600;
  wire tmp7601;
  wire tmp7602;
  wire tmp7603;
  wire tmp7604;
  wire tmp7605;
  wire tmp7606;
  wire tmp7607;
  wire tmp7608;
  wire tmp7609;
  wire tmp7610;
  wire tmp7611;
  wire tmp7612;
  wire tmp7613;
  wire tmp7614;
  wire tmp7615;
  wire tmp7616;
  wire tmp7617;
  wire tmp7618;
  wire tmp7619;
  wire tmp7620;
  wire tmp7621;
  wire tmp7622;
  wire tmp7623;
  wire tmp7624;
  wire tmp7625;
  wire tmp7626;
  wire tmp7627;
  wire tmp7628;
  wire tmp7629;
  wire tmp7630;
  wire tmp7631;
  wire tmp7632;
  wire tmp7633;
  wire tmp7634;
  wire tmp7635;
  wire tmp7636;
  wire tmp7637;
  wire tmp7638;
  wire tmp7639;
  wire tmp7640;
  wire tmp7641;
  wire tmp7642;
  wire tmp7643;
  wire tmp7644;
  wire tmp7645;
  wire tmp7646;
  wire tmp7647;
  wire tmp7648;
  wire tmp7649;
  wire tmp7650;
  wire tmp7651;
  wire tmp7652;
  wire tmp7653;
  wire tmp7654;
  wire tmp7655;
  wire tmp7656;
  wire tmp7657;
  wire tmp7658;
  wire tmp7659;
  wire tmp7660;
  wire tmp7661;
  wire tmp7662;
  wire tmp7663;
  wire tmp7664;
  wire tmp7665;
  wire tmp7666;
  wire tmp7667;
  wire tmp7668;
  wire tmp7669;
  wire tmp7670;
  wire tmp7671;
  wire tmp7672;
  wire tmp7673;
  wire tmp7674;
  wire tmp7675;
  wire tmp7676;
  wire tmp7677;
  wire tmp7678;
  wire tmp7679;
  wire tmp7680;
  wire tmp7681;
  wire tmp7682;
  wire tmp7683;
  wire tmp7684;
  wire tmp7685;
  wire tmp7686;
  wire tmp7687;
  wire tmp7688;
  wire tmp7689;
  wire tmp7690;
  wire tmp7691;
  wire tmp7692;
  wire tmp7693;
  wire tmp7694;
  wire tmp7695;
  wire tmp7696;
  wire tmp7697;
  wire tmp7698;
  wire tmp7699;
  wire tmp7700;
  wire tmp7701;
  wire tmp7702;
  wire tmp7703;
  wire tmp7704;
  wire tmp7705;
  wire tmp7706;
  wire tmp7707;
  wire tmp7708;
  wire tmp7709;
  wire tmp7710;
  wire tmp7711;
  wire tmp7712;
  wire tmp7713;
  wire tmp7714;
  wire tmp7715;
  wire tmp7716;
  wire tmp7717;
  wire tmp7718;
  wire tmp7719;
  wire tmp7720;
  wire tmp7721;
  wire tmp7722;
  wire tmp7723;
  wire tmp7724;
  wire tmp7725;
  wire tmp7726;
  wire tmp7727;
  wire tmp7728;
  wire tmp7729;
  wire tmp7730;
  wire tmp7731;
  wire tmp7732;
  wire tmp7733;
  wire tmp7734;
  wire tmp7735;
  wire tmp7736;
  wire tmp7737;
  wire tmp7738;
  wire tmp7739;
  wire tmp7740;
  wire tmp7741;
  wire tmp7742;
  wire tmp7743;
  wire tmp7744;
  wire tmp7745;
  wire tmp7746;
  wire tmp7747;
  wire tmp7748;
  wire tmp7749;
  wire tmp7750;
  wire tmp7751;
  wire tmp7752;
  wire tmp7753;
  wire tmp7754;
  wire tmp7755;
  wire tmp7756;
  wire tmp7757;
  wire tmp7758;
  wire tmp7759;
  wire tmp7760;
  wire tmp7761;
  wire tmp7762;
  wire tmp7763;
  wire tmp7764;
  wire tmp7765;
  wire tmp7766;
  wire tmp7767;
  wire tmp7768;
  wire tmp7769;
  wire tmp7770;
  wire tmp7771;
  wire tmp7772;
  wire tmp7773;
  wire tmp7774;
  wire tmp7775;
  wire tmp7776;
  wire tmp7777;
  wire tmp7778;
  wire tmp7779;
  wire tmp7780;
  wire tmp7781;
  wire tmp7782;
  wire tmp7783;
  wire tmp7784;
  wire tmp7785;
  wire tmp7786;
  wire tmp7787;
  wire tmp7788;
  wire tmp7789;
  wire tmp7790;
  wire tmp7791;
  wire tmp7792;
  wire tmp7793;
  wire tmp7794;
  wire tmp7795;
  wire tmp7796;
  wire tmp7797;
  wire tmp7798;
  wire tmp7799;
  wire tmp7800;
  wire tmp7801;
  wire tmp7802;
  wire tmp7803;
  wire tmp7804;
  wire tmp7805;
  wire tmp7806;
  wire tmp7807;
  wire tmp7808;
  wire tmp7809;
  wire tmp7810;
  wire tmp7811;
  wire tmp7812;
  wire tmp7813;
  wire tmp7814;
  wire tmp7815;
  wire tmp7816;
  wire tmp7817;
  wire tmp7818;
  wire tmp7819;
  wire tmp7820;
  wire tmp7821;
  wire tmp7822;
  wire tmp7823;
  wire tmp7824;
  wire tmp7825;
  wire tmp7826;
  wire tmp7827;
  wire tmp7828;
  wire tmp7829;
  wire tmp7830;
  wire tmp7831;
  wire tmp7832;
  wire tmp7833;
  wire tmp7834;
  wire tmp7835;
  wire tmp7836;
  wire tmp7837;
  wire tmp7838;
  wire tmp7839;
  wire tmp7840;
  wire tmp7841;
  wire tmp7842;
  wire tmp7843;
  wire tmp7844;
  wire tmp7845;
  wire tmp7846;
  wire tmp7847;
  wire tmp7848;
  wire tmp7849;
  wire tmp7850;
  wire tmp7851;
  wire tmp7852;
  wire tmp7853;
  wire tmp7854;
  wire tmp7855;
  wire tmp7856;
  wire tmp7857;
  wire tmp7858;
  wire tmp7859;
  wire tmp7860;
  wire tmp7861;
  wire tmp7862;
  wire tmp7863;
  wire tmp7864;
  wire tmp7865;
  wire tmp7866;
  wire tmp7867;
  wire tmp7868;
  wire tmp7869;
  wire tmp7870;
  wire tmp7871;
  wire tmp7872;
  wire tmp7873;
  wire tmp7874;
  wire tmp7875;
  wire tmp7876;
  wire tmp7877;
  wire tmp7878;
  wire tmp7879;
  wire tmp7880;
  wire tmp7881;
  wire tmp7882;
  wire tmp7883;
  wire tmp7884;
  wire tmp7885;
  wire tmp7886;
  wire tmp7887;
  wire tmp7888;
  wire tmp7889;
  wire tmp7890;
  wire tmp7891;
  wire tmp7892;
  wire tmp7893;
  wire tmp7894;
  wire tmp7895;
  wire tmp7896;
  wire tmp7897;
  wire tmp7898;
  wire tmp7899;
  wire tmp7900;
  wire tmp7901;
  wire tmp7902;
  wire tmp7903;
  wire tmp7904;
  wire tmp7905;
  wire tmp7906;
  wire tmp7907;
  wire tmp7908;
  wire tmp7909;
  wire tmp7910;
  wire tmp7911;
  wire tmp7912;
  wire tmp7913;
  wire tmp7914;
  wire tmp7915;
  wire tmp7916;
  wire tmp7917;
  wire tmp7918;
  wire tmp7919;
  wire tmp7920;
  wire tmp7921;
  wire tmp7922;
  wire tmp7923;
  wire tmp7924;
  wire tmp7925;
  wire tmp7926;
  wire tmp7927;
  wire tmp7928;
  wire tmp7929;
  wire tmp7930;
  wire tmp7931;
  wire tmp7932;
  wire tmp7933;
  wire tmp7934;
  wire tmp7935;
  wire tmp7936;
  wire tmp7937;
  wire tmp7938;
  wire tmp7939;
  wire tmp7940;
  wire tmp7941;
  wire tmp7942;
  wire tmp7943;
  wire tmp7944;
  wire tmp7945;
  wire tmp7946;
  wire tmp7947;
  wire tmp7948;
  wire tmp7949;
  wire tmp7950;
  wire tmp7951;
  wire tmp7952;
  wire tmp7953;
  wire tmp7954;
  wire tmp7955;
  wire tmp7956;
  wire tmp7957;
  wire tmp7958;
  wire tmp7959;
  wire tmp7960;
  wire tmp7961;
  wire tmp7962;
  wire tmp7963;
  wire tmp7964;
  wire tmp7965;
  wire tmp7966;
  wire tmp7967;
  wire tmp7968;
  wire tmp7969;
  wire tmp7970;
  wire tmp7971;
  wire tmp7972;
  wire tmp7973;
  wire tmp7974;
  wire tmp7975;
  wire tmp7976;
  wire tmp7977;
  wire tmp7978;
  wire tmp7979;
  wire tmp7980;
  wire tmp7981;
  wire tmp7982;
  wire tmp7983;
  wire tmp7984;
  wire tmp7985;
  wire tmp7986;
  wire tmp7987;
  wire tmp7988;
  wire tmp7989;
  wire tmp7990;
  wire tmp7991;
  wire tmp7992;
  wire tmp7993;
  wire tmp7994;
  wire tmp7995;
  wire tmp7996;
  wire tmp7997;
  wire tmp7998;
  wire tmp7999;
  wire tmp8000;
  wire tmp8001;
  wire tmp8002;
  wire tmp8003;
  wire tmp8004;
  wire tmp8005;
  wire tmp8006;
  wire tmp8007;
  wire tmp8008;
  wire tmp8009;
  wire tmp8010;
  wire tmp8011;
  wire tmp8012;
  wire tmp8013;
  wire tmp8014;
  wire tmp8015;
  wire tmp8016;
  wire tmp8017;
  wire tmp8018;
  wire tmp8019;
  wire tmp8020;
  wire tmp8021;
  wire tmp8022;
  wire tmp8023;
  wire tmp8024;
  wire tmp8025;
  wire tmp8026;
  wire tmp8027;
  wire tmp8028;
  wire tmp8029;
  wire tmp8030;
  wire tmp8031;
  wire tmp8032;
  wire tmp8033;
  wire tmp8034;
  wire tmp8035;
  wire tmp8036;
  wire tmp8037;
  wire tmp8038;
  wire tmp8039;
  wire tmp8040;
  wire tmp8041;
  wire tmp8042;
  wire tmp8043;
  wire tmp8044;
  wire tmp8045;
  wire tmp8046;
  wire tmp8047;
  wire tmp8048;
  wire tmp8049;
  wire tmp8050;
  wire tmp8051;
  wire tmp8052;
  wire tmp8053;
  wire tmp8054;
  wire tmp8055;
  wire tmp8056;
  wire tmp8057;
  wire tmp8058;
  wire tmp8059;
  wire tmp8060;
  wire tmp8061;
  wire tmp8062;
  wire tmp8063;
  wire tmp8064;
  wire tmp8065;
  wire tmp8066;
  wire tmp8067;
  wire tmp8068;
  wire tmp8069;
  wire tmp8070;
  wire tmp8071;
  wire tmp8072;
  wire tmp8073;
  wire tmp8074;
  wire tmp8075;
  wire tmp8076;
  wire tmp8077;
  wire tmp8078;
  wire tmp8079;
  wire tmp8080;
  wire tmp8081;
  wire tmp8082;
  wire tmp8083;
  wire tmp8084;
  wire tmp8085;
  wire tmp8086;
  wire tmp8087;
  wire tmp8088;
  wire tmp8089;
  wire tmp8090;
  wire tmp8091;
  wire tmp8092;
  wire tmp8093;
  wire tmp8094;
  wire tmp8095;
  wire tmp8096;
  wire tmp8097;
  wire tmp8098;
  wire tmp8099;
  wire tmp8100;
  wire tmp8101;
  wire tmp8102;
  wire tmp8103;
  wire tmp8104;
  wire tmp8105;
  wire tmp8106;
  wire tmp8107;
  wire tmp8108;
  wire tmp8109;
  wire tmp8110;
  wire tmp8111;
  wire tmp8112;
  wire tmp8113;
  wire tmp8114;
  wire tmp8115;
  wire tmp8116;
  wire tmp8117;
  wire tmp8118;
  wire tmp8119;
  wire tmp8120;
  wire tmp8121;
  wire tmp8122;
  wire tmp8123;
  wire tmp8124;
  wire tmp8125;
  wire tmp8126;
  wire tmp8127;
  wire tmp8128;
  wire tmp8129;
  wire tmp8130;
  wire tmp8131;
  wire tmp8132;
  wire tmp8133;
  wire tmp8134;
  wire tmp8135;
  wire tmp8136;
  wire tmp8137;
  wire tmp8138;
  wire tmp8139;
  wire tmp8140;
  wire tmp8141;
  wire tmp8142;
  wire tmp8143;
  wire tmp8144;
  wire tmp8145;
  wire tmp8146;
  wire tmp8147;
  wire tmp8148;
  wire tmp8149;
  wire tmp8150;
  wire tmp8151;
  wire tmp8152;
  wire tmp8153;
  wire tmp8154;
  wire tmp8155;
  wire tmp8156;
  wire tmp8157;
  wire tmp8158;
  wire tmp8159;
  wire tmp8160;
  wire tmp8161;
  wire tmp8162;
  wire tmp8163;
  wire tmp8164;
  wire tmp8165;
  wire tmp8166;
  wire tmp8167;
  wire tmp8168;
  wire tmp8169;
  wire tmp8170;
  wire tmp8171;
  wire tmp8172;
  wire tmp8173;
  wire tmp8174;
  wire tmp8175;
  wire tmp8176;
  wire tmp8177;
  wire tmp8178;
  wire tmp8179;
  wire tmp8180;
  wire tmp8181;
  wire tmp8182;
  wire tmp8183;
  wire tmp8184;
  wire tmp8185;
  wire tmp8186;
  wire tmp8187;
  wire tmp8188;
  wire tmp8189;
  wire tmp8190;
  wire tmp8191;
  wire tmp8192;
  wire tmp8193;
  wire tmp8194;
  wire tmp8195;
  wire tmp8196;
  wire tmp8197;
  wire tmp8198;
  wire tmp8199;
  wire tmp8200;
  wire tmp8201;
  wire tmp8202;
  wire tmp8203;
  wire tmp8204;
  wire tmp8205;
  wire tmp8206;
  wire tmp8207;
  wire tmp8208;
  wire tmp8209;
  wire tmp8210;
  wire tmp8211;
  wire tmp8212;
  wire tmp8213;
  wire tmp8214;
  wire tmp8215;
  wire tmp8216;
  wire tmp8217;
  wire tmp8218;
  wire tmp8219;
  wire tmp8220;
  wire tmp8221;
  wire tmp8222;
  wire tmp8223;
  wire tmp8224;
  wire tmp8225;
  wire tmp8226;
  wire tmp8227;
  wire tmp8228;
  wire tmp8229;
  wire tmp8230;
  wire tmp8231;
  wire tmp8232;
  wire tmp8233;
  wire tmp8234;
  wire tmp8235;
  wire tmp8236;
  wire tmp8237;
  wire tmp8238;
  wire tmp8239;
  wire tmp8240;
  wire tmp8241;
  wire tmp8242;
  wire tmp8243;
  wire tmp8244;
  wire tmp8245;
  wire tmp8246;
  wire tmp8247;
  wire tmp8248;
  wire tmp8249;
  wire tmp8250;
  wire tmp8251;
  wire tmp8252;
  wire tmp8253;
  wire tmp8254;
  wire tmp8255;
  wire tmp8256;
  wire tmp8257;
  wire tmp8258;
  wire tmp8259;
  wire tmp8260;
  wire tmp8261;
  wire tmp8262;
  wire tmp8263;
  wire tmp8264;
  wire tmp8265;
  wire tmp8266;
  wire tmp8267;
  wire tmp8268;
  wire tmp8269;
  wire tmp8270;
  wire tmp8271;
  wire tmp8272;
  wire tmp8273;
  wire tmp8274;
  wire tmp8275;
  wire tmp8276;
  wire tmp8277;
  wire tmp8278;
  wire tmp8279;
  wire tmp8280;
  wire tmp8281;
  wire tmp8282;
  wire tmp8283;
  wire tmp8284;
  wire tmp8285;
  wire tmp8286;
  wire tmp8287;
  wire tmp8288;
  wire tmp8289;
  wire tmp8290;
  wire tmp8291;
  wire tmp8292;
  wire tmp8293;
  wire tmp8294;
  wire tmp8295;
  wire tmp8296;
  wire tmp8297;
  wire tmp8298;
  wire tmp8299;
  wire tmp8300;
  wire tmp8301;
  wire tmp8302;
  wire tmp8303;
  wire tmp8304;
  wire tmp8305;
  wire tmp8306;
  wire tmp8307;
  wire tmp8308;
  wire tmp8309;
  wire tmp8310;
  wire tmp8311;
  wire tmp8312;
  wire tmp8313;
  wire tmp8314;
  wire tmp8315;
  wire tmp8316;
  wire tmp8317;
  wire tmp8318;
  wire tmp8319;
  wire tmp8320;
  wire tmp8321;
  wire tmp8322;
  wire tmp8323;
  wire tmp8324;
  wire tmp8325;
  wire tmp8326;
  wire tmp8327;
  wire tmp8328;
  wire tmp8329;
  wire tmp8330;
  wire tmp8331;
  wire tmp8332;
  wire tmp8333;
  wire tmp8334;
  wire tmp8335;
  wire tmp8336;
  wire tmp8337;
  wire tmp8338;
  wire tmp8339;
  wire tmp8340;
  wire tmp8341;
  wire tmp8342;
  wire tmp8343;
  wire tmp8344;
  wire tmp8345;
  wire tmp8346;
  wire tmp8347;
  wire tmp8348;
  wire tmp8349;
  wire tmp8350;
  wire tmp8351;
  wire tmp8352;
  wire tmp8353;
  wire tmp8354;
  wire tmp8355;
  wire tmp8356;
  wire tmp8357;
  wire tmp8358;
  wire tmp8359;
  wire tmp8360;
  wire tmp8361;
  wire tmp8362;
  wire tmp8363;
  wire tmp8364;
  wire tmp8365;
  wire tmp8366;
  wire tmp8367;
  wire tmp8368;
  wire tmp8369;
  wire tmp8370;
  wire tmp8371;
  wire tmp8372;
  wire tmp8373;
  wire tmp8374;
  wire tmp8375;
  wire tmp8376;
  wire tmp8377;
  wire tmp8378;
  wire tmp8379;
  wire tmp8380;
  wire tmp8381;
  wire tmp8382;
  wire tmp8383;
  wire tmp8384;
  wire tmp8385;
  wire tmp8386;
  wire tmp8387;
  wire tmp8388;
  wire tmp8389;
  wire tmp8390;
  wire tmp8391;
  wire tmp8392;
  wire tmp8393;
  wire tmp8394;
  wire tmp8395;
  wire tmp8396;
  wire tmp8397;
  wire tmp8398;
  wire tmp8399;
  wire tmp8400;
  wire tmp8401;
  wire tmp8402;
  wire tmp8403;
  wire tmp8404;
  wire tmp8405;
  wire tmp8406;
  wire tmp8407;
  wire tmp8408;
  wire tmp8409;
  wire tmp8410;
  wire tmp8411;
  wire tmp8412;
  wire tmp8413;
  wire tmp8414;
  wire tmp8415;
  wire tmp8416;
  wire tmp8417;
  wire tmp8418;
  wire tmp8419;
  wire tmp8420;
  wire tmp8421;
  wire tmp8422;
  wire tmp8423;
  wire tmp8424;
  wire tmp8425;
  wire tmp8426;
  wire tmp8427;
  wire tmp8428;
  wire tmp8429;
  wire tmp8430;
  wire tmp8431;
  wire tmp8432;
  wire tmp8433;
  wire tmp8434;
  wire tmp8435;
  wire tmp8436;
  wire tmp8437;
  wire tmp8438;
  wire tmp8439;
  wire tmp8440;
  wire tmp8441;
  wire tmp8442;
  wire tmp8443;
  wire tmp8444;
  wire tmp8445;
  wire tmp8446;
  wire tmp8447;
  wire tmp8448;
  wire tmp8449;
  wire tmp8450;
  wire tmp8451;
  wire tmp8452;
  wire tmp8453;
  wire tmp8454;
  wire tmp8455;
  wire tmp8456;
  wire tmp8457;
  wire tmp8458;
  wire tmp8459;
  wire tmp8460;
  wire tmp8461;
  wire tmp8462;
  wire tmp8463;
  wire tmp8464;
  wire tmp8465;
  wire tmp8466;
  wire tmp8467;
  wire tmp8468;
  wire tmp8469;
  wire tmp8470;
  wire tmp8471;
  wire tmp8472;
  wire tmp8473;
  wire tmp8474;
  wire tmp8475;
  wire tmp8476;
  wire tmp8477;
  wire tmp8478;
  wire tmp8479;
  wire tmp8480;
  wire tmp8481;
  wire tmp8482;
  wire tmp8483;
  wire tmp8484;
  wire tmp8485;
  wire tmp8486;
  wire tmp8487;
  wire tmp8488;
  wire tmp8489;
  wire tmp8490;
  wire tmp8491;
  wire tmp8492;
  wire tmp8493;
  wire tmp8494;
  wire tmp8495;
  wire tmp8496;
  wire tmp8497;
  wire tmp8498;
  wire tmp8499;
  wire tmp8500;
  wire tmp8501;
  wire tmp8502;
  wire tmp8503;
  wire tmp8504;
  wire tmp8505;
  wire tmp8506;
  wire tmp8507;
  wire tmp8508;
  wire tmp8509;
  wire tmp8510;
  wire tmp8511;
  wire tmp8512;
  wire tmp8513;
  wire tmp8514;
  wire tmp8515;
  wire tmp8516;
  wire tmp8517;
  wire tmp8518;
  wire tmp8519;
  wire tmp8520;
  wire tmp8521;
  wire tmp8522;
  wire tmp8523;
  wire tmp8524;
  wire tmp8525;
  wire tmp8526;
  wire tmp8527;
  wire tmp8528;
  wire tmp8529;
  wire tmp8530;
  wire tmp8531;
  wire tmp8532;
  wire tmp8533;
  wire tmp8534;
  wire tmp8535;
  wire tmp8536;
  wire tmp8537;
  wire tmp8538;
  wire tmp8539;
  wire tmp8540;
  wire tmp8541;
  wire tmp8542;
  wire tmp8543;
  wire tmp8544;
  wire tmp8545;
  wire tmp8546;
  wire tmp8547;
  wire tmp8548;
  wire tmp8549;
  wire tmp8550;
  wire tmp8551;
  wire tmp8552;
  wire tmp8553;
  wire tmp8554;
  wire tmp8555;
  wire tmp8556;
  wire tmp8557;
  wire tmp8558;
  wire tmp8559;
  wire tmp8560;
  wire tmp8561;
  wire tmp8562;
  wire tmp8563;
  wire tmp8564;
  wire tmp8565;
  wire tmp8566;
  wire tmp8567;
  wire tmp8568;
  wire tmp8569;
  wire tmp8570;
  wire tmp8571;
  wire tmp8572;
  wire tmp8573;
  wire tmp8574;
  wire tmp8575;
  wire tmp8576;
  wire tmp8577;
  wire tmp8578;
  wire tmp8579;
  wire tmp8580;
  wire tmp8581;
  wire tmp8582;
  wire tmp8583;
  wire tmp8584;
  wire tmp8585;
  wire tmp8586;
  wire tmp8587;
  wire tmp8588;
  wire tmp8589;
  wire tmp8590;
  wire tmp8591;
  wire tmp8592;
  wire tmp8593;
  wire tmp8594;
  wire tmp8595;
  wire tmp8596;
  wire tmp8597;
  wire tmp8598;
  wire tmp8599;
  wire tmp8600;
  wire tmp8601;
  wire tmp8602;
  wire tmp8603;
  wire tmp8604;
  wire tmp8605;
  wire tmp8606;
  wire tmp8607;
  wire tmp8608;
  wire tmp8609;
  wire tmp8610;
  wire tmp8611;
  wire tmp8612;
  wire tmp8613;
  wire tmp8614;
  wire tmp8615;
  wire tmp8616;
  wire tmp8617;
  wire tmp8618;
  wire tmp8619;
  wire tmp8620;
  wire tmp8621;
  wire tmp8622;
  wire tmp8623;
  wire tmp8624;
  wire tmp8625;
  wire tmp8626;
  wire tmp8627;
  wire tmp8628;
  wire tmp8629;
  wire tmp8630;
  wire tmp8631;
  wire tmp8632;
  wire tmp8633;
  wire tmp8634;
  wire tmp8635;
  wire tmp8636;
  wire tmp8637;
  wire tmp8638;
  wire tmp8639;
  wire tmp8640;
  wire tmp8641;
  wire tmp8642;
  wire tmp8643;
  wire tmp8644;
  wire tmp8645;
  wire tmp8646;
  wire tmp8647;
  wire tmp8648;
  wire tmp8649;
  wire tmp8650;
  wire tmp8651;
  wire tmp8652;
  wire tmp8653;
  wire tmp8654;
  wire tmp8655;
  wire tmp8656;
  wire tmp8657;
  wire tmp8658;
  wire tmp8659;
  wire tmp8660;
  wire tmp8661;
  wire tmp8662;
  wire tmp8663;
  wire tmp8664;
  wire tmp8665;
  wire tmp8666;
  wire tmp8667;
  wire tmp8668;
  wire tmp8669;
  wire tmp8670;
  wire tmp8671;
  wire tmp8672;
  wire tmp8673;
  wire tmp8674;
  wire tmp8675;
  wire tmp8676;
  wire tmp8677;
  wire tmp8678;
  wire tmp8679;
  wire tmp8680;
  wire tmp8681;
  wire tmp8682;
  wire tmp8683;
  wire tmp8684;
  wire tmp8685;
  wire tmp8686;
  wire tmp8687;
  wire tmp8688;
  wire tmp8689;
  wire tmp8690;
  wire tmp8691;
  wire tmp8692;
  wire tmp8693;
  wire tmp8694;
  wire tmp8695;
  wire tmp8696;
  wire tmp8697;
  wire tmp8698;
  wire tmp8699;
  wire tmp8700;
  wire tmp8701;
  wire tmp8702;
  wire tmp8703;
  wire tmp8704;
  wire tmp8705;
  wire tmp8706;
  wire tmp8707;
  wire tmp8708;
  wire tmp8709;
  wire tmp8710;
  wire tmp8711;
  wire tmp8712;
  wire tmp8713;
  wire tmp8714;
  wire tmp8715;
  wire tmp8716;
  wire tmp8717;
  wire tmp8718;
  wire tmp8719;
  wire tmp8720;
  wire tmp8721;
  wire tmp8722;
  wire tmp8723;
  wire tmp8724;
  wire tmp8725;
  wire tmp8726;
  wire tmp8727;
  wire tmp8728;
  wire tmp8729;
  wire tmp8730;
  wire tmp8731;
  wire tmp8732;
  wire tmp8733;
  wire tmp8734;
  wire tmp8735;
  wire tmp8736;
  wire tmp8737;
  wire tmp8738;
  wire tmp8739;
  wire tmp8740;
  wire tmp8741;
  wire tmp8742;
  wire tmp8743;
  wire tmp8744;
  wire tmp8745;
  wire tmp8746;
  wire tmp8747;
  wire tmp8748;
  wire tmp8749;
  wire tmp8750;
  wire tmp8751;
  wire tmp8752;
  wire tmp8753;
  wire tmp8754;
  wire tmp8755;
  wire tmp8756;
  wire tmp8757;
  wire tmp8758;
  wire tmp8759;
  wire tmp8760;
  wire tmp8761;
  wire tmp8762;
  wire tmp8763;
  wire tmp8764;
  wire tmp8765;
  wire tmp8766;
  wire tmp8767;
  wire tmp8768;
  wire tmp8769;
  wire tmp8770;
  wire tmp8771;
  wire tmp8772;
  wire tmp8773;
  wire tmp8774;
  wire tmp8775;
  wire tmp8776;
  wire tmp8777;
  wire tmp8778;
  wire tmp8779;
  wire tmp8780;
  wire tmp8781;
  wire tmp8782;
  wire tmp8783;
  wire tmp8784;
  wire tmp8785;
  wire tmp8786;
  wire tmp8787;
  wire tmp8788;
  wire tmp8789;
  wire tmp8790;
  wire tmp8791;
  wire tmp8792;
  wire tmp8793;
  wire tmp8794;
  wire tmp8795;
  wire tmp8796;
  wire tmp8797;
  wire tmp8798;
  wire tmp8799;
  wire tmp8800;
  wire tmp8801;
  wire tmp8802;
  wire tmp8803;
  wire tmp8804;
  wire tmp8805;
  wire tmp8806;
  wire tmp8807;
  wire tmp8808;
  wire tmp8809;
  wire tmp8810;
  wire tmp8811;
  wire tmp8812;
  wire tmp8813;
  wire tmp8814;
  wire tmp8815;
  wire tmp8816;
  wire tmp8817;
  wire tmp8818;
  wire tmp8819;
  wire tmp8820;
  wire tmp8821;
  wire tmp8822;
  wire tmp8823;
  wire tmp8824;
  wire tmp8825;
  wire tmp8826;
  wire tmp8827;
  wire tmp8828;
  wire tmp8829;
  wire tmp8830;
  wire tmp8831;
  wire tmp8832;
  wire tmp8833;
  wire tmp8834;
  wire tmp8835;
  wire tmp8836;
  wire tmp8837;
  wire tmp8838;
  wire tmp8839;
  wire tmp8840;
  wire tmp8841;
  wire tmp8842;
  wire tmp8843;
  wire tmp8844;
  wire tmp8845;
  wire tmp8846;
  wire tmp8847;
  wire tmp8848;
  wire tmp8849;
  wire tmp8850;
  wire tmp8851;
  wire tmp8852;
  wire tmp8853;
  wire tmp8854;
  wire tmp8855;
  wire tmp8856;
  wire tmp8857;
  wire tmp8858;
  wire tmp8859;
  wire tmp8860;
  wire tmp8861;
  wire tmp8862;
  wire tmp8863;
  wire tmp8864;
  wire tmp8865;
  wire tmp8866;
  wire tmp8867;
  wire tmp8868;
  wire tmp8869;
  wire tmp8870;
  wire tmp8871;
  wire tmp8872;
  wire tmp8873;
  wire tmp8874;
  wire tmp8875;
  wire tmp8876;
  wire tmp8877;
  wire tmp8878;
  wire tmp8879;
  wire tmp8880;
  wire tmp8881;
  wire tmp8882;
  wire tmp8883;
  wire tmp8884;
  wire tmp8885;
  wire tmp8886;
  wire tmp8887;
  wire tmp8888;
  wire tmp8889;
  wire tmp8890;
  wire tmp8891;
  wire tmp8892;
  wire tmp8893;
  wire tmp8894;
  wire tmp8895;
  wire tmp8896;
  wire tmp8897;
  wire tmp8898;
  wire tmp8899;
  wire tmp8900;
  wire tmp8901;
  wire tmp8902;
  wire tmp8903;
  wire tmp8904;
  wire tmp8905;
  wire tmp8906;
  wire tmp8907;
  wire tmp8908;
  wire tmp8909;
  wire tmp8910;
  wire tmp8911;
  wire tmp8912;
  wire tmp8913;
  wire tmp8914;
  wire tmp8915;
  wire tmp8916;
  wire tmp8917;
  wire tmp8918;
  wire tmp8919;
  wire tmp8920;
  wire tmp8921;
  wire tmp8922;
  wire tmp8923;
  wire tmp8924;
  wire tmp8925;
  wire tmp8926;
  wire tmp8927;
  wire tmp8928;
  wire tmp8929;
  wire tmp8930;
  wire tmp8931;
  wire tmp8932;
  wire tmp8933;
  wire tmp8934;
  wire tmp8935;
  wire tmp8936;
  wire tmp8937;
  wire tmp8938;
  wire tmp8939;
  wire tmp8940;
  wire tmp8941;
  wire tmp8942;
  wire tmp8943;
  wire tmp8944;
  wire tmp8945;
  wire tmp8946;
  wire tmp8947;
  wire tmp8948;
  wire tmp8949;
  wire tmp8950;
  wire tmp8951;
  wire tmp8952;
  wire tmp8953;
  wire tmp8954;
  wire tmp8955;
  wire tmp8956;
  wire tmp8957;
  wire tmp8958;
  wire tmp8959;
  wire tmp8960;
  wire tmp8961;
  wire tmp8962;
  wire tmp8963;
  wire tmp8964;
  wire tmp8965;
  wire tmp8966;
  wire tmp8967;
  wire tmp8968;
  wire tmp8969;
  wire tmp8970;
  wire tmp8971;
  wire tmp8972;
  wire tmp8973;
  wire tmp8974;
  wire tmp8975;
  wire tmp8976;
  wire tmp8977;
  wire tmp8978;
  wire tmp8979;
  wire tmp8980;
  wire tmp8981;
  wire tmp8982;
  wire tmp8983;
  wire tmp8984;
  wire tmp8985;
  wire tmp8986;
  wire tmp8987;
  wire tmp8988;
  wire tmp8989;
  wire tmp8990;
  wire tmp8991;
  wire tmp8992;
  wire tmp8993;
  wire tmp8994;
  wire tmp8995;
  wire tmp8996;
  wire tmp8997;
  wire tmp8998;
  wire tmp8999;
  wire tmp9000;
  wire tmp9001;
  wire tmp9002;
  wire tmp9003;
  wire tmp9004;
  wire tmp9005;
  wire tmp9006;
  wire tmp9007;
  wire tmp9008;
  wire tmp9009;
  wire tmp9010;
  wire tmp9011;
  wire tmp9012;
  wire tmp9013;
  wire tmp9014;
  wire tmp9015;
  wire tmp9016;
  wire tmp9017;
  wire tmp9018;
  wire tmp9019;
  wire tmp9020;
  wire tmp9021;
  wire tmp9022;
  wire tmp9023;
  wire tmp9024;
  wire tmp9025;
  wire tmp9026;
  wire tmp9027;
  wire tmp9028;
  wire tmp9029;
  wire tmp9030;
  wire tmp9031;
  wire tmp9032;
  wire tmp9033;
  wire tmp9034;
  wire tmp9035;
  wire tmp9036;
  wire tmp9037;
  wire tmp9038;
  wire tmp9039;
  wire tmp9040;
  wire tmp9041;
  wire tmp9042;
  wire tmp9043;
  wire tmp9044;
  wire tmp9045;
  wire tmp9046;
  wire tmp9047;
  wire tmp9048;
  wire tmp9049;
  wire tmp9050;
  wire tmp9051;
  wire tmp9052;
  wire tmp9053;
  wire tmp9054;
  wire tmp9055;
  wire tmp9056;
  wire tmp9057;
  wire tmp9058;
  wire tmp9059;
  wire tmp9060;
  wire tmp9061;
  wire tmp9062;
  wire tmp9063;
  wire tmp9064;
  wire tmp9065;
  wire tmp9066;
  wire tmp9067;
  wire tmp9068;
  wire tmp9069;
  wire tmp9070;
  wire tmp9071;
  wire tmp9072;
  wire tmp9073;
  wire tmp9074;
  wire tmp9075;
  wire tmp9076;
  wire tmp9077;
  wire tmp9078;
  wire tmp9079;
  wire tmp9080;
  wire tmp9081;
  wire tmp9082;
  wire tmp9083;
  wire tmp9084;
  wire tmp9085;
  wire tmp9086;
  wire tmp9087;
  wire tmp9088;
  wire tmp9089;
  wire tmp9090;
  wire tmp9091;
  wire tmp9092;
  wire tmp9093;
  wire tmp9094;
  wire tmp9095;
  wire tmp9096;
  wire tmp9097;
  wire tmp9098;
  wire tmp9099;
  wire tmp9100;
  wire tmp9101;
  wire tmp9102;
  wire tmp9103;
  wire tmp9104;
  wire tmp9105;
  wire tmp9106;
  wire tmp9107;
  wire tmp9108;
  wire tmp9109;
  wire tmp9110;
  wire tmp9111;
  wire tmp9112;
  wire tmp9113;
  wire tmp9114;
  wire tmp9115;
  wire tmp9116;
  wire tmp9117;
  wire tmp9118;
  wire tmp9119;
  wire tmp9120;
  wire tmp9121;
  wire tmp9122;
  wire tmp9123;
  wire tmp9124;
  wire tmp9125;
  wire tmp9126;
  wire tmp9127;
  wire tmp9128;
  wire tmp9129;
  wire tmp9130;
  wire tmp9131;
  wire tmp9132;
  wire tmp9133;
  wire tmp9134;
  wire tmp9135;
  wire tmp9136;
  wire tmp9137;
  wire tmp9138;
  wire tmp9139;
  wire tmp9140;
  wire tmp9141;
  wire tmp9142;
  wire tmp9143;
  wire tmp9144;
  wire tmp9145;
  wire tmp9146;
  wire tmp9147;
  wire tmp9148;
  wire tmp9149;
  wire tmp9150;
  wire tmp9151;
  wire tmp9152;
  wire tmp9153;
  wire tmp9154;
  wire tmp9155;
  wire tmp9156;
  wire tmp9157;
  wire tmp9158;
  wire tmp9159;
  wire tmp9160;
  wire tmp9161;
  wire tmp9162;
  wire tmp9163;
  wire tmp9164;
  wire tmp9165;
  wire tmp9166;
  wire tmp9167;
  wire tmp9168;
  wire tmp9169;
  wire tmp9170;
  wire tmp9171;
  wire tmp9172;
  wire tmp9173;
  wire tmp9174;
  wire tmp9175;
  wire tmp9176;
  wire tmp9177;
  wire tmp9178;
  wire tmp9179;
  wire tmp9180;
  wire tmp9181;
  wire tmp9182;
  wire tmp9183;
  wire tmp9184;
  wire tmp9185;
  wire tmp9186;
  wire tmp9187;
  wire tmp9188;
  wire tmp9189;
  wire tmp9190;
  wire tmp9191;
  wire tmp9192;
  wire tmp9193;
  wire tmp9194;
  wire tmp9195;
  wire tmp9196;
  wire tmp9197;
  wire tmp9198;
  wire tmp9199;
  wire tmp9200;
  wire tmp9201;
  wire tmp9202;
  wire tmp9203;
  wire tmp9204;
  wire tmp9205;
  wire tmp9206;
  wire tmp9207;
  wire tmp9208;
  wire tmp9209;
  wire tmp9210;
  wire tmp9211;
  wire tmp9212;
  wire tmp9213;
  wire tmp9214;
  wire tmp9215;
  wire tmp9216;
  wire tmp9217;
  wire tmp9218;
  wire tmp9219;
  wire tmp9220;
  wire tmp9221;
  wire tmp9222;
  wire tmp9223;
  wire tmp9224;
  wire tmp9225;
  wire tmp9226;
  wire tmp9227;
  wire tmp9228;
  wire tmp9229;
  wire tmp9230;
  wire tmp9231;
  wire tmp9232;
  wire tmp9233;
  wire tmp9234;
  wire tmp9235;
  wire tmp9236;
  wire tmp9237;
  wire tmp9238;
  wire tmp9239;
  wire tmp9240;
  wire tmp9241;
  wire tmp9242;
  wire tmp9243;
  wire tmp9244;
  wire tmp9245;
  wire tmp9246;
  wire tmp9247;
  wire tmp9248;
  wire tmp9249;
  wire tmp9250;
  wire tmp9251;
  wire tmp9252;
  wire tmp9253;
  wire tmp9254;
  wire tmp9255;
  wire tmp9256;
  wire tmp9257;
  wire tmp9258;
  wire tmp9259;
  wire tmp9260;
  wire tmp9261;
  wire tmp9262;
  wire tmp9263;
  wire tmp9264;
  wire tmp9265;
  wire tmp9266;
  wire tmp9267;
  wire tmp9268;
  wire tmp9269;
  wire tmp9270;
  wire tmp9271;
  wire tmp9272;
  wire tmp9273;
  wire tmp9274;
  wire tmp9275;
  wire tmp9276;
  wire tmp9277;
  wire tmp9278;
  wire tmp9279;
  wire tmp9280;
  wire tmp9281;
  wire tmp9282;
  wire tmp9283;
  wire tmp9284;
  wire tmp9285;
  wire tmp9286;
  wire tmp9287;
  wire tmp9288;
  wire tmp9289;
  wire tmp9290;
  wire tmp9291;
  wire tmp9292;
  wire tmp9293;
  wire tmp9294;
  wire tmp9295;
  wire tmp9296;
  wire tmp9297;
  wire tmp9298;
  wire tmp9299;
  wire tmp9300;
  wire tmp9301;
  wire tmp9302;
  wire tmp9303;
  wire tmp9304;
  wire tmp9305;
  wire tmp9306;
  wire tmp9307;
  wire tmp9308;
  wire tmp9309;
  wire tmp9310;
  wire tmp9311;
  wire tmp9312;
  wire tmp9313;
  wire tmp9314;
  wire tmp9315;
  wire tmp9316;
  wire tmp9317;
  wire tmp9318;
  wire tmp9319;
  wire tmp9320;
  wire tmp9321;
  wire tmp9322;
  wire tmp9323;
  wire tmp9324;
  wire tmp9325;
  wire tmp9326;
  wire tmp9327;
  wire tmp9328;
  wire tmp9329;
  wire tmp9330;
  wire tmp9331;
  wire tmp9332;
  wire tmp9333;
  wire tmp9334;
  wire tmp9335;
  wire tmp9336;
  wire tmp9337;
  wire tmp9338;
  wire tmp9339;
  wire tmp9340;
  wire tmp9341;
  wire tmp9342;
  wire tmp9343;
  wire tmp9344;
  wire tmp9345;
  wire tmp9346;
  wire tmp9347;
  wire tmp9348;
  wire tmp9349;
  wire tmp9350;
  wire tmp9351;
  wire tmp9352;
  wire tmp9353;
  wire tmp9354;
  wire tmp9355;
  wire tmp9356;
  wire tmp9357;
  wire tmp9358;
  wire tmp9359;
  wire tmp9360;
  wire tmp9361;
  wire tmp9362;
  wire tmp9363;
  wire tmp9364;
  wire tmp9365;
  wire tmp9366;
  wire tmp9367;
  wire tmp9368;
  wire tmp9369;
  wire tmp9370;
  wire tmp9371;
  wire tmp9372;
  wire tmp9373;
  wire tmp9374;
  wire tmp9375;
  wire tmp9376;
  wire tmp9377;
  wire tmp9378;
  wire tmp9379;
  wire tmp9380;
  wire tmp9381;
  wire tmp9382;
  wire tmp9383;
  wire tmp9384;
  wire tmp9385;
  wire tmp9386;
  wire tmp9387;
  wire tmp9388;
  wire tmp9389;
  wire tmp9390;
  wire tmp9391;
  wire tmp9392;
  wire tmp9393;
  wire tmp9394;
  wire tmp9395;
  wire tmp9396;
  wire tmp9397;
  wire tmp9398;
  wire tmp9399;
  wire tmp9400;
  wire tmp9401;
  wire tmp9402;
  wire tmp9403;
  wire tmp9404;
  wire tmp9405;
  wire tmp9406;
  wire tmp9407;
  wire tmp9408;
  wire tmp9409;
  wire tmp9410;
  wire tmp9411;
  wire tmp9412;
  wire tmp9413;
  wire tmp9414;
  wire tmp9415;
  wire tmp9416;
  wire tmp9417;
  wire tmp9418;
  wire tmp9419;
  wire tmp9420;
  wire tmp9421;
  wire tmp9422;
  wire tmp9423;
  wire tmp9424;
  wire tmp9425;
  wire tmp9426;
  wire tmp9427;
  wire tmp9428;
  wire tmp9429;
  wire tmp9430;
  wire tmp9431;
  wire tmp9432;
  wire tmp9433;
  wire tmp9434;
  wire tmp9435;
  wire tmp9436;
  wire tmp9437;
  wire tmp9438;
  wire tmp9439;
  wire tmp9440;
  wire tmp9441;
  wire tmp9442;
  wire tmp9443;
  wire tmp9444;
  wire tmp9445;
  wire tmp9446;
  wire tmp9447;
  wire tmp9448;
  wire tmp9449;
  wire tmp9450;
  wire tmp9451;
  wire tmp9452;
  wire tmp9453;
  wire tmp9454;
  wire tmp9455;
  wire tmp9456;
  wire tmp9457;
  wire tmp9458;
  wire tmp9459;
  wire tmp9460;
  wire tmp9461;
  wire tmp9462;
  wire tmp9463;
  wire tmp9464;
  wire tmp9465;
  wire tmp9466;
  wire tmp9467;
  wire tmp9468;
  wire tmp9469;
  wire tmp9470;
  wire tmp9471;
  wire tmp9472;
  wire tmp9473;
  wire tmp9474;
  wire tmp9475;
  wire tmp9476;
  wire tmp9477;
  wire tmp9478;
  wire tmp9479;
  wire tmp9480;
  wire tmp9481;
  wire tmp9482;
  wire tmp9483;
  wire tmp9484;
  wire tmp9485;
  wire tmp9486;
  wire tmp9487;
  wire tmp9488;
  wire tmp9489;
  wire tmp9490;
  wire tmp9491;
  wire tmp9492;
  wire tmp9493;
  wire tmp9494;
  wire tmp9495;
  wire tmp9496;
  wire tmp9497;
  wire tmp9498;
  wire tmp9499;
  wire tmp9500;
  wire tmp9501;
  wire tmp9502;
  wire tmp9503;
  wire tmp9504;
  wire tmp9505;
  wire tmp9506;
  wire tmp9507;
  wire tmp9508;
  wire tmp9509;
  wire tmp9510;
  wire tmp9511;
  wire tmp9512;
  wire tmp9513;
  wire tmp9514;
  wire tmp9515;
  wire tmp9516;
  wire tmp9517;
  wire tmp9518;
  wire tmp9519;
  wire tmp9520;
  wire tmp9521;
  wire tmp9522;
  wire tmp9523;
  wire tmp9524;
  wire tmp9525;
  wire tmp9526;
  wire tmp9527;
  wire tmp9528;
  wire tmp9529;
  wire tmp9530;
  wire tmp9531;
  wire tmp9532;
  wire tmp9533;
  wire tmp9534;
  wire tmp9535;
  wire tmp9536;
  wire tmp9537;
  wire tmp9538;
  wire tmp9539;
  wire tmp9540;
  wire tmp9541;
  wire tmp9542;
  wire tmp9543;
  wire tmp9544;
  wire tmp9545;
  wire tmp9546;
  wire tmp9547;
  wire tmp9548;
  wire tmp9549;
  wire tmp9550;
  wire tmp9551;
  wire tmp9552;
  wire tmp9553;
  wire tmp9554;
  wire tmp9555;
  wire tmp9556;
  wire tmp9557;
  wire tmp9558;
  wire tmp9559;
  wire tmp9560;
  wire tmp9561;
  wire tmp9562;
  wire tmp9563;
  wire tmp9564;
  wire tmp9565;
  wire tmp9566;
  wire tmp9567;
  wire tmp9568;
  wire tmp9569;
  wire tmp9570;
  wire tmp9571;
  wire tmp9572;
  wire tmp9573;
  wire tmp9574;
  wire tmp9575;
  wire tmp9576;
  wire tmp9577;
  wire tmp9578;
  wire tmp9579;
  wire tmp9580;
  wire tmp9581;
  wire tmp9582;
  wire tmp9583;
  wire tmp9584;
  wire tmp9585;
  wire tmp9586;
  wire tmp9587;
  wire tmp9588;
  wire tmp9589;
  wire tmp9590;
  wire tmp9591;
  wire tmp9592;
  wire tmp9593;
  wire tmp9594;
  wire tmp9595;
  wire tmp9596;
  wire tmp9597;
  wire tmp9598;
  wire tmp9599;
  wire tmp9600;
  wire tmp9601;
  wire tmp9602;
  wire tmp9603;
  wire tmp9604;
  wire tmp9605;
  wire tmp9606;
  wire tmp9607;
  wire tmp9608;
  wire tmp9609;
  wire tmp9610;
  wire tmp9611;
  wire tmp9612;
  wire tmp9613;
  wire tmp9614;
  wire tmp9615;
  wire tmp9616;
  wire tmp9617;
  wire tmp9618;
  wire tmp9619;
  wire tmp9620;
  wire tmp9621;
  wire tmp9622;
  wire tmp9623;
  wire tmp9624;
  wire tmp9625;
  wire tmp9626;
  wire tmp9627;
  wire tmp9628;
  wire tmp9629;
  wire tmp9630;
  wire tmp9631;
  wire tmp9632;
  wire tmp9633;
  wire tmp9634;
  wire tmp9635;
  wire tmp9636;
  wire tmp9637;
  wire tmp9638;
  wire tmp9639;
  wire tmp9640;
  wire tmp9641;
  wire tmp9642;
  wire tmp9643;
  wire tmp9644;
  wire tmp9645;
  wire tmp9646;
  wire tmp9647;
  wire tmp9648;
  wire tmp9649;
  wire tmp9650;
  wire tmp9651;
  wire tmp9652;
  wire tmp9653;
  wire tmp9654;
  wire tmp9655;
  wire tmp9656;
  wire tmp9657;
  wire tmp9658;
  wire tmp9659;
  wire tmp9660;
  wire tmp9661;
  wire tmp9662;
  wire tmp9663;
  wire tmp9664;
  wire tmp9665;
  wire tmp9666;
  wire tmp9667;
  wire tmp9668;
  wire tmp9669;
  wire tmp9670;
  wire tmp9671;
  wire tmp9672;
  wire tmp9673;
  wire tmp9674;
  wire tmp9675;
  wire tmp9676;
  wire tmp9677;
  wire tmp9678;
  wire tmp9679;
  wire tmp9680;
  wire tmp9681;
  wire tmp9682;
  wire tmp9683;
  wire tmp9684;
  wire tmp9685;
  wire tmp9686;
  wire tmp9687;
  wire tmp9688;
  wire tmp9689;
  wire tmp9690;
  wire tmp9691;
  wire tmp9692;
  wire tmp9693;
  wire tmp9694;
  wire tmp9695;
  wire tmp9696;
  wire tmp9697;
  wire tmp9698;
  wire tmp9699;
  wire tmp9700;
  wire tmp9701;
  wire tmp9702;
  wire tmp9703;
  wire tmp9704;
  wire tmp9705;
  wire tmp9706;
  wire tmp9707;
  wire tmp9708;
  wire tmp9709;
  wire tmp9710;
  wire tmp9711;
  wire tmp9712;
  wire tmp9713;
  wire tmp9714;
  wire tmp9715;
  wire tmp9716;
  wire tmp9717;
  wire tmp9718;
  wire tmp9719;
  wire tmp9720;
  wire tmp9721;
  wire tmp9722;
  wire tmp9723;
  wire tmp9724;
  wire tmp9725;
  wire tmp9726;
  wire tmp9727;
  wire tmp9728;
  wire tmp9729;
  wire tmp9730;
  wire tmp9731;
  wire tmp9732;
  wire tmp9733;
  wire tmp9734;
  wire tmp9735;
  wire tmp9736;
  wire tmp9737;
  wire tmp9738;
  wire tmp9739;
  wire tmp9740;
  wire tmp9741;
  wire tmp9742;
  wire tmp9743;
  wire tmp9744;
  wire tmp9745;
  wire tmp9746;
  wire tmp9747;
  wire tmp9748;
  wire tmp9749;
  wire tmp9750;
  wire tmp9751;
  wire tmp9752;
  wire tmp9753;
  wire tmp9754;
  wire tmp9755;
  wire tmp9756;
  wire tmp9757;
  wire tmp9758;
  wire tmp9759;
  wire tmp9760;
  wire tmp9761;
  wire tmp9762;
  wire tmp9763;
  wire tmp9764;
  wire tmp9765;
  wire tmp9766;
  wire tmp9767;
  wire tmp9768;
  wire tmp9769;
  wire tmp9770;
  wire tmp9771;
  wire tmp9772;
  wire tmp9773;
  wire tmp9774;
  wire tmp9775;
  wire tmp9776;
  wire tmp9777;
  wire tmp9778;
  wire tmp9779;
  wire tmp9780;
  wire tmp9781;
  wire tmp9782;
  wire tmp9783;
  wire tmp9784;
  wire tmp9785;
  wire tmp9786;
  wire tmp9787;
  wire tmp9788;
  wire tmp9789;
  wire tmp9790;
  wire tmp9791;
  wire tmp9792;
  wire tmp9793;
  wire tmp9794;
  wire tmp9795;
  wire tmp9796;
  wire tmp9797;
  wire tmp9798;
  wire tmp9799;
  wire tmp9800;
  wire tmp9801;
  wire tmp9802;
  wire tmp9803;
  wire tmp9804;
  wire tmp9805;
  wire tmp9806;
  wire tmp9807;
  wire tmp9808;
  wire tmp9809;
  wire tmp9810;
  wire tmp9811;
  wire tmp9812;
  wire tmp9813;
  wire tmp9814;
  wire tmp9815;
  wire tmp9816;
  wire tmp9817;
  wire tmp9818;
  wire tmp9819;
  wire tmp9820;
  wire tmp9821;
  wire tmp9822;
  wire tmp9823;
  wire tmp9824;
  wire tmp9825;
  wire tmp9826;
  wire tmp9827;
  wire tmp9828;
  wire tmp9829;
  wire tmp9830;
  wire tmp9831;
  wire tmp9832;
  wire tmp9833;
  wire tmp9834;
  wire tmp9835;
  wire tmp9836;
  wire tmp9837;
  wire tmp9838;
  wire tmp9839;
  wire tmp9840;
  wire tmp9841;
  wire tmp9842;
  wire tmp9843;
  wire tmp9844;
  wire tmp9845;
  wire tmp9846;
  wire tmp9847;
  wire tmp9848;
  wire tmp9849;
  wire tmp9850;
  wire tmp9851;
  wire tmp9852;
  wire tmp9853;
  wire tmp9854;
  wire tmp9855;
  wire tmp9856;
  wire tmp9857;
  wire tmp9858;
  wire tmp9859;
  wire tmp9860;
  wire tmp9861;
  wire tmp9862;
  wire tmp9863;
  wire tmp9864;
  wire tmp9865;
  wire tmp9866;
  wire tmp9867;
  wire tmp9868;
  wire tmp9869;
  wire tmp9870;
  wire tmp9871;
  wire tmp9872;
  wire tmp9873;
  wire tmp9874;
  wire tmp9875;
  wire tmp9876;
  wire tmp9877;
  wire tmp9878;
  wire tmp9879;
  wire tmp9880;
  wire tmp9881;
  wire tmp9882;
  wire tmp9883;
  wire tmp9884;
  wire tmp9885;
  wire tmp9886;
  wire tmp9887;
  wire tmp9888;
  wire tmp9889;
  wire tmp9890;
  wire tmp9891;
  wire tmp9892;
  wire tmp9893;
  wire tmp9894;
  wire tmp9895;
  wire tmp9896;
  wire tmp9897;
  wire tmp9898;
  wire tmp9899;
  wire tmp9900;
  wire tmp9901;
  wire tmp9902;
  wire tmp9903;
  wire tmp9904;
  wire tmp9905;
  wire tmp9906;
  wire tmp9907;
  wire tmp9908;
  wire tmp9909;
  wire tmp9910;
  wire tmp9911;
  wire tmp9912;
  wire tmp9913;
  wire tmp9914;
  wire tmp9915;
  wire tmp9916;
  wire tmp9917;
  wire tmp9918;
  wire tmp9919;
  wire tmp9920;
  wire tmp9921;
  wire tmp9922;
  wire tmp9923;
  wire tmp9924;
  wire tmp9925;
  wire tmp9926;
  wire tmp9927;
  wire tmp9928;
  wire tmp9929;
  wire tmp9930;
  wire tmp9931;
  wire tmp9932;
  wire tmp9933;
  wire tmp9934;
  wire tmp9935;
  wire tmp9936;
  wire tmp9937;
  wire tmp9938;
  wire tmp9939;
  wire tmp9940;
  wire tmp9941;
  wire tmp9942;
  wire tmp9943;
  wire tmp9944;
  wire tmp9945;
  wire tmp9946;
  wire tmp9947;
  wire tmp9948;
  wire tmp9949;
  wire tmp9950;
  wire tmp9951;
  wire tmp9952;
  wire tmp9953;
  wire tmp9954;
  wire tmp9955;
  wire tmp9956;
  wire tmp9957;
  wire tmp9958;
  wire tmp9959;
  wire tmp9960;
  wire tmp9961;
  wire tmp9962;
  wire tmp9963;
  wire tmp9964;
  wire tmp9965;
  wire tmp9966;
  wire tmp9967;
  wire tmp9968;
  wire tmp9969;
  wire tmp9970;
  wire tmp9971;
  wire tmp9972;
  wire tmp9973;
  wire tmp9974;
  wire tmp9975;
  wire tmp9976;
  wire tmp9977;
  wire tmp9978;
  wire tmp9979;
  wire tmp9980;
  wire tmp9981;
  wire tmp9982;
  wire tmp9983;
  wire tmp9984;
  wire tmp9985;
  wire tmp9986;
  wire tmp9987;
  wire tmp9988;
  wire tmp9989;
  wire tmp9990;
  wire tmp9991;
  wire tmp9992;
  wire tmp9993;
  wire tmp9994;
  wire tmp9995;
  wire tmp9996;
  wire tmp9997;
  wire tmp9998;
  wire tmp9999;
  wire tmp10000;
  wire tmp10001;
  wire tmp10002;
  wire tmp10003;
  wire tmp10004;
  wire tmp10005;
  wire tmp10006;
  wire tmp10007;
  wire tmp10008;
  wire tmp10009;
  wire tmp10010;
  wire tmp10011;
  wire tmp10012;
  wire tmp10013;
  wire tmp10014;
  wire tmp10015;
  wire tmp10016;
  wire tmp10017;
  wire tmp10018;
  wire tmp10019;
  wire tmp10020;
  wire tmp10021;
  wire tmp10022;
  wire tmp10023;
  wire tmp10024;
  wire tmp10025;
  wire tmp10026;
  wire tmp10027;
  wire tmp10028;
  wire tmp10029;
  wire tmp10030;
  wire tmp10031;
  wire tmp10032;
  wire tmp10033;
  wire tmp10034;
  wire tmp10035;
  wire tmp10036;
  wire tmp10037;
  wire tmp10038;
  wire tmp10039;
  wire tmp10040;
  wire tmp10041;
  wire tmp10042;
  wire tmp10043;
  wire tmp10044;
  wire tmp10045;
  wire tmp10046;
  wire tmp10047;
  wire tmp10048;
  wire tmp10049;
  wire tmp10050;
  wire tmp10051;
  wire tmp10052;
  wire tmp10053;
  wire tmp10054;
  wire tmp10055;
  wire tmp10056;
  wire tmp10057;
  wire tmp10058;
  wire tmp10059;
  wire tmp10060;
  wire tmp10061;
  wire tmp10062;
  wire tmp10063;
  wire tmp10064;
  wire tmp10065;
  wire tmp10066;
  wire tmp10067;
  wire tmp10068;
  wire tmp10069;
  wire tmp10070;
  wire tmp10071;
  wire tmp10072;
  wire tmp10073;
  wire tmp10074;
  wire tmp10075;
  wire tmp10076;
  wire tmp10077;
  wire tmp10078;
  wire tmp10079;
  wire tmp10080;
  wire tmp10081;
  wire tmp10082;
  wire tmp10083;
  wire tmp10084;
  wire tmp10085;
  wire tmp10086;
  wire tmp10087;
  wire tmp10088;
  wire tmp10089;
  wire tmp10090;
  wire tmp10091;
  wire tmp10092;
  wire tmp10093;
  wire tmp10094;
  wire tmp10095;
  wire tmp10096;
  wire tmp10097;
  wire tmp10098;
  wire tmp10099;
  wire tmp10100;
  wire tmp10101;
  wire tmp10102;
  wire tmp10103;
  wire tmp10104;
  wire tmp10105;
  wire tmp10106;
  wire tmp10107;
  wire tmp10108;
  wire tmp10109;
  wire tmp10110;
  wire tmp10111;
  wire tmp10112;
  wire tmp10113;
  wire tmp10114;
  wire tmp10115;
  wire tmp10116;
  wire tmp10117;
  wire tmp10118;
  wire tmp10119;
  wire tmp10120;
  wire tmp10121;
  wire tmp10122;
  wire tmp10123;
  wire tmp10124;
  wire tmp10125;
  wire tmp10126;
  wire tmp10127;
  wire tmp10128;
  wire tmp10129;
  wire tmp10130;
  wire tmp10131;
  wire tmp10132;
  wire tmp10133;
  wire tmp10134;
  wire tmp10135;
  wire tmp10136;
  wire tmp10137;
  wire tmp10138;
  wire tmp10139;
  wire tmp10140;
  wire tmp10141;
  wire tmp10142;
  wire tmp10143;
  wire tmp10144;
  wire tmp10145;
  wire tmp10146;
  wire tmp10147;
  wire tmp10148;
  wire tmp10149;
  wire tmp10150;
  wire tmp10151;
  wire tmp10152;
  wire tmp10153;
  wire tmp10154;
  wire tmp10155;
  wire tmp10156;
  wire tmp10157;
  wire tmp10158;
  wire tmp10159;
  wire tmp10160;
  wire tmp10161;
  wire tmp10162;
  wire tmp10163;
  wire tmp10164;
  wire tmp10165;
  wire tmp10166;
  wire tmp10167;
  wire tmp10168;
  wire tmp10169;
  wire tmp10170;
  wire tmp10171;
  wire tmp10172;
  wire tmp10173;
  wire tmp10174;
  wire tmp10175;
  wire tmp10176;
  wire tmp10177;
  wire tmp10178;
  wire tmp10179;
  wire tmp10180;
  wire tmp10181;
  wire tmp10182;
  wire tmp10183;
  wire tmp10184;
  wire tmp10185;
  wire tmp10186;
  wire tmp10187;
  wire tmp10188;
  wire tmp10189;
  wire tmp10190;
  wire tmp10191;
  wire tmp10192;
  wire tmp10193;
  wire tmp10194;
  wire tmp10195;
  wire tmp10196;
  wire tmp10197;
  wire tmp10198;
  wire tmp10199;
  wire tmp10200;
  wire tmp10201;
  wire tmp10202;
  wire tmp10203;
  wire tmp10204;
  wire tmp10205;
  wire tmp10206;
  wire tmp10207;
  wire tmp10208;
  wire tmp10209;
  wire tmp10210;
  wire tmp10211;
  wire tmp10212;
  wire tmp10213;
  wire tmp10214;
  wire tmp10215;
  wire tmp10216;
  wire tmp10217;
  wire tmp10218;
  wire tmp10219;
  wire tmp10220;
  wire tmp10221;
  wire tmp10222;
  wire tmp10223;
  wire tmp10224;
  wire tmp10225;
  wire tmp10226;
  wire tmp10227;
  wire tmp10228;
  wire tmp10229;
  wire tmp10230;
  wire tmp10231;
  wire tmp10232;
  wire tmp10233;
  wire tmp10234;
  wire tmp10235;
  wire tmp10236;
  wire tmp10237;
  wire tmp10238;
  wire tmp10239;
  wire tmp10240;
  wire tmp10241;
  wire tmp10242;
  wire tmp10243;
  wire tmp10244;
  wire tmp10245;
  wire tmp10246;
  wire tmp10247;
  wire tmp10248;
  wire tmp10249;
  wire tmp10250;
  wire tmp10251;
  wire tmp10252;
  wire tmp10253;
  wire tmp10254;
  wire tmp10255;
  wire tmp10256;
  wire tmp10257;
  wire tmp10258;
  wire tmp10259;
  wire tmp10260;
  wire tmp10261;
  wire tmp10262;
  wire tmp10263;
  wire tmp10264;
  wire tmp10265;
  wire tmp10266;
  wire tmp10267;
  wire tmp10268;
  wire tmp10269;
  wire tmp10270;
  wire tmp10271;
  wire tmp10272;
  wire tmp10273;
  wire tmp10274;
  wire tmp10275;
  wire tmp10276;
  wire tmp10277;
  wire tmp10278;
  wire tmp10279;
  wire tmp10280;
  wire tmp10281;
  wire tmp10282;
  wire tmp10283;
  wire tmp10284;
  wire tmp10285;
  wire tmp10286;
  wire tmp10287;
  wire tmp10288;
  wire tmp10289;
  wire tmp10290;
  wire tmp10291;
  wire tmp10292;
  wire tmp10293;
  wire tmp10294;
  wire tmp10295;
  wire tmp10296;
  wire tmp10297;
  wire tmp10298;
  wire tmp10299;
  wire tmp10300;
  wire tmp10301;
  wire tmp10302;
  wire tmp10303;
  wire tmp10304;
  wire tmp10305;
  wire tmp10306;
  wire tmp10307;
  wire tmp10308;
  wire tmp10309;
  wire tmp10310;
  wire tmp10311;
  wire tmp10312;
  wire tmp10313;
  wire tmp10314;
  wire tmp10315;
  wire tmp10316;
  wire tmp10317;
  wire tmp10318;
  wire tmp10319;
  wire tmp10320;
  wire tmp10321;
  wire tmp10322;
  wire tmp10323;
  wire tmp10324;
  wire tmp10325;
  wire tmp10326;
  wire tmp10327;
  wire tmp10328;
  wire tmp10329;
  wire tmp10330;
  wire tmp10331;
  wire tmp10332;
  wire tmp10333;
  wire tmp10334;
  wire tmp10335;
  wire tmp10336;
  wire tmp10337;
  wire tmp10338;
  wire tmp10339;
  wire tmp10340;
  wire tmp10341;
  wire tmp10342;
  wire tmp10343;
  wire tmp10344;
  wire tmp10345;
  wire tmp10346;
  wire tmp10347;
  wire tmp10348;
  wire tmp10349;
  wire tmp10350;
  wire tmp10351;
  wire tmp10352;
  wire tmp10353;
  wire tmp10354;
  wire tmp10355;
  wire tmp10356;
  wire tmp10357;
  wire tmp10358;
  wire tmp10359;
  wire tmp10360;
  wire tmp10361;
  wire tmp10362;
  wire tmp10363;
  wire tmp10364;
  wire tmp10365;
  wire tmp10366;
  wire tmp10367;
  wire tmp10368;
  wire tmp10369;
  wire tmp10370;
  wire tmp10371;
  wire tmp10372;
  wire tmp10373;
  wire tmp10374;
  wire tmp10375;
  wire tmp10376;
  wire tmp10377;
  wire tmp10378;
  wire tmp10379;
  wire tmp10380;
  wire tmp10381;
  wire tmp10382;
  wire tmp10383;
  wire tmp10384;
  wire tmp10385;
  wire tmp10386;
  wire tmp10387;
  wire tmp10388;
  wire tmp10389;
  wire tmp10390;
  wire tmp10391;
  wire tmp10392;
  wire tmp10393;
  wire tmp10394;
  wire tmp10395;
  wire tmp10396;
  wire tmp10397;
  wire tmp10398;
  wire tmp10399;
  wire tmp10400;
  wire tmp10401;
  wire tmp10402;
  wire tmp10403;
  wire tmp10404;
  wire tmp10405;
  wire tmp10406;
  wire tmp10407;
  wire tmp10408;
  wire tmp10409;
  wire tmp10410;
  wire tmp10411;
  wire tmp10412;
  wire tmp10413;
  wire tmp10414;
  wire tmp10415;
  wire tmp10416;
  wire tmp10417;
  wire tmp10418;
  wire tmp10419;
  wire tmp10420;
  wire tmp10421;
  wire tmp10422;
  wire tmp10423;
  wire tmp10424;
  wire tmp10425;
  wire tmp10426;
  wire tmp10427;
  wire tmp10428;
  wire tmp10429;
  wire tmp10430;
  wire tmp10431;
  wire tmp10432;
  wire tmp10433;
  wire tmp10434;
  wire tmp10435;
  wire tmp10436;
  wire tmp10437;
  wire tmp10438;
  wire tmp10439;
  wire tmp10440;
  wire tmp10441;
  wire tmp10442;
  wire tmp10443;
  wire tmp10444;
  wire tmp10445;
  wire tmp10446;
  wire tmp10447;
  wire tmp10448;
  wire tmp10449;
  wire tmp10450;
  wire tmp10451;
  wire tmp10452;
  wire tmp10453;
  wire tmp10454;
  wire tmp10455;
  wire tmp10456;
  wire tmp10457;
  wire tmp10458;
  wire tmp10459;
  wire tmp10460;
  wire tmp10461;
  wire tmp10462;
  wire tmp10463;
  wire tmp10464;
  wire tmp10465;
  wire tmp10466;
  wire tmp10467;
  wire tmp10468;
  wire tmp10469;
  wire tmp10470;
  wire tmp10471;
  wire tmp10472;
  wire tmp10473;
  wire tmp10474;
  wire tmp10475;
  wire tmp10476;
  wire tmp10477;
  wire tmp10478;
  wire tmp10479;
  wire tmp10480;
  wire tmp10481;
  wire tmp10482;
  wire tmp10483;
  wire tmp10484;
  wire tmp10485;
  wire tmp10486;
  wire tmp10487;
  wire tmp10488;
  wire tmp10489;
  wire tmp10490;
  wire tmp10491;
  wire tmp10492;
  wire tmp10493;
  wire tmp10494;
  wire tmp10495;
  wire tmp10496;
  wire tmp10497;
  wire tmp10498;
  wire tmp10499;
  wire tmp10500;
  wire tmp10501;
  wire tmp10502;
  wire tmp10503;
  wire tmp10504;
  wire tmp10505;
  wire tmp10506;
  wire tmp10507;
  wire tmp10508;
  wire tmp10509;
  wire tmp10510;
  wire tmp10511;
  wire tmp10512;
  wire tmp10513;
  wire tmp10514;
  wire tmp10515;
  wire tmp10516;
  wire tmp10517;
  wire tmp10518;
  wire tmp10519;
  wire tmp10520;
  wire tmp10521;
  wire tmp10522;
  wire tmp10523;
  wire tmp10524;
  wire tmp10525;
  wire tmp10526;
  wire tmp10527;
  wire tmp10528;
  wire tmp10529;
  wire tmp10530;
  wire tmp10531;
  wire tmp10532;
  wire tmp10533;
  wire tmp10534;
  wire tmp10535;
  wire tmp10536;
  wire tmp10537;
  wire tmp10538;
  wire tmp10539;
  wire tmp10540;
  wire tmp10541;
  wire tmp10542;
  wire tmp10543;
  wire tmp10544;
  wire tmp10545;
  wire tmp10546;
  wire tmp10547;
  wire tmp10548;
  wire tmp10549;
  wire tmp10550;
  wire tmp10551;
  wire tmp10552;
  wire tmp10553;
  wire tmp10554;
  wire tmp10555;
  wire tmp10556;
  wire tmp10557;
  wire tmp10558;
  wire tmp10559;
  wire tmp10560;
  wire tmp10561;
  wire tmp10562;
  wire tmp10563;
  wire tmp10564;
  wire tmp10565;
  wire tmp10566;
  wire tmp10567;
  wire tmp10568;
  wire tmp10569;
  wire tmp10570;
  wire tmp10571;
  wire tmp10572;
  wire tmp10573;
  wire tmp10574;
  wire tmp10575;
  wire tmp10576;
  wire tmp10577;
  wire tmp10578;
  wire tmp10579;
  wire tmp10580;
  wire tmp10581;
  wire tmp10582;
  wire tmp10583;
  wire tmp10584;
  wire tmp10585;
  wire tmp10586;
  wire tmp10587;
  wire tmp10588;
  wire tmp10589;
  wire tmp10590;
  wire tmp10591;
  wire tmp10592;
  wire tmp10593;
  wire tmp10594;
  wire tmp10595;
  wire tmp10596;
  wire tmp10597;
  wire tmp10598;
  wire tmp10599;
  wire tmp10600;
  wire tmp10601;
  wire tmp10602;
  wire tmp10603;
  wire tmp10604;
  wire tmp10605;
  wire tmp10606;
  wire tmp10607;
  wire tmp10608;
  wire tmp10609;
  wire tmp10610;
  wire tmp10611;
  wire tmp10612;
  wire tmp10613;
  wire tmp10614;
  wire tmp10615;
  wire tmp10616;
  wire tmp10617;
  wire tmp10618;
  wire tmp10619;
  wire tmp10620;
  wire tmp10621;
  wire tmp10622;
  wire tmp10623;
  wire tmp10624;
  wire tmp10625;
  wire tmp10626;
  wire tmp10627;
  wire tmp10628;
  wire tmp10629;
  wire tmp10630;
  wire tmp10631;
  wire tmp10632;
  wire tmp10633;
  wire tmp10634;
  wire tmp10635;
  wire tmp10636;
  wire tmp10637;
  wire tmp10638;
  wire tmp10639;
  wire tmp10640;
  wire tmp10641;
  wire tmp10642;
  wire tmp10643;
  wire tmp10644;
  wire tmp10645;
  wire tmp10646;
  wire tmp10647;
  wire tmp10648;
  wire tmp10649;
  wire tmp10650;
  wire tmp10651;
  wire tmp10652;
  wire tmp10653;
  wire tmp10654;
  wire tmp10655;
  wire tmp10656;
  wire tmp10657;
  wire tmp10658;
  wire tmp10659;
  wire tmp10660;
  wire tmp10661;
  wire tmp10662;
  wire tmp10663;
  wire tmp10664;
  wire tmp10665;
  wire tmp10666;
  wire tmp10667;
  wire tmp10668;
  wire tmp10669;
  wire tmp10670;
  wire tmp10671;
  wire tmp10672;
  wire tmp10673;
  wire tmp10674;
  wire tmp10675;
  wire tmp10676;
  wire tmp10677;
  wire tmp10678;
  wire tmp10679;
  wire tmp10680;
  wire tmp10681;
  wire tmp10682;
  wire tmp10683;
  wire tmp10684;
  wire tmp10685;
  wire tmp10686;
  wire tmp10687;
  wire tmp10688;
  wire tmp10689;
  wire tmp10690;
  wire tmp10691;
  wire tmp10692;
  wire tmp10693;
  wire tmp10694;
  wire tmp10695;
  wire tmp10696;
  wire tmp10697;
  wire tmp10698;
  wire tmp10699;
  wire tmp10700;
  wire tmp10701;
  wire tmp10702;
  wire tmp10703;
  wire tmp10704;
  wire tmp10705;
  wire tmp10706;
  wire tmp10707;
  wire tmp10708;
  wire tmp10709;
  wire tmp10710;
  wire tmp10711;
  wire tmp10712;
  wire tmp10713;
  wire tmp10714;
  wire tmp10715;
  wire tmp10716;
  wire tmp10717;
  wire tmp10718;
  wire tmp10719;
  wire tmp10720;
  wire tmp10721;
  wire tmp10722;
  wire tmp10723;
  wire tmp10724;
  wire tmp10725;
  wire tmp10726;
  wire tmp10727;
  wire tmp10728;
  wire tmp10729;
  wire tmp10730;
  wire tmp10731;
  wire tmp10732;
  wire tmp10733;
  wire tmp10734;
  wire tmp10735;
  wire tmp10736;
  wire tmp10737;
  wire tmp10738;
  wire tmp10739;
  wire tmp10740;
  wire tmp10741;
  wire tmp10742;
  wire tmp10743;
  wire tmp10744;
  wire tmp10745;
  wire tmp10746;
  wire tmp10747;
  wire tmp10748;
  wire tmp10749;
  wire tmp10750;
  wire tmp10751;
  wire tmp10752;
  wire tmp10753;
  wire tmp10754;
  wire tmp10755;
  wire tmp10756;
  wire tmp10757;
  wire tmp10758;
  wire tmp10759;
  wire tmp10760;
  wire tmp10761;
  wire tmp10762;
  wire tmp10763;
  wire tmp10764;
  wire tmp10765;
  wire tmp10766;
  wire tmp10767;
  wire tmp10768;
  wire tmp10769;
  wire tmp10770;
  wire tmp10771;
  wire tmp10772;
  wire tmp10773;
  wire tmp10774;
  wire tmp10775;
  wire tmp10776;
  wire tmp10777;
  wire tmp10778;
  wire tmp10779;
  wire tmp10780;
  wire tmp10781;
  wire tmp10782;
  wire tmp10783;
  wire tmp10784;
  wire tmp10785;
  wire tmp10786;
  wire tmp10787;
  wire tmp10788;
  wire tmp10789;
  wire tmp10790;
  wire tmp10791;
  wire tmp10792;
  wire tmp10793;
  wire tmp10794;
  wire tmp10795;
  wire tmp10796;
  wire tmp10797;
  wire tmp10798;
  wire tmp10799;
  wire tmp10800;
  wire tmp10801;
  wire tmp10802;
  wire tmp10803;
  wire tmp10804;
  wire tmp10805;
  wire tmp10806;
  wire tmp10807;
  wire tmp10808;
  wire tmp10809;
  wire tmp10810;
  wire tmp10811;
  wire tmp10812;
  wire tmp10813;
  wire tmp10814;
  wire tmp10815;
  wire tmp10816;
  wire tmp10817;
  wire tmp10818;
  wire tmp10819;
  wire tmp10820;
  wire tmp10821;
  wire tmp10822;
  wire tmp10823;
  wire tmp10824;
  wire tmp10825;
  wire tmp10826;
  wire tmp10827;
  wire tmp10828;
  wire tmp10829;
  wire tmp10830;
  wire tmp10831;
  wire tmp10832;
  wire tmp10833;
  wire tmp10834;
  wire tmp10835;
  wire tmp10836;
  wire tmp10837;
  wire tmp10838;
  wire tmp10839;
  wire tmp10840;
  wire tmp10841;
  wire tmp10842;
  wire tmp10843;
  wire tmp10844;
  wire tmp10845;
  wire tmp10846;
  wire tmp10847;
  wire tmp10848;
  wire tmp10849;
  wire tmp10850;
  wire tmp10851;
  wire tmp10852;
  wire tmp10853;
  wire tmp10854;
  wire tmp10855;
  wire tmp10856;
  wire tmp10857;
  wire tmp10858;
  wire tmp10859;
  wire tmp10860;
  wire tmp10861;
  wire tmp10862;
  wire tmp10863;
  wire tmp10864;
  wire tmp10865;
  wire tmp10866;
  wire tmp10867;
  wire tmp10868;
  wire tmp10869;
  wire tmp10870;
  wire tmp10871;
  wire tmp10872;
  wire tmp10873;
  wire tmp10874;
  wire tmp10875;
  wire tmp10876;
  wire tmp10877;
  wire tmp10878;
  wire tmp10879;
  wire tmp10880;
  wire tmp10881;
  wire tmp10882;
  wire tmp10883;
  wire tmp10884;
  wire tmp10885;
  wire tmp10886;
  wire tmp10887;
  wire tmp10888;
  wire tmp10889;
  wire tmp10890;
  wire tmp10891;
  wire tmp10892;
  wire tmp10893;
  wire tmp10894;
  wire tmp10895;
  wire tmp10896;
  wire tmp10897;
  wire tmp10898;
  wire tmp10899;
  wire tmp10900;
  wire tmp10901;
  wire tmp10902;
  wire tmp10903;
  wire tmp10904;
  wire tmp10905;
  wire tmp10906;
  wire tmp10907;
  wire tmp10908;
  wire tmp10909;
  wire tmp10910;
  wire tmp10911;
  wire tmp10912;
  wire tmp10913;
  wire tmp10914;
  wire tmp10915;
  wire tmp10916;
  wire tmp10917;
  wire tmp10918;
  wire tmp10919;
  wire tmp10920;
  wire tmp10921;
  wire tmp10922;
  wire tmp10923;
  wire tmp10924;
  wire tmp10925;
  wire tmp10926;
  wire tmp10927;
  wire tmp10928;
  wire tmp10929;
  wire tmp10930;
  wire tmp10931;
  wire tmp10932;
  wire tmp10933;
  wire tmp10934;
  wire tmp10935;
  wire tmp10936;
  wire tmp10937;
  wire tmp10938;
  wire tmp10939;
  wire tmp10940;
  wire tmp10941;
  wire tmp10942;
  wire tmp10943;
  wire tmp10944;
  wire tmp10945;
  wire tmp10946;
  wire tmp10947;
  wire tmp10948;
  wire tmp10949;
  wire tmp10950;
  wire tmp10951;
  wire tmp10952;
  wire tmp10953;
  wire tmp10954;
  wire tmp10955;
  wire tmp10956;
  wire tmp10957;
  wire tmp10958;
  wire tmp10959;
  wire tmp10960;
  wire tmp10961;
  wire tmp10962;
  wire tmp10963;
  wire tmp10964;
  wire tmp10965;
  wire tmp10966;
  wire tmp10967;
  wire tmp10968;
  wire tmp10969;
  wire tmp10970;
  wire tmp10971;
  wire tmp10972;
  wire tmp10973;
  wire tmp10974;
  wire tmp10975;
  wire tmp10976;
  wire tmp10977;
  wire tmp10978;
  wire tmp10979;
  wire tmp10980;
  wire tmp10981;
  wire tmp10982;
  wire tmp10983;
  wire tmp10984;
  wire tmp10985;
  wire tmp10986;
  wire tmp10987;
  wire tmp10988;
  wire tmp10989;
  wire tmp10990;
  wire tmp10991;
  wire tmp10992;
  wire tmp10993;
  wire tmp10994;
  wire tmp10995;
  wire tmp10996;
  wire tmp10997;
  wire tmp10998;
  wire tmp10999;
  wire tmp11000;
  wire tmp11001;
  wire tmp11002;
  wire tmp11003;
  wire tmp11004;
  wire tmp11005;
  wire tmp11006;
  wire tmp11007;
  wire tmp11008;
  wire tmp11009;
  wire tmp11010;
  wire tmp11011;
  wire tmp11012;
  wire tmp11013;
  wire tmp11014;
  wire tmp11015;
  wire tmp11016;
  wire tmp11017;
  wire tmp11018;
  wire tmp11019;
  wire tmp11020;
  wire tmp11021;
  wire tmp11022;
  wire tmp11023;
  wire tmp11024;
  wire tmp11025;
  wire tmp11026;
  wire tmp11027;
  wire tmp11028;
  wire tmp11029;
  wire tmp11030;
  wire tmp11031;
  wire tmp11032;
  wire tmp11033;
  wire tmp11034;
  wire tmp11035;
  wire tmp11036;
  wire tmp11037;
  wire tmp11038;
  wire tmp11039;
  wire tmp11040;
  wire tmp11041;
  wire tmp11042;
  wire tmp11043;
  wire tmp11044;
  wire tmp11045;
  wire tmp11046;
  wire tmp11047;
  wire tmp11048;
  wire tmp11049;
  wire tmp11050;
  wire tmp11051;
  wire tmp11052;
  wire tmp11053;
  wire tmp11054;
  wire tmp11055;
  wire tmp11056;
  wire tmp11057;
  wire tmp11058;
  wire tmp11059;
  wire tmp11060;
  wire tmp11061;
  wire tmp11062;
  wire tmp11063;
  wire tmp11064;
  wire tmp11065;
  wire tmp11066;
  wire tmp11067;
  wire tmp11068;
  wire tmp11069;
  wire tmp11070;
  wire tmp11071;
  wire tmp11072;
  wire tmp11073;
  wire tmp11074;
  wire tmp11075;
  wire tmp11076;
  wire tmp11077;
  wire tmp11078;
  wire tmp11079;
  wire tmp11080;
  wire tmp11081;
  wire tmp11082;
  wire tmp11083;
  wire tmp11084;
  wire tmp11085;
  wire tmp11086;
  wire tmp11087;
  wire tmp11088;
  wire tmp11089;
  wire tmp11090;
  wire tmp11091;
  wire tmp11092;
  wire tmp11093;
  wire tmp11094;
  wire tmp11095;
  wire tmp11096;
  wire tmp11097;
  wire tmp11098;
  wire tmp11099;
  wire tmp11100;
  wire tmp11101;
  wire tmp11102;
  wire tmp11103;
  wire tmp11104;
  wire tmp11105;
  wire tmp11106;
  wire tmp11107;
  wire tmp11108;
  wire tmp11109;
  wire tmp11110;
  wire tmp11111;
  wire tmp11112;
  wire tmp11113;
  wire tmp11114;
  wire tmp11115;
  wire tmp11116;
  wire tmp11117;
  wire tmp11118;
  wire tmp11119;
  wire tmp11120;
  wire tmp11121;
  wire tmp11122;
  wire tmp11123;
  wire tmp11124;
  wire tmp11125;
  wire tmp11126;
  wire tmp11127;
  wire tmp11128;
  wire tmp11129;
  wire tmp11130;
  wire tmp11131;
  wire tmp11132;
  wire tmp11133;
  wire tmp11134;
  wire tmp11135;
  wire tmp11136;
  wire tmp11137;
  wire tmp11138;
  wire tmp11139;
  wire tmp11140;
  wire tmp11141;
  wire tmp11142;
  wire tmp11143;
  wire tmp11144;
  wire tmp11145;
  wire tmp11146;
  wire tmp11147;
  wire tmp11148;
  wire tmp11149;
  wire tmp11150;
  wire tmp11151;
  wire tmp11152;
  wire tmp11153;
  wire tmp11154;
  wire tmp11155;
  wire tmp11156;
  wire tmp11157;
  wire tmp11158;
  wire tmp11159;
  wire tmp11160;
  wire tmp11161;
  wire tmp11162;
  wire tmp11163;
  wire tmp11164;
  wire tmp11165;
  wire tmp11166;
  wire tmp11167;
  wire tmp11168;
  wire tmp11169;
  wire tmp11170;
  wire tmp11171;
  wire tmp11172;
  wire tmp11173;
  wire tmp11174;
  wire tmp11175;
  wire tmp11176;
  wire tmp11177;
  wire tmp11178;
  wire tmp11179;
  wire tmp11180;
  wire tmp11181;
  wire tmp11182;
  wire tmp11183;
  wire tmp11184;
  wire tmp11185;
  wire tmp11186;
  wire tmp11187;
  wire tmp11188;
  wire tmp11189;
  wire tmp11190;
  wire tmp11191;
  wire tmp11192;
  wire tmp11193;
  wire tmp11194;
  wire tmp11195;
  wire tmp11196;
  wire tmp11197;
  wire tmp11198;
  wire tmp11199;
  wire tmp11200;
  wire tmp11201;
  wire tmp11202;
  wire tmp11203;
  wire tmp11204;
  wire tmp11205;
  wire tmp11206;
  wire tmp11207;
  wire tmp11208;
  wire tmp11209;
  wire tmp11210;
  wire tmp11211;
  wire tmp11212;
  wire tmp11213;
  wire tmp11214;
  wire tmp11215;
  wire tmp11216;
  wire tmp11217;
  wire tmp11218;
  wire tmp11219;
  wire tmp11220;
  wire tmp11221;
  wire tmp11222;
  wire tmp11223;
  wire tmp11224;
  wire tmp11225;
  wire tmp11226;
  wire tmp11227;
  wire tmp11228;
  wire tmp11229;
  wire tmp11230;
  wire tmp11231;
  wire tmp11232;
  wire tmp11233;
  wire tmp11234;
  wire tmp11235;
  wire tmp11236;
  wire tmp11237;
  wire tmp11238;
  wire tmp11239;
  wire tmp11240;
  wire tmp11241;
  wire tmp11242;
  wire tmp11243;
  wire tmp11244;
  wire tmp11245;
  wire tmp11246;
  wire tmp11247;
  wire tmp11248;
  wire tmp11249;
  wire tmp11250;
  wire tmp11251;
  wire tmp11252;
  wire tmp11253;
  wire tmp11254;
  wire tmp11255;
  wire tmp11256;
  wire tmp11257;
  wire tmp11258;
  wire tmp11259;
  wire tmp11260;
  wire tmp11261;
  wire tmp11262;
  wire tmp11263;
  wire tmp11264;
  wire tmp11265;
  wire tmp11266;
  wire tmp11267;
  wire tmp11268;
  wire tmp11269;
  wire tmp11270;
  wire tmp11271;
  wire tmp11272;
  wire tmp11273;
  wire tmp11274;
  wire tmp11275;
  wire tmp11276;
  wire tmp11277;
  wire tmp11278;
  wire tmp11279;
  wire tmp11280;
  wire tmp11281;
  wire tmp11282;
  wire tmp11283;
  wire tmp11284;
  wire tmp11285;
  wire tmp11286;
  wire tmp11287;
  wire tmp11288;
  wire tmp11289;
  wire tmp11290;
  wire tmp11291;
  wire tmp11292;
  wire tmp11293;
  wire tmp11294;
  wire tmp11295;
  wire tmp11296;
  wire tmp11297;
  wire tmp11298;
  wire tmp11299;
  wire tmp11300;
  wire tmp11301;
  wire tmp11302;
  wire tmp11303;
  wire tmp11304;
  wire tmp11305;
  wire tmp11306;
  wire tmp11307;
  wire tmp11308;
  wire tmp11309;
  wire tmp11310;
  wire tmp11311;
  wire tmp11312;
  wire tmp11313;
  wire tmp11314;
  wire tmp11315;
  wire tmp11316;
  wire tmp11317;
  wire tmp11318;
  wire tmp11319;
  wire tmp11320;
  wire tmp11321;
  wire tmp11322;
  wire tmp11323;
  wire tmp11324;
  wire tmp11325;
  wire tmp11326;
  wire tmp11327;
  wire tmp11328;
  wire tmp11329;
  wire tmp11330;
  wire tmp11331;
  wire tmp11332;
  wire tmp11333;
  wire tmp11334;
  wire tmp11335;
  wire tmp11336;
  wire tmp11337;
  wire tmp11338;
  wire tmp11339;
  wire tmp11340;
  wire tmp11341;
  wire tmp11342;
  wire tmp11343;
  wire tmp11344;
  wire tmp11345;
  wire tmp11346;
  wire tmp11347;
  wire tmp11348;
  wire tmp11349;
  wire tmp11350;
  wire tmp11351;
  wire tmp11352;
  wire tmp11353;
  wire tmp11354;
  wire tmp11355;
  wire tmp11356;
  wire tmp11357;
  wire tmp11358;
  wire tmp11359;
  wire tmp11360;
  wire tmp11361;
  wire tmp11362;
  wire tmp11363;
  wire tmp11364;
  wire tmp11365;
  wire tmp11366;
  wire tmp11367;
  wire tmp11368;
  wire tmp11369;
  wire tmp11370;
  wire tmp11371;
  wire tmp11372;
  wire tmp11373;
  wire tmp11374;
  wire tmp11375;
  wire tmp11376;
  wire tmp11377;
  wire tmp11378;
  wire tmp11379;
  wire tmp11380;
  wire tmp11381;
  wire tmp11382;
  wire tmp11383;
  wire tmp11384;
  wire tmp11385;
  wire tmp11386;
  wire tmp11387;
  wire tmp11388;
  wire tmp11389;
  wire tmp11390;
  wire tmp11391;
  wire tmp11392;
  wire tmp11393;
  wire tmp11394;
  wire tmp11395;
  wire tmp11396;
  wire tmp11397;
  wire tmp11398;
  wire tmp11399;
  wire tmp11400;
  wire tmp11401;
  wire tmp11402;
  wire tmp11403;
  wire tmp11404;
  wire tmp11405;
  wire tmp11406;
  wire tmp11407;
  wire tmp11408;
  wire tmp11409;
  wire tmp11410;
  wire tmp11411;
  wire tmp11412;
  wire tmp11413;
  wire tmp11414;
  wire tmp11415;
  wire tmp11416;
  wire tmp11417;
  wire tmp11418;
  wire tmp11419;
  wire tmp11420;
  wire tmp11421;
  wire tmp11422;
  wire tmp11423;
  wire tmp11424;
  wire tmp11425;
  wire tmp11426;
  wire tmp11427;
  wire tmp11428;
  wire tmp11429;
  wire tmp11430;
  wire tmp11431;
  wire tmp11432;
  wire tmp11433;
  wire tmp11434;
  wire tmp11435;
  wire tmp11436;
  wire tmp11437;
  wire tmp11438;
  wire tmp11439;
  wire tmp11440;
  wire tmp11441;
  wire tmp11442;
  wire tmp11443;
  wire tmp11444;
  wire tmp11445;
  wire tmp11446;
  wire tmp11447;
  wire tmp11448;
  wire tmp11449;
  wire tmp11450;
  wire tmp11451;
  wire tmp11452;
  wire tmp11453;
  wire tmp11454;
  wire tmp11455;
  wire tmp11456;
  wire tmp11457;
  wire tmp11458;
  wire tmp11459;
  wire tmp11460;
  wire tmp11461;
  wire tmp11462;
  wire tmp11463;
  wire tmp11464;
  wire tmp11465;
  wire tmp11466;
  wire tmp11467;
  wire tmp11468;
  wire tmp11469;
  wire tmp11470;
  wire tmp11471;
  wire tmp11472;
  wire tmp11473;
  wire tmp11474;
  wire tmp11475;
  wire tmp11476;
  wire tmp11477;
  wire tmp11478;
  wire tmp11479;
  wire tmp11480;
  wire tmp11481;
  wire tmp11482;
  wire tmp11483;
  wire tmp11484;
  wire tmp11485;
  wire tmp11486;
  wire tmp11487;
  wire tmp11488;
  wire tmp11489;
  wire tmp11490;
  wire tmp11491;
  wire tmp11492;
  wire tmp11493;
  wire tmp11494;
  wire tmp11495;
  wire tmp11496;
  wire tmp11497;
  wire tmp11498;
  wire tmp11499;
  wire tmp11500;
  wire tmp11501;
  wire tmp11502;
  wire tmp11503;
  wire tmp11504;
  wire tmp11505;
  wire tmp11506;
  wire tmp11507;
  wire tmp11508;
  wire tmp11509;
  wire tmp11510;
  wire tmp11511;
  wire tmp11512;
  wire tmp11513;
  wire tmp11514;
  wire tmp11515;
  wire tmp11516;
  wire tmp11517;
  wire tmp11518;
  wire tmp11519;
  wire tmp11520;
  wire tmp11521;
  wire tmp11522;
  wire tmp11523;
  wire tmp11524;
  wire tmp11525;
  wire tmp11526;
  wire tmp11527;
  wire tmp11528;
  wire tmp11529;
  wire tmp11530;
  wire tmp11531;
  wire tmp11532;
  wire tmp11533;
  wire tmp11534;
  wire tmp11535;
  wire tmp11536;
  wire tmp11537;
  wire tmp11538;
  wire tmp11539;
  wire tmp11540;
  wire tmp11541;
  wire tmp11542;
  wire tmp11543;
  wire tmp11544;
  wire tmp11545;
  wire tmp11546;
  wire tmp11547;
  wire tmp11548;
  wire tmp11549;
  wire tmp11550;
  wire tmp11551;
  wire tmp11552;
  wire tmp11553;
  wire tmp11554;
  wire tmp11555;
  wire tmp11556;
  wire tmp11557;
  wire tmp11558;
  wire tmp11559;
  wire tmp11560;
  wire tmp11561;
  wire tmp11562;
  wire tmp11563;
  wire tmp11564;
  wire tmp11565;
  wire tmp11566;
  wire tmp11567;
  wire tmp11568;
  wire tmp11569;
  wire tmp11570;
  wire tmp11571;
  wire tmp11572;
  wire tmp11573;
  wire tmp11574;
  wire tmp11575;
  wire tmp11576;
  wire tmp11577;
  wire tmp11578;
  wire tmp11579;
  wire tmp11580;
  wire tmp11581;
  wire tmp11582;
  wire tmp11583;
  wire tmp11584;
  wire tmp11585;
  wire tmp11586;
  wire tmp11587;
  wire tmp11588;
  wire tmp11589;
  wire tmp11590;
  wire tmp11591;
  wire tmp11592;
  wire tmp11593;
  wire tmp11594;
  wire tmp11595;
  wire tmp11596;
  wire tmp11597;
  wire tmp11598;
  wire tmp11599;
  wire tmp11600;
  wire tmp11601;
  wire tmp11602;
  wire tmp11603;
  wire tmp11604;
  wire tmp11605;
  wire tmp11606;
  wire tmp11607;
  wire tmp11608;
  wire tmp11609;
  wire tmp11610;
  wire tmp11611;
  wire tmp11612;
  wire tmp11613;
  wire tmp11614;
  wire tmp11615;
  wire tmp11616;
  wire tmp11617;
  wire tmp11618;
  wire tmp11619;
  wire tmp11620;
  wire tmp11621;
  wire tmp11622;
  wire tmp11623;
  wire tmp11624;
  wire tmp11625;
  wire tmp11626;
  wire tmp11627;
  wire tmp11628;
  wire tmp11629;
  wire tmp11630;
  wire tmp11631;
  wire tmp11632;
  wire tmp11633;
  wire tmp11634;
  wire tmp11635;
  wire tmp11636;
  wire tmp11637;
  wire tmp11638;
  wire tmp11639;
  wire tmp11640;
  wire tmp11641;
  wire tmp11642;
  wire tmp11643;
  wire tmp11644;
  wire tmp11645;
  wire tmp11646;
  wire tmp11647;
  wire tmp11648;
  wire tmp11649;
  wire tmp11650;
  wire tmp11651;
  wire tmp11652;
  wire tmp11653;
  wire tmp11654;
  wire tmp11655;
  wire tmp11656;
  wire tmp11657;
  wire tmp11658;
  wire tmp11659;
  wire tmp11660;
  wire tmp11661;
  wire tmp11662;
  wire tmp11663;
  wire tmp11664;
  wire tmp11665;
  wire tmp11666;
  wire tmp11667;
  wire tmp11668;
  wire tmp11669;
  wire tmp11670;
  wire tmp11671;
  wire tmp11672;
  wire tmp11673;
  wire tmp11674;
  wire tmp11675;
  wire tmp11676;
  wire tmp11677;
  wire tmp11678;
  wire tmp11679;
  wire tmp11680;
  wire tmp11681;
  wire tmp11682;
  wire tmp11683;
  wire tmp11684;
  wire tmp11685;
  wire tmp11686;
  wire tmp11687;
  wire tmp11688;
  wire tmp11689;
  wire tmp11690;
  wire tmp11691;
  wire tmp11692;
  wire tmp11693;
  wire tmp11694;
  wire tmp11695;
  wire tmp11696;
  wire tmp11697;
  wire tmp11698;
  wire tmp11699;
  wire tmp11700;
  wire tmp11701;
  wire tmp11702;
  wire tmp11703;
  wire tmp11704;
  wire tmp11705;
  wire tmp11706;
  wire tmp11707;
  wire tmp11708;
  wire tmp11709;
  wire tmp11710;
  wire tmp11711;
  wire tmp11712;
  wire tmp11713;
  wire tmp11714;
  wire tmp11715;
  wire tmp11716;
  wire tmp11717;
  wire tmp11718;
  wire tmp11719;
  wire tmp11720;
  wire tmp11721;
  wire tmp11722;
  wire tmp11723;
  wire tmp11724;
  wire tmp11725;
  wire tmp11726;
  wire tmp11727;
  wire tmp11728;
  wire tmp11729;
  wire tmp11730;
  wire tmp11731;
  wire tmp11732;
  wire tmp11733;
  wire tmp11734;
  wire tmp11735;
  wire tmp11736;
  wire tmp11737;
  wire tmp11738;
  wire tmp11739;
  wire tmp11740;
  wire tmp11741;
  wire tmp11742;
  wire tmp11743;
  wire tmp11744;
  wire tmp11745;
  wire tmp11746;
  wire tmp11747;
  wire tmp11748;
  wire tmp11749;
  wire tmp11750;
  wire tmp11751;
  wire tmp11752;
  wire tmp11753;
  wire tmp11754;
  wire tmp11755;
  wire tmp11756;
  wire tmp11757;
  wire tmp11758;
  wire tmp11759;
  wire tmp11760;
  wire tmp11761;
  wire tmp11762;
  wire tmp11763;
  wire tmp11764;
  wire tmp11765;
  wire tmp11766;
  wire tmp11767;
  wire tmp11768;
  wire tmp11769;
  wire tmp11770;
  wire tmp11771;
  wire tmp11772;
  wire tmp11773;
  wire tmp11774;
  wire tmp11775;
  wire tmp11776;
  wire tmp11777;
  wire tmp11778;
  wire tmp11779;
  wire tmp11780;
  wire tmp11781;
  wire tmp11782;
  wire tmp11783;
  wire tmp11784;
  wire tmp11785;
  wire tmp11786;
  wire tmp11787;
  wire tmp11788;
  wire tmp11789;
  wire tmp11790;
  wire tmp11791;
  wire tmp11792;
  wire tmp11793;
  wire tmp11794;
  wire tmp11795;
  wire tmp11796;
  wire tmp11797;
  wire tmp11798;
  wire tmp11799;
  wire tmp11800;
  wire tmp11801;
  wire tmp11802;
  wire tmp11803;
  wire tmp11804;
  wire tmp11805;
  wire tmp11806;
  wire tmp11807;
  wire tmp11808;
  wire tmp11809;
  wire tmp11810;
  wire tmp11811;
  wire tmp11812;
  wire tmp11813;
  wire tmp11814;
  wire tmp11815;
  wire tmp11816;
  wire tmp11817;
  wire tmp11818;
  wire tmp11819;
  wire tmp11820;
  wire tmp11821;
  wire tmp11822;
  wire tmp11823;
  wire tmp11824;
  wire tmp11825;
  wire tmp11826;
  wire tmp11827;
  wire tmp11828;
  wire tmp11829;
  wire tmp11830;
  wire tmp11831;
  wire tmp11832;
  wire tmp11833;
  wire tmp11834;
  wire tmp11835;
  wire tmp11836;
  wire tmp11837;
  wire tmp11838;
  wire tmp11839;
  wire tmp11840;
  wire tmp11841;
  wire tmp11842;
  wire tmp11843;
  wire tmp11844;
  wire tmp11845;
  wire tmp11846;
  wire tmp11847;
  wire tmp11848;
  wire tmp11849;
  wire tmp11850;
  wire tmp11851;
  wire tmp11852;
  wire tmp11853;
  wire tmp11854;
  wire tmp11855;
  wire tmp11856;
  wire tmp11857;
  wire tmp11858;
  wire tmp11859;
  wire tmp11860;
  wire tmp11861;
  wire tmp11862;
  wire tmp11863;
  wire tmp11864;
  wire tmp11865;
  wire tmp11866;
  wire tmp11867;
  wire tmp11868;
  wire tmp11869;
  wire tmp11870;
  wire tmp11871;
  wire tmp11872;
  wire tmp11873;
  wire tmp11874;
  wire tmp11875;
  wire tmp11876;
  wire tmp11877;
  wire tmp11878;
  wire tmp11879;
  wire tmp11880;
  wire tmp11881;
  wire tmp11882;
  wire tmp11883;
  wire tmp11884;
  wire tmp11885;
  wire tmp11886;
  wire tmp11887;
  wire tmp11888;
  wire tmp11889;
  wire tmp11890;
  wire tmp11891;
  wire tmp11892;
  wire tmp11893;
  wire tmp11894;
  wire tmp11895;
  wire tmp11896;
  wire tmp11897;
  wire tmp11898;
  wire tmp11899;
  wire tmp11900;
  wire tmp11901;
  wire tmp11902;
  wire tmp11903;
  wire tmp11904;
  wire tmp11905;
  wire tmp11906;
  wire tmp11907;
  wire tmp11908;
  wire tmp11909;
  wire tmp11910;
  wire tmp11911;
  wire tmp11912;
  wire tmp11913;
  wire tmp11914;
  wire tmp11915;
  wire tmp11916;
  wire tmp11917;
  wire tmp11918;
  wire tmp11919;
  wire tmp11920;
  wire tmp11921;
  wire tmp11922;
  wire tmp11923;
  wire tmp11924;
  wire tmp11925;
  wire tmp11926;
  wire tmp11927;
  wire tmp11928;
  wire tmp11929;
  wire tmp11930;
  wire tmp11931;
  wire tmp11932;
  wire tmp11933;
  wire tmp11934;
  wire tmp11935;
  wire tmp11936;
  wire tmp11937;
  wire tmp11938;
  wire tmp11939;
  wire tmp11940;
  wire tmp11941;
  wire tmp11942;
  wire tmp11943;
  wire tmp11944;
  wire tmp11945;
  wire tmp11946;
  wire tmp11947;
  wire tmp11948;
  wire tmp11949;
  wire tmp11950;
  wire tmp11951;
  wire tmp11952;
  wire tmp11953;
  wire tmp11954;
  wire tmp11955;
  wire tmp11956;
  wire tmp11957;
  wire tmp11958;
  wire tmp11959;
  wire tmp11960;
  wire tmp11961;
  wire tmp11962;
  wire tmp11963;
  wire tmp11964;
  wire tmp11965;
  wire tmp11966;
  wire tmp11967;
  wire tmp11968;
  wire tmp11969;
  wire tmp11970;
  wire tmp11971;
  wire tmp11972;
  wire tmp11973;
  wire tmp11974;
  wire tmp11975;
  wire tmp11976;
  wire tmp11977;
  wire tmp11978;
  wire tmp11979;
  wire tmp11980;
  wire tmp11981;
  wire tmp11982;
  wire tmp11983;
  wire tmp11984;
  wire tmp11985;
  wire tmp11986;
  wire tmp11987;
  wire tmp11988;
  wire tmp11989;
  wire tmp11990;
  wire tmp11991;
  wire tmp11992;
  wire tmp11993;
  wire tmp11994;
  wire tmp11995;
  wire tmp11996;
  wire tmp11997;
  wire tmp11998;
  wire tmp11999;
  wire tmp12000;
  wire tmp12001;
  wire tmp12002;
  wire tmp12003;
  wire tmp12004;
  wire tmp12005;
  wire tmp12006;
  wire tmp12007;
  wire tmp12008;
  wire tmp12009;
  wire tmp12010;
  wire tmp12011;
  wire tmp12012;
  wire tmp12013;
  wire tmp12014;
  wire tmp12015;
  wire tmp12016;
  wire tmp12017;
  wire tmp12018;
  wire tmp12019;
  wire tmp12020;
  wire tmp12021;
  wire tmp12022;
  wire tmp12023;
  wire tmp12024;
  wire tmp12025;
  wire tmp12026;
  wire tmp12027;
  wire tmp12028;
  wire tmp12029;
  wire tmp12030;
  wire tmp12031;
  wire tmp12032;
  wire tmp12033;
  wire tmp12034;
  wire tmp12035;
  wire tmp12036;
  wire tmp12037;
  wire tmp12038;
  wire tmp12039;
  wire tmp12040;
  wire tmp12041;
  wire tmp12042;
  wire tmp12043;
  wire tmp12044;
  wire tmp12045;
  wire tmp12046;
  wire tmp12047;
  wire tmp12048;
  wire tmp12049;
  wire tmp12050;
  wire tmp12051;
  wire tmp12052;
  wire tmp12053;
  wire tmp12054;
  wire tmp12055;
  wire tmp12056;
  wire tmp12057;
  wire tmp12058;
  wire tmp12059;
  wire tmp12060;
  wire tmp12061;
  wire tmp12062;
  wire tmp12063;
  wire tmp12064;
  wire tmp12065;
  wire tmp12066;
  wire tmp12067;
  wire tmp12068;
  wire tmp12069;
  wire tmp12070;
  wire tmp12071;
  wire tmp12072;
  wire tmp12073;
  wire tmp12074;
  wire tmp12075;
  wire tmp12076;
  wire tmp12077;
  wire tmp12078;
  wire tmp12079;
  wire tmp12080;
  wire tmp12081;
  wire tmp12082;
  wire tmp12083;
  wire tmp12084;
  wire tmp12085;
  wire tmp12086;
  wire tmp12087;
  wire tmp12088;
  wire tmp12089;
  wire tmp12090;
  wire tmp12091;
  wire tmp12092;
  wire tmp12093;
  wire tmp12094;
  wire tmp12095;
  wire tmp12096;
  wire tmp12097;
  wire tmp12098;
  wire tmp12099;
  wire tmp12100;
  wire tmp12101;
  wire tmp12102;
  wire tmp12103;
  wire tmp12104;
  wire tmp12105;
  wire tmp12106;
  wire tmp12107;
  wire tmp12108;
  wire tmp12109;
  wire tmp12110;
  wire tmp12111;
  wire tmp12112;
  wire tmp12113;
  wire tmp12114;
  wire tmp12115;
  wire tmp12116;
  wire tmp12117;
  wire tmp12118;
  wire tmp12119;
  wire tmp12120;
  wire tmp12121;
  wire tmp12122;
  wire tmp12123;
  wire tmp12124;
  wire tmp12125;
  wire tmp12126;
  wire tmp12127;
  wire tmp12128;
  wire tmp12129;
  wire tmp12130;
  wire tmp12131;
  wire tmp12132;
  wire tmp12133;
  wire tmp12134;
  wire tmp12135;
  wire tmp12136;
  wire tmp12137;
  wire tmp12138;
  wire tmp12139;
  wire tmp12140;
  wire tmp12141;
  wire tmp12142;
  wire tmp12143;
  wire tmp12144;
  wire tmp12145;
  wire tmp12146;
  wire tmp12147;
  wire tmp12148;
  wire tmp12149;
  wire tmp12150;
  wire tmp12151;
  wire tmp12152;
  wire tmp12153;
  wire tmp12154;
  wire tmp12155;
  wire tmp12156;
  wire tmp12157;
  wire tmp12158;
  wire tmp12159;
  wire tmp12160;
  wire tmp12161;
  wire tmp12162;
  wire tmp12163;
  wire tmp12164;
  wire tmp12165;
  wire tmp12166;
  wire tmp12167;
  wire tmp12168;
  wire tmp12169;
  wire tmp12170;
  wire tmp12171;
  wire tmp12172;
  wire tmp12173;
  wire tmp12174;
  wire tmp12175;
  wire tmp12176;
  wire tmp12177;
  wire tmp12178;
  wire tmp12179;
  wire tmp12180;
  wire tmp12181;
  wire tmp12182;
  wire tmp12183;
  wire tmp12184;
  wire tmp12185;
  wire tmp12186;
  wire tmp12187;
  wire tmp12188;
  wire tmp12189;
  wire tmp12190;
  wire tmp12191;
  wire tmp12192;
  wire tmp12193;
  wire tmp12194;
  wire tmp12195;
  wire tmp12196;
  wire tmp12197;
  wire tmp12198;
  wire tmp12199;
  wire tmp12200;
  wire tmp12201;
  wire tmp12202;
  wire tmp12203;
  wire tmp12204;
  wire tmp12205;
  wire tmp12206;
  wire tmp12207;
  wire tmp12208;
  wire tmp12209;
  wire tmp12210;
  wire tmp12211;
  wire tmp12212;
  wire tmp12213;
  wire tmp12214;
  wire tmp12215;
  wire tmp12216;
  wire tmp12217;
  wire tmp12218;
  wire tmp12219;
  wire tmp12220;
  wire tmp12221;
  wire tmp12222;
  wire tmp12223;
  wire tmp12224;
  wire tmp12225;
  wire tmp12226;
  wire tmp12227;
  wire tmp12228;
  wire tmp12229;
  wire tmp12230;
  wire tmp12231;
  wire tmp12232;
  wire tmp12233;
  wire tmp12234;
  wire tmp12235;
  wire tmp12236;
  wire tmp12237;
  wire tmp12238;
  wire tmp12239;
  wire tmp12240;
  wire tmp12241;
  wire tmp12242;
  wire tmp12243;
  wire tmp12244;
  wire tmp12245;
  wire tmp12246;
  wire tmp12247;
  wire tmp12248;
  wire tmp12249;
  wire tmp12250;
  wire tmp12251;
  wire tmp12252;
  wire tmp12253;
  wire tmp12254;
  wire tmp12255;
  wire tmp12256;
  wire tmp12257;
  wire tmp12258;
  wire tmp12259;
  wire tmp12260;
  wire tmp12261;
  wire tmp12262;
  wire tmp12263;
  wire tmp12264;
  wire tmp12265;
  wire tmp12266;
  wire tmp12267;
  wire tmp12268;
  wire tmp12269;
  wire tmp12270;
  wire tmp12271;
  wire tmp12272;
  wire tmp12273;
  wire tmp12274;
  wire tmp12275;
  wire tmp12276;
  wire tmp12277;
  wire tmp12278;
  wire tmp12279;
  wire tmp12280;
  wire tmp12281;
  wire tmp12282;
  wire tmp12283;
  wire tmp12284;
  wire tmp12285;
  wire tmp12286;
  wire tmp12287;
  wire tmp12288;
  wire tmp12289;
  wire tmp12290;
  wire tmp12291;
  wire tmp12292;
  wire tmp12293;
  wire tmp12294;
  wire tmp12295;
  wire tmp12296;
  wire tmp12297;
  wire tmp12298;
  wire tmp12299;
  wire tmp12300;
  wire tmp12301;
  wire tmp12302;
  wire tmp12303;
  wire tmp12304;
  wire tmp12305;
  wire tmp12306;
  wire tmp12307;
  wire tmp12308;
  wire tmp12309;
  wire tmp12310;
  wire tmp12311;
  wire tmp12312;
  wire tmp12313;
  wire tmp12314;
  wire tmp12315;
  wire tmp12316;
  wire tmp12317;
  wire tmp12318;
  wire tmp12319;
  wire tmp12320;
  wire tmp12321;
  wire tmp12322;
  wire tmp12323;
  wire tmp12324;
  wire tmp12325;
  wire tmp12326;
  wire tmp12327;
  wire tmp12328;
  wire tmp12329;
  wire tmp12330;
  wire tmp12331;
  wire tmp12332;
  wire tmp12333;
  wire tmp12334;
  wire tmp12335;
  wire tmp12336;
  wire tmp12337;
  wire tmp12338;
  wire tmp12339;
  wire tmp12340;
  wire tmp12341;
  wire tmp12342;
  wire tmp12343;
  wire tmp12344;
  wire tmp12345;
  wire tmp12346;
  wire tmp12347;
  wire tmp12348;
  wire tmp12349;
  wire tmp12350;
  wire tmp12351;
  wire tmp12352;
  wire tmp12353;
  wire tmp12354;
  wire tmp12355;
  wire tmp12356;
  wire tmp12357;
  wire tmp12358;
  wire tmp12359;
  wire tmp12360;
  wire tmp12361;
  wire tmp12362;
  wire tmp12363;
  wire tmp12364;
  wire tmp12365;
  wire tmp12366;
  wire tmp12367;
  wire tmp12368;
  wire tmp12369;
  wire tmp12370;
  wire tmp12371;
  wire tmp12372;
  wire tmp12373;
  wire tmp12374;
  wire tmp12375;
  wire tmp12376;
  wire tmp12377;
  wire tmp12378;
  wire tmp12379;
  wire tmp12380;
  wire tmp12381;
  wire tmp12382;
  wire tmp12383;
  wire tmp12384;
  wire tmp12385;
  wire tmp12386;
  wire tmp12387;
  wire tmp12388;
  wire tmp12389;
  wire tmp12390;
  wire tmp12391;
  wire tmp12392;
  wire tmp12393;
  wire tmp12394;
  wire tmp12395;
  wire tmp12396;
  wire tmp12397;
  wire tmp12398;
  wire tmp12399;
  wire tmp12400;
  wire tmp12401;
  wire tmp12402;
  wire tmp12403;
  wire tmp12404;
  wire tmp12405;
  wire tmp12406;
  wire tmp12407;
  wire tmp12408;
  wire tmp12409;
  wire tmp12410;
  wire tmp12411;
  wire tmp12412;
  wire tmp12413;
  wire tmp12414;
  wire tmp12415;
  wire tmp12416;
  wire tmp12417;
  wire tmp12418;
  wire tmp12419;
  wire tmp12420;
  wire tmp12421;
  wire tmp12422;
  wire tmp12423;
  wire tmp12424;
  wire tmp12425;
  wire tmp12426;
  wire tmp12427;
  wire tmp12428;
  wire tmp12429;
  wire tmp12430;
  wire tmp12431;
  wire tmp12432;
  wire tmp12433;
  wire tmp12434;
  wire tmp12435;
  wire tmp12436;
  wire tmp12437;
  wire tmp12438;
  wire tmp12439;
  wire tmp12440;
  wire tmp12441;
  wire tmp12442;
  wire tmp12443;
  wire tmp12444;
  wire tmp12445;
  wire tmp12446;
  wire tmp12447;
  wire tmp12448;
  wire tmp12449;
  wire tmp12450;
  wire tmp12451;
  wire tmp12452;
  wire tmp12453;
  wire tmp12454;
  wire tmp12455;
  wire tmp12456;
  wire tmp12457;
  wire tmp12458;
  wire tmp12459;
  wire tmp12460;
  wire tmp12461;
  wire tmp12462;
  wire tmp12463;
  wire tmp12464;
  wire tmp12465;
  wire tmp12466;
  wire tmp12467;
  wire tmp12468;
  wire tmp12469;
  wire tmp12470;
  wire tmp12471;
  wire tmp12472;
  wire tmp12473;
  wire tmp12474;
  wire tmp12475;
  wire tmp12476;
  wire tmp12477;
  wire tmp12478;
  wire tmp12479;
  wire tmp12480;
  wire tmp12481;
  wire tmp12482;
  wire tmp12483;
  wire tmp12484;
  wire tmp12485;
  wire tmp12486;
  wire tmp12487;
  wire tmp12488;
  wire tmp12489;
  wire tmp12490;
  wire tmp12491;
  wire tmp12492;
  wire tmp12493;
  wire tmp12494;
  wire tmp12495;
  wire tmp12496;
  wire tmp12497;
  wire tmp12498;
  wire tmp12499;
  wire tmp12500;
  wire tmp12501;
  wire tmp12502;
  wire tmp12503;
  wire tmp12504;
  wire tmp12505;
  wire tmp12506;
  wire tmp12507;
  wire tmp12508;
  wire tmp12509;
  wire tmp12510;
  wire tmp12511;
  wire tmp12512;
  wire tmp12513;
  wire tmp12514;
  wire tmp12515;
  wire tmp12516;
  wire tmp12517;
  wire tmp12518;
  wire tmp12519;
  wire tmp12520;
  wire tmp12521;
  wire tmp12522;
  wire tmp12523;
  wire tmp12524;
  wire tmp12525;
  wire tmp12526;
  wire tmp12527;
  wire tmp12528;
  wire tmp12529;
  wire tmp12530;
  wire tmp12531;
  wire tmp12532;
  wire tmp12533;
  wire tmp12534;
  wire tmp12535;
  wire tmp12536;
  wire tmp12537;
  wire tmp12538;
  wire tmp12539;
  wire tmp12540;
  wire tmp12541;
  wire tmp12542;
  wire tmp12543;
  wire tmp12544;
  wire tmp12545;
  wire tmp12546;
  wire tmp12547;
  wire tmp12548;
  wire tmp12549;
  wire tmp12550;
  wire tmp12551;
  wire tmp12552;
  wire tmp12553;
  wire tmp12554;
  wire tmp12555;
  wire tmp12556;
  wire tmp12557;
  wire tmp12558;
  wire tmp12559;
  wire tmp12560;
  wire tmp12561;
  wire tmp12562;
  wire tmp12563;
  wire tmp12564;
  wire tmp12565;
  wire tmp12566;
  wire tmp12567;
  wire tmp12568;
  wire tmp12569;
  wire tmp12570;
  wire tmp12571;
  wire tmp12572;
  wire tmp12573;
  wire tmp12574;
  wire tmp12575;
  wire tmp12576;
  wire tmp12577;
  wire tmp12578;
  wire tmp12579;
  wire tmp12580;
  wire tmp12581;
  wire tmp12582;
  wire tmp12583;
  wire tmp12584;
  wire tmp12585;
  wire tmp12586;
  wire tmp12587;
  wire tmp12588;
  wire tmp12589;
  wire tmp12590;
  wire tmp12591;
  wire tmp12592;
  wire tmp12593;
  wire tmp12594;
  wire tmp12595;
  wire tmp12596;
  wire tmp12597;
  wire tmp12598;
  wire tmp12599;
  wire tmp12600;
  wire tmp12601;
  wire tmp12602;
  wire tmp12603;
  wire tmp12604;
  wire tmp12605;
  wire tmp12606;
  wire tmp12607;
  wire tmp12608;
  wire tmp12609;
  wire tmp12610;
  wire tmp12611;
  wire tmp12612;
  wire tmp12613;
  wire tmp12614;
  wire tmp12615;
  wire tmp12616;
  wire tmp12617;
  wire tmp12618;
  wire tmp12619;
  wire tmp12620;
  wire tmp12621;
  wire tmp12622;
  wire tmp12623;
  wire tmp12624;
  wire tmp12625;
  wire tmp12626;
  wire tmp12627;
  wire tmp12628;
  wire tmp12629;
  wire tmp12630;
  wire tmp12631;
  wire tmp12632;
  wire tmp12633;
  wire tmp12634;
  wire tmp12635;
  wire tmp12636;
  wire tmp12637;
  wire tmp12638;
  wire tmp12639;
  wire tmp12640;
  wire tmp12641;
  wire tmp12642;
  wire tmp12643;
  wire tmp12644;
  wire tmp12645;
  wire tmp12646;
  wire tmp12647;
  wire tmp12648;
  wire tmp12649;
  wire tmp12650;
  wire tmp12651;
  wire tmp12652;
  wire tmp12653;
  wire tmp12654;
  wire tmp12655;
  wire tmp12656;
  wire tmp12657;
  wire tmp12658;
  wire tmp12659;
  wire tmp12660;
  wire tmp12661;
  wire tmp12662;
  wire tmp12663;
  wire tmp12664;
  wire tmp12665;
  wire tmp12666;
  wire tmp12667;
  wire tmp12668;
  wire tmp12669;
  wire tmp12670;
  wire tmp12671;
  wire tmp12672;
  wire tmp12673;
  wire tmp12674;
  wire tmp12675;
  wire tmp12676;
  wire tmp12677;
  wire tmp12678;
  wire tmp12679;
  wire tmp12680;
  wire tmp12681;
  wire tmp12682;
  wire tmp12683;
  wire tmp12684;
  wire tmp12685;
  wire tmp12686;
  wire tmp12687;
  wire tmp12688;
  wire tmp12689;
  wire tmp12690;
  wire tmp12691;
  wire tmp12692;
  wire tmp12693;
  wire tmp12694;
  wire tmp12695;
  wire tmp12696;
  wire tmp12697;
  wire tmp12698;
  wire tmp12699;
  wire tmp12700;
  wire tmp12701;
  wire tmp12702;
  wire tmp12703;
  wire tmp12704;
  wire tmp12705;
  wire tmp12706;
  wire tmp12707;
  wire tmp12708;
  wire tmp12709;
  wire tmp12710;
  wire tmp12711;
  wire tmp12712;
  wire tmp12713;
  wire tmp12714;
  wire tmp12715;
  wire tmp12716;
  wire tmp12717;
  wire tmp12718;
  wire tmp12719;
  wire tmp12720;
  wire tmp12721;
  wire tmp12722;
  wire tmp12723;
  wire tmp12724;
  wire tmp12725;
  wire tmp12726;
  wire tmp12727;
  wire tmp12728;
  wire tmp12729;
  wire tmp12730;
  wire tmp12731;
  wire tmp12732;
  wire tmp12733;
  wire tmp12734;
  wire tmp12735;
  wire tmp12736;
  wire tmp12737;
  wire tmp12738;
  wire tmp12739;
  wire tmp12740;
  wire tmp12741;
  wire tmp12742;
  wire tmp12743;
  wire tmp12744;
  wire tmp12745;
  wire tmp12746;
  wire tmp12747;
  wire tmp12748;
  wire tmp12749;
  wire tmp12750;
  wire tmp12751;
  wire tmp12752;
  wire tmp12753;
  wire tmp12754;
  wire tmp12755;
  wire tmp12756;
  wire tmp12757;
  wire tmp12758;
  wire tmp12759;
  wire tmp12760;
  wire tmp12761;
  wire tmp12762;
  wire tmp12763;
  wire tmp12764;
  wire tmp12765;
  wire tmp12766;
  wire tmp12767;
  wire tmp12768;
  wire tmp12769;
  wire tmp12770;
  wire tmp12771;
  wire tmp12772;
  wire tmp12773;
  wire tmp12774;
  wire tmp12775;
  wire tmp12776;
  wire tmp12777;
  wire tmp12778;
  wire tmp12779;
  wire tmp12780;
  wire tmp12781;
  wire tmp12782;
  wire tmp12783;
  wire tmp12784;
  wire tmp12785;
  wire tmp12786;
  wire tmp12787;
  wire tmp12788;
  wire tmp12789;
  wire tmp12790;
  wire tmp12791;
  wire tmp12792;
  wire tmp12793;
  wire tmp12794;
  wire tmp12795;
  wire tmp12796;
  wire tmp12797;
  wire tmp12798;
  wire tmp12799;
  wire tmp12800;
  wire tmp12801;
  wire tmp12802;
  wire tmp12803;
  wire tmp12804;
  wire tmp12805;
  wire tmp12806;
  wire tmp12807;
  wire tmp12808;
  wire tmp12809;
  wire tmp12810;
  wire tmp12811;
  wire tmp12812;
  wire tmp12813;
  wire tmp12814;
  wire tmp12815;
  wire tmp12816;
  wire tmp12817;
  wire tmp12818;
  wire tmp12819;
  wire tmp12820;
  wire tmp12821;
  wire tmp12822;
  wire tmp12823;
  wire tmp12824;
  wire tmp12825;
  wire tmp12826;
  wire tmp12827;
  wire tmp12828;
  wire tmp12829;
  wire tmp12830;
  wire tmp12831;
  wire tmp12832;
  wire tmp12833;
  wire tmp12834;
  wire tmp12835;
  wire tmp12836;
  wire tmp12837;
  wire tmp12838;
  wire tmp12839;
  wire tmp12840;
  wire tmp12841;
  wire tmp12842;
  wire tmp12843;
  wire tmp12844;
  wire tmp12845;
  wire tmp12846;
  wire tmp12847;
  wire tmp12848;
  wire tmp12849;
  wire tmp12850;
  wire tmp12851;
  wire tmp12852;
  wire tmp12853;
  wire tmp12854;
  wire tmp12855;
  wire tmp12856;
  wire tmp12857;
  wire tmp12858;
  wire tmp12859;
  wire tmp12860;
  wire tmp12861;
  wire tmp12862;
  wire tmp12863;
  wire tmp12864;
  wire tmp12865;
  wire tmp12866;
  wire tmp12867;
  wire tmp12868;
  wire tmp12869;
  wire tmp12870;
  wire tmp12871;
  wire tmp12872;
  wire tmp12873;
  wire tmp12874;
  wire tmp12875;
  wire tmp12876;
  wire tmp12877;
  wire tmp12878;
  wire tmp12879;
  wire tmp12880;
  wire tmp12881;
  wire tmp12882;
  wire tmp12883;
  wire tmp12884;
  wire tmp12885;
  wire tmp12886;
  wire tmp12887;
  wire tmp12888;
  wire tmp12889;
  wire tmp12890;
  wire tmp12891;
  wire tmp12892;
  wire tmp12893;
  wire tmp12894;
  wire tmp12895;
  wire tmp12896;
  wire tmp12897;
  wire tmp12898;
  wire tmp12899;
  wire tmp12900;
  wire tmp12901;
  wire tmp12902;
  wire tmp12903;
  wire tmp12904;
  wire tmp12905;
  wire tmp12906;
  wire tmp12907;
  wire tmp12908;
  wire tmp12909;
  wire tmp12910;
  wire tmp12911;
  wire tmp12912;
  wire tmp12913;
  wire tmp12914;
  wire tmp12915;
  wire tmp12916;
  wire tmp12917;
  wire tmp12918;
  wire tmp12919;
  wire tmp12920;
  wire tmp12921;
  wire tmp12922;
  wire tmp12923;
  wire tmp12924;
  wire tmp12925;
  wire tmp12926;
  wire tmp12927;
  wire tmp12928;
  wire tmp12929;
  wire tmp12930;
  wire tmp12931;
  wire tmp12932;
  wire tmp12933;
  wire tmp12934;
  wire tmp12935;
  wire tmp12936;
  wire tmp12937;
  wire tmp12938;
  wire tmp12939;
  wire tmp12940;
  wire tmp12941;
  wire tmp12942;
  wire tmp12943;
  wire tmp12944;
  wire tmp12945;
  wire tmp12946;
  wire tmp12947;
  wire tmp12948;
  wire tmp12949;
  wire tmp12950;
  wire tmp12951;
  wire tmp12952;
  wire tmp12953;
  wire tmp12954;
  wire tmp12955;
  wire tmp12956;
  wire tmp12957;
  wire tmp12958;
  wire tmp12959;
  wire tmp12960;
  wire tmp12961;
  wire tmp12962;
  wire tmp12963;
  wire tmp12964;
  wire tmp12965;
  wire tmp12966;
  wire tmp12967;
  wire tmp12968;
  wire tmp12969;
  wire tmp12970;
  wire tmp12971;
  wire tmp12972;
  wire tmp12973;
  wire tmp12974;
  wire tmp12975;
  wire tmp12976;
  wire tmp12977;
  wire tmp12978;
  wire tmp12979;
  wire tmp12980;
  wire tmp12981;
  wire tmp12982;
  wire tmp12983;
  wire tmp12984;
  wire tmp12985;
  wire tmp12986;
  wire tmp12987;
  wire tmp12988;
  wire tmp12989;
  wire tmp12990;
  wire tmp12991;
  wire tmp12992;
  wire tmp12993;
  wire tmp12994;
  wire tmp12995;
  wire tmp12996;
  wire tmp12997;
  wire tmp12998;
  wire tmp12999;
  wire tmp13000;
  wire tmp13001;
  wire tmp13002;
  wire tmp13003;
  wire tmp13004;
  wire tmp13005;
  wire tmp13006;
  wire tmp13007;
  wire tmp13008;
  wire tmp13009;
  wire tmp13010;
  wire tmp13011;
  wire tmp13012;
  wire tmp13013;
  wire tmp13014;
  wire tmp13015;
  wire tmp13016;
  wire tmp13017;
  wire tmp13018;
  wire tmp13019;
  wire tmp13020;
  wire tmp13021;
  wire tmp13022;
  wire tmp13023;
  wire tmp13024;
  wire tmp13025;
  wire tmp13026;
  wire tmp13027;
  wire tmp13028;
  wire tmp13029;
  wire tmp13030;
  wire tmp13031;
  wire tmp13032;
  wire tmp13033;
  wire tmp13034;
  wire tmp13035;
  wire tmp13036;
  wire tmp13037;
  wire tmp13038;
  wire tmp13039;
  wire tmp13040;
  wire tmp13041;
  wire tmp13042;
  wire tmp13043;
  wire tmp13044;
  wire tmp13045;
  wire tmp13046;
  wire tmp13047;
  wire tmp13048;
  wire tmp13049;
  wire tmp13050;
  wire tmp13051;
  wire tmp13052;
  wire tmp13053;
  wire tmp13054;
  wire tmp13055;
  wire tmp13056;
  wire tmp13057;
  wire tmp13058;
  wire tmp13059;
  wire tmp13060;
  wire tmp13061;
  wire tmp13062;
  wire tmp13063;
  wire tmp13064;
  wire tmp13065;
  wire tmp13066;
  wire tmp13067;
  wire tmp13068;
  wire tmp13069;
  wire tmp13070;
  wire tmp13071;
  wire tmp13072;
  wire tmp13073;
  wire tmp13074;
  wire tmp13075;
  wire tmp13076;
  wire tmp13077;
  wire tmp13078;
  wire tmp13079;
  wire tmp13080;
  wire tmp13081;
  wire tmp13082;
  wire tmp13083;
  wire tmp13084;
  wire tmp13085;
  wire tmp13086;
  wire tmp13087;
  wire tmp13088;
  wire tmp13089;
  wire tmp13090;
  wire tmp13091;
  wire tmp13092;
  wire tmp13093;
  wire tmp13094;
  wire tmp13095;
  wire tmp13096;
  wire tmp13097;
  wire tmp13098;
  wire tmp13099;
  wire tmp13100;
  wire tmp13101;
  wire tmp13102;
  wire tmp13103;
  wire tmp13104;
  wire tmp13105;
  wire tmp13106;
  wire tmp13107;
  wire tmp13108;
  wire tmp13109;
  wire tmp13110;
  wire tmp13111;
  wire tmp13112;
  wire tmp13113;
  wire tmp13114;
  wire tmp13115;
  wire tmp13116;
  wire tmp13117;
  wire tmp13118;
  wire tmp13119;
  wire tmp13120;
  wire tmp13121;
  wire tmp13122;
  wire tmp13123;
  wire tmp13124;
  wire tmp13125;
  wire tmp13126;
  wire tmp13127;
  wire tmp13128;
  wire tmp13129;
  wire tmp13130;
  wire tmp13131;
  wire tmp13132;
  wire tmp13133;
  wire tmp13134;
  wire tmp13135;
  wire tmp13136;
  wire tmp13137;
  wire tmp13138;
  wire tmp13139;
  wire tmp13140;
  wire tmp13141;
  wire tmp13142;
  wire tmp13143;
  wire tmp13144;
  wire tmp13145;
  wire tmp13146;
  wire tmp13147;
  wire tmp13148;
  wire tmp13149;
  wire tmp13150;
  wire tmp13151;
  wire tmp13152;
  wire tmp13153;
  wire tmp13154;
  wire tmp13155;
  wire tmp13156;
  wire tmp13157;
  wire tmp13158;
  wire tmp13159;
  wire tmp13160;
  wire tmp13161;
  wire tmp13162;
  wire tmp13163;
  wire tmp13164;
  wire tmp13165;
  wire tmp13166;
  wire tmp13167;
  wire tmp13168;
  wire tmp13169;
  wire tmp13170;
  wire tmp13171;
  wire tmp13172;
  wire tmp13173;
  wire tmp13174;
  wire tmp13175;
  wire tmp13176;
  wire tmp13177;
  wire tmp13178;
  wire tmp13179;
  wire tmp13180;
  wire tmp13181;
  wire tmp13182;
  wire tmp13183;
  wire tmp13184;
  wire tmp13185;
  wire tmp13186;
  wire tmp13187;
  wire tmp13188;
  wire tmp13189;
  wire tmp13190;
  wire tmp13191;
  wire tmp13192;
  wire tmp13193;
  wire tmp13194;
  wire tmp13195;
  wire tmp13196;
  wire tmp13197;
  wire tmp13198;
  wire tmp13199;
  wire tmp13200;
  wire tmp13201;
  wire tmp13202;
  wire tmp13203;
  wire tmp13204;
  wire tmp13205;
  wire tmp13206;
  wire tmp13207;
  wire tmp13208;
  wire tmp13209;
  wire tmp13210;
  wire tmp13211;
  wire tmp13212;
  wire tmp13213;
  wire tmp13214;
  wire tmp13215;
  wire tmp13216;
  wire tmp13217;
  wire tmp13218;
  wire tmp13219;
  wire tmp13220;
  wire tmp13221;
  wire tmp13222;
  wire tmp13223;
  wire tmp13224;
  wire tmp13225;
  wire tmp13226;
  wire tmp13227;
  wire tmp13228;
  wire tmp13229;
  wire tmp13230;
  wire tmp13231;
  wire tmp13232;
  wire tmp13233;
  wire tmp13234;
  wire tmp13235;
  wire tmp13236;
  wire tmp13237;
  wire tmp13238;
  wire tmp13239;
  wire tmp13240;
  wire tmp13241;
  wire tmp13242;
  wire tmp13243;
  wire tmp13244;
  wire tmp13245;
  wire tmp13246;
  wire tmp13247;
  wire tmp13248;
  wire tmp13249;
  wire tmp13250;
  wire tmp13251;
  wire tmp13252;
  wire tmp13253;
  wire tmp13254;
  wire tmp13255;
  wire tmp13256;
  wire tmp13257;
  wire tmp13258;
  wire tmp13259;
  wire tmp13260;
  wire tmp13261;
  wire tmp13262;
  wire tmp13263;
  wire tmp13264;
  wire tmp13265;
  wire tmp13266;
  wire tmp13267;
  wire tmp13268;
  wire tmp13269;
  wire tmp13270;
  wire tmp13271;
  wire tmp13272;
  wire tmp13273;
  wire tmp13274;
  wire tmp13275;
  wire tmp13276;
  wire tmp13277;
  wire tmp13278;
  wire tmp13279;
  wire tmp13280;
  wire tmp13281;
  wire tmp13282;
  wire tmp13283;
  wire tmp13284;
  wire tmp13285;
  wire tmp13286;
  wire tmp13287;
  wire tmp13288;
  wire tmp13289;
  wire tmp13290;
  wire tmp13291;
  wire tmp13292;
  wire tmp13293;
  wire tmp13294;
  wire tmp13295;
  wire tmp13296;
  wire tmp13297;
  wire tmp13298;
  wire tmp13299;
  wire tmp13300;
  wire tmp13301;
  wire tmp13302;
  wire tmp13303;
  wire tmp13304;
  wire tmp13305;
  wire tmp13306;
  wire tmp13307;
  wire tmp13308;
  wire tmp13309;
  wire tmp13310;
  wire tmp13311;
  wire tmp13312;
  wire tmp13313;
  wire tmp13314;
  wire tmp13315;
  wire tmp13316;
  wire tmp13317;
  wire tmp13318;
  wire tmp13319;
  wire tmp13320;
  wire tmp13321;
  wire tmp13322;
  wire tmp13323;
  wire tmp13324;
  wire tmp13325;
  wire tmp13326;
  wire tmp13327;
  wire tmp13328;
  wire tmp13329;
  wire tmp13330;
  wire tmp13331;
  wire tmp13332;
  wire tmp13333;
  wire tmp13334;
  wire tmp13335;
  wire tmp13336;
  wire tmp13337;
  wire tmp13338;
  wire tmp13339;
  wire tmp13340;
  wire tmp13341;
  wire tmp13342;
  wire tmp13343;
  wire tmp13344;
  wire tmp13345;
  wire tmp13346;
  wire tmp13347;
  wire tmp13348;
  wire tmp13349;
  wire tmp13350;
  wire tmp13351;
  wire tmp13352;
  wire tmp13353;
  wire tmp13354;
  wire tmp13355;
  wire tmp13356;
  wire tmp13357;
  wire tmp13358;
  wire tmp13359;
  wire tmp13360;
  wire tmp13361;
  wire tmp13362;
  wire tmp13363;
  wire tmp13364;
  wire tmp13365;
  wire tmp13366;
  wire tmp13367;
  wire tmp13368;
  wire tmp13369;
  wire tmp13370;
  wire tmp13371;
  wire tmp13372;
  wire tmp13373;
  wire tmp13374;
  wire tmp13375;
  wire tmp13376;
  wire tmp13377;
  wire tmp13378;
  wire tmp13379;
  wire tmp13380;
  wire tmp13381;
  wire tmp13382;
  wire tmp13383;
  wire tmp13384;
  wire tmp13385;
  wire tmp13386;
  wire tmp13387;
  wire tmp13388;
  wire tmp13389;
  wire tmp13390;
  wire tmp13391;
  wire tmp13392;
  wire tmp13393;
  wire tmp13394;
  wire tmp13395;
  wire tmp13396;
  wire tmp13397;
  wire tmp13398;
  wire tmp13399;
  wire tmp13400;
  wire tmp13401;
  wire tmp13402;
  wire tmp13403;
  wire tmp13404;
  wire tmp13405;
  wire tmp13406;
  wire tmp13407;
  wire tmp13408;
  wire tmp13409;
  wire tmp13410;
  wire tmp13411;
  wire tmp13412;
  wire tmp13413;
  wire tmp13414;
  wire tmp13415;
  wire tmp13416;
  wire tmp13417;
  wire tmp13418;
  wire tmp13419;
  wire tmp13420;
  wire tmp13421;
  wire tmp13422;
  wire tmp13423;
  wire tmp13424;
  wire tmp13425;
  wire tmp13426;
  wire tmp13427;
  wire tmp13428;
  wire tmp13429;
  wire tmp13430;
  wire tmp13431;
  wire tmp13432;
  wire tmp13433;
  wire tmp13434;
  wire tmp13435;
  wire tmp13436;
  wire tmp13437;
  wire tmp13438;
  wire tmp13439;
  wire tmp13440;
  wire tmp13441;
  wire tmp13442;
  wire tmp13443;
  wire tmp13444;
  wire tmp13445;
  wire tmp13446;
  wire tmp13447;
  wire tmp13448;
  wire tmp13449;
  wire tmp13450;
  wire tmp13451;
  wire tmp13452;
  wire tmp13453;
  wire tmp13454;
  wire tmp13455;
  wire tmp13456;
  wire tmp13457;
  wire tmp13458;
  wire tmp13459;
  wire tmp13460;
  wire tmp13461;
  wire tmp13462;
  wire tmp13463;
  wire tmp13464;
  wire tmp13465;
  wire tmp13466;
  wire tmp13467;
  wire tmp13468;
  wire tmp13469;
  wire tmp13470;
  wire tmp13471;
  wire tmp13472;
  wire tmp13473;
  wire tmp13474;
  wire tmp13475;
  wire tmp13476;
  wire tmp13477;
  wire tmp13478;
  wire tmp13479;
  wire tmp13480;
  wire tmp13481;
  wire tmp13482;
  wire tmp13483;
  wire tmp13484;
  wire tmp13485;
  wire tmp13486;
  wire tmp13487;
  wire tmp13488;
  wire tmp13489;
  wire tmp13490;
  wire tmp13491;
  wire tmp13492;
  wire tmp13493;
  wire tmp13494;
  wire tmp13495;
  wire tmp13496;
  wire tmp13497;
  wire tmp13498;
  wire tmp13499;
  wire tmp13500;
  wire tmp13501;
  wire tmp13502;
  wire tmp13503;
  wire tmp13504;
  wire tmp13505;
  wire tmp13506;
  wire tmp13507;
  wire tmp13508;
  wire tmp13509;
  wire tmp13510;
  wire tmp13511;
  wire tmp13512;
  wire tmp13513;
  wire tmp13514;
  wire tmp13515;
  wire tmp13516;
  wire tmp13517;
  wire tmp13518;
  wire tmp13519;
  wire tmp13520;
  wire tmp13521;
  wire tmp13522;
  wire tmp13523;
  wire tmp13524;
  wire tmp13525;
  wire tmp13526;
  wire tmp13527;
  wire tmp13528;
  wire tmp13529;
  wire tmp13530;
  wire tmp13531;
  wire tmp13532;
  wire tmp13533;
  wire tmp13534;
  wire tmp13535;
  wire tmp13536;
  wire tmp13537;
  wire tmp13538;
  wire tmp13539;
  wire tmp13540;
  wire tmp13541;
  wire tmp13542;
  wire tmp13543;
  wire tmp13544;
  wire tmp13545;
  wire tmp13546;
  wire tmp13547;
  wire tmp13548;
  wire tmp13549;
  wire tmp13550;
  wire tmp13551;
  wire tmp13552;
  wire tmp13553;
  wire tmp13554;
  wire tmp13555;
  wire tmp13556;
  wire tmp13557;
  wire tmp13558;
  wire tmp13559;
  wire tmp13560;
  wire tmp13561;
  wire tmp13562;
  wire tmp13563;
  wire tmp13564;
  wire tmp13565;
  wire tmp13566;
  wire tmp13567;
  wire tmp13568;
  wire tmp13569;
  wire tmp13570;
  wire tmp13571;
  wire tmp13572;
  wire tmp13573;
  wire tmp13574;
  wire tmp13575;
  wire tmp13576;
  wire tmp13577;
  wire tmp13578;
  wire tmp13579;
  wire tmp13580;
  wire tmp13581;
  wire tmp13582;
  wire tmp13583;
  wire tmp13584;
  wire tmp13585;
  wire tmp13586;
  wire tmp13587;
  wire tmp13588;
  wire tmp13589;
  wire tmp13590;
  wire tmp13591;
  wire tmp13592;
  wire tmp13593;
  wire tmp13594;
  wire tmp13595;
  wire tmp13596;
  wire tmp13597;
  wire tmp13598;
  wire tmp13599;
  wire tmp13600;
  wire tmp13601;
  wire tmp13602;
  wire tmp13603;
  wire tmp13604;
  wire tmp13605;
  wire tmp13606;
  wire tmp13607;
  wire tmp13608;
  wire tmp13609;
  wire tmp13610;
  wire tmp13611;
  wire tmp13612;
  wire tmp13613;
  wire tmp13614;
  wire tmp13615;
  wire tmp13616;
  wire tmp13617;
  wire tmp13618;
  wire tmp13619;
  wire tmp13620;
  wire tmp13621;
  wire tmp13622;
  wire tmp13623;
  wire tmp13624;
  wire tmp13625;
  wire tmp13626;
  wire tmp13627;
  wire tmp13628;
  wire tmp13629;
  wire tmp13630;
  wire tmp13631;
  wire tmp13632;
  wire tmp13633;
  wire tmp13634;
  wire tmp13635;
  wire tmp13636;
  wire tmp13637;
  wire tmp13638;
  wire tmp13639;
  wire tmp13640;
  wire tmp13641;
  wire tmp13642;
  wire tmp13643;
  wire tmp13644;
  wire tmp13645;
  wire tmp13646;
  wire tmp13647;
  wire tmp13648;
  wire tmp13649;
  wire tmp13650;
  wire tmp13651;
  wire tmp13652;
  wire tmp13653;
  wire tmp13654;
  wire tmp13655;
  wire tmp13656;
  wire tmp13657;
  wire tmp13658;
  wire tmp13659;
  wire tmp13660;
  wire tmp13661;
  wire tmp13662;
  wire tmp13663;
  wire tmp13664;
  wire tmp13665;
  wire tmp13666;
  wire tmp13667;
  wire tmp13668;
  wire tmp13669;
  wire tmp13670;
  wire tmp13671;
  wire tmp13672;
  wire tmp13673;
  wire tmp13674;
  wire tmp13675;
  wire tmp13676;
  wire tmp13677;
  wire tmp13678;
  wire tmp13679;
  wire tmp13680;
  wire tmp13681;
  wire tmp13682;
  wire tmp13683;
  wire tmp13684;
  wire tmp13685;
  wire tmp13686;
  wire tmp13687;
  wire tmp13688;
  wire tmp13689;
  wire tmp13690;
  wire tmp13691;
  wire tmp13692;
  wire tmp13693;
  wire tmp13694;
  wire tmp13695;
  wire tmp13696;
  wire tmp13697;
  wire tmp13698;
  wire tmp13699;
  wire tmp13700;
  wire tmp13701;
  wire tmp13702;
  wire tmp13703;
  wire tmp13704;
  wire tmp13705;
  wire tmp13706;
  wire tmp13707;
  wire tmp13708;
  wire tmp13709;
  wire tmp13710;
  wire tmp13711;
  wire tmp13712;
  wire tmp13713;
  wire tmp13714;
  wire tmp13715;
  wire tmp13716;
  wire tmp13717;
  wire tmp13718;
  wire tmp13719;
  wire tmp13720;
  wire tmp13721;
  wire tmp13722;
  wire tmp13723;
  wire tmp13724;
  wire tmp13725;
  wire tmp13726;
  wire tmp13727;
  wire tmp13728;
  wire tmp13729;
  wire tmp13730;
  wire tmp13731;
  wire tmp13732;
  wire tmp13733;
  wire tmp13734;
  wire tmp13735;
  wire tmp13736;
  wire tmp13737;
  wire tmp13738;
  wire tmp13739;
  wire tmp13740;
  wire tmp13741;
  wire tmp13742;
  wire tmp13743;
  wire tmp13744;
  wire tmp13745;
  wire tmp13746;
  wire tmp13747;
  wire tmp13748;
  wire tmp13749;
  wire tmp13750;
  wire tmp13751;
  wire tmp13752;
  wire tmp13753;
  wire tmp13754;
  wire tmp13755;
  wire tmp13756;
  wire tmp13757;
  wire tmp13758;
  wire tmp13759;
  wire tmp13760;
  wire tmp13761;
  wire tmp13762;
  wire tmp13763;
  wire tmp13764;
  wire tmp13765;
  wire tmp13766;
  wire tmp13767;
  wire tmp13768;
  wire tmp13769;
  wire tmp13770;
  wire tmp13771;
  wire tmp13772;
  wire tmp13773;
  wire tmp13774;
  wire tmp13775;
  wire tmp13776;
  wire tmp13777;
  wire tmp13778;
  wire tmp13779;
  wire tmp13780;
  wire tmp13781;
  wire tmp13782;
  wire tmp13783;
  wire tmp13784;
  wire tmp13785;
  wire tmp13786;
  wire tmp13787;
  wire tmp13788;
  wire tmp13789;
  wire tmp13790;
  wire tmp13791;
  wire tmp13792;
  wire tmp13793;
  wire tmp13794;
  wire tmp13795;
  wire tmp13796;
  wire tmp13797;
  wire tmp13798;
  wire tmp13799;
  wire tmp13800;
  wire tmp13801;
  wire tmp13802;
  wire tmp13803;
  wire tmp13804;
  wire tmp13805;
  wire tmp13806;
  wire tmp13807;
  wire tmp13808;
  wire tmp13809;
  wire tmp13810;
  wire tmp13811;
  wire tmp13812;
  wire tmp13813;
  wire tmp13814;
  wire tmp13815;
  wire tmp13816;
  wire tmp13817;
  wire tmp13818;
  wire tmp13819;
  wire tmp13820;
  wire tmp13821;
  wire tmp13822;
  wire tmp13823;
  wire tmp13824;
  wire tmp13825;
  wire tmp13826;
  wire tmp13827;
  wire tmp13828;
  wire tmp13829;
  wire tmp13830;
  wire tmp13831;
  wire tmp13832;
  wire tmp13833;
  wire tmp13834;
  wire tmp13835;
  wire tmp13836;
  wire tmp13837;
  wire tmp13838;
  wire tmp13839;
  wire tmp13840;
  wire tmp13841;
  wire tmp13842;
  wire tmp13843;
  wire tmp13844;
  wire tmp13845;
  wire tmp13846;
  wire tmp13847;
  wire tmp13848;
  wire tmp13849;
  wire tmp13850;
  wire tmp13851;
  wire tmp13852;
  wire tmp13853;
  wire tmp13854;
  wire tmp13855;
  wire tmp13856;
  wire tmp13857;
  wire tmp13858;
  wire tmp13859;
  wire tmp13860;
  wire tmp13861;
  wire tmp13862;
  wire tmp13863;
  wire tmp13864;
  wire tmp13865;
  wire tmp13866;
  wire tmp13867;
  wire tmp13868;
  wire tmp13869;
  wire tmp13870;
  wire tmp13871;
  wire tmp13872;
  wire tmp13873;
  wire tmp13874;
  wire tmp13875;
  wire tmp13876;
  wire tmp13877;
  wire tmp13878;
  wire tmp13879;
  wire tmp13880;
  wire tmp13881;
  wire tmp13882;
  wire tmp13883;
  wire tmp13884;
  wire tmp13885;
  wire tmp13886;
  wire tmp13887;
  wire tmp13888;
  wire tmp13889;
  wire tmp13890;
  wire tmp13891;
  wire tmp13892;
  wire tmp13893;
  wire tmp13894;
  wire tmp13895;
  wire tmp13896;
  wire tmp13897;
  wire tmp13898;
  wire tmp13899;
  wire tmp13900;
  wire tmp13901;
  wire tmp13902;
  wire tmp13903;
  wire tmp13904;
  wire tmp13905;
  wire tmp13906;
  wire tmp13907;
  wire tmp13908;
  wire tmp13909;
  wire tmp13910;
  wire tmp13911;
  wire tmp13912;
  wire tmp13913;
  wire tmp13914;
  wire tmp13915;
  wire tmp13916;
  wire tmp13917;
  wire tmp13918;
  wire tmp13919;
  wire tmp13920;
  wire tmp13921;
  wire tmp13922;
  wire tmp13923;
  wire tmp13924;
  wire tmp13925;
  wire tmp13926;
  wire tmp13927;
  wire tmp13928;
  wire tmp13929;
  wire tmp13930;
  wire tmp13931;
  wire tmp13932;
  wire tmp13933;
  wire tmp13934;
  wire tmp13935;
  wire tmp13936;
  wire tmp13937;
  wire tmp13938;
  wire tmp13939;
  wire tmp13940;
  wire tmp13941;
  wire tmp13942;
  wire tmp13943;
  wire tmp13944;
  wire tmp13945;
  wire tmp13946;
  wire tmp13947;
  wire tmp13948;
  wire tmp13949;
  wire tmp13950;
  wire tmp13951;
  wire tmp13952;
  wire tmp13953;
  wire tmp13954;
  wire tmp13955;
  wire tmp13956;
  wire tmp13957;
  wire tmp13958;
  wire tmp13959;
  wire tmp13960;
  wire tmp13961;
  wire tmp13962;
  wire tmp13963;
  wire tmp13964;
  wire tmp13965;
  wire tmp13966;
  wire tmp13967;
  wire tmp13968;
  wire tmp13969;
  wire tmp13970;
  wire tmp13971;
  wire tmp13972;
  wire tmp13973;
  wire tmp13974;
  wire tmp13975;
  wire tmp13976;
  wire tmp13977;
  wire tmp13978;
  wire tmp13979;
  wire tmp13980;
  wire tmp13981;
  wire tmp13982;
  wire tmp13983;
  wire tmp13984;
  wire tmp13985;
  wire tmp13986;
  wire tmp13987;
  wire tmp13988;
  wire tmp13989;
  wire tmp13990;
  wire tmp13991;
  wire tmp13992;
  wire tmp13993;
  wire tmp13994;
  wire tmp13995;
  wire tmp13996;
  wire tmp13997;
  wire tmp13998;
  wire tmp13999;
  wire tmp14000;
  wire tmp14001;
  wire tmp14002;
  wire tmp14003;
  wire tmp14004;
  wire tmp14005;
  wire tmp14006;
  wire tmp14007;
  wire tmp14008;
  wire tmp14009;
  wire tmp14010;
  wire tmp14011;
  wire tmp14012;
  wire tmp14013;
  wire tmp14014;
  wire tmp14015;
  wire tmp14016;
  wire tmp14017;
  wire tmp14018;
  wire tmp14019;
  wire tmp14020;
  wire tmp14021;
  wire tmp14022;
  wire tmp14023;
  wire tmp14024;
  wire tmp14025;
  wire tmp14026;
  wire tmp14027;
  wire tmp14028;
  wire tmp14029;
  wire tmp14030;
  wire tmp14031;
  wire tmp14032;
  wire tmp14033;
  wire tmp14034;
  wire tmp14035;
  wire tmp14036;
  wire tmp14037;
  wire tmp14038;
  wire tmp14039;
  wire tmp14040;
  wire tmp14041;
  wire tmp14042;
  wire tmp14043;
  wire tmp14044;
  wire tmp14045;
  wire tmp14046;
  wire tmp14047;
  wire tmp14048;
  wire tmp14049;
  wire tmp14050;
  wire tmp14051;
  wire tmp14052;
  wire tmp14053;
  wire tmp14054;
  wire tmp14055;
  wire tmp14056;
  wire tmp14057;
  wire tmp14058;
  wire tmp14059;
  wire tmp14060;
  wire tmp14061;
  wire tmp14062;
  wire tmp14063;
  wire tmp14064;
  wire tmp14065;
  wire tmp14066;
  wire tmp14067;
  wire tmp14068;
  wire tmp14069;
  wire tmp14070;
  wire tmp14071;
  wire tmp14072;
  wire tmp14073;
  wire tmp14074;
  wire tmp14075;
  wire tmp14076;
  wire tmp14077;
  wire tmp14078;
  wire tmp14079;
  wire tmp14080;
  wire tmp14081;
  wire tmp14082;
  wire tmp14083;
  wire tmp14084;
  wire tmp14085;
  wire tmp14086;
  wire tmp14087;
  wire tmp14088;
  wire tmp14089;
  wire tmp14090;
  wire tmp14091;
  wire tmp14092;
  wire tmp14093;
  wire tmp14094;
  wire tmp14095;
  wire tmp14096;
  wire tmp14097;
  wire tmp14098;
  wire tmp14099;
  wire tmp14100;
  wire tmp14101;
  wire tmp14102;
  wire tmp14103;
  wire tmp14104;
  wire tmp14105;
  wire tmp14106;
  wire tmp14107;
  wire tmp14108;
  wire tmp14109;
  wire tmp14110;
  wire tmp14111;
  wire tmp14112;
  wire tmp14113;
  wire tmp14114;
  wire tmp14115;
  wire tmp14116;
  wire tmp14117;
  wire tmp14118;
  wire tmp14119;
  wire tmp14120;
  wire tmp14121;
  wire tmp14122;
  wire tmp14123;
  wire tmp14124;
  wire tmp14125;
  wire tmp14126;
  wire tmp14127;
  wire tmp14128;
  wire tmp14129;
  wire tmp14130;
  wire tmp14131;
  wire tmp14132;
  wire tmp14133;
  wire tmp14134;
  wire tmp14135;
  wire tmp14136;
  wire tmp14137;
  wire tmp14138;
  wire tmp14139;
  wire tmp14140;
  wire tmp14141;
  wire tmp14142;
  wire tmp14143;
  wire tmp14144;
  wire tmp14145;
  wire tmp14146;
  wire tmp14147;
  wire tmp14148;
  wire tmp14149;
  wire tmp14150;
  wire tmp14151;
  wire tmp14152;
  wire tmp14153;
  wire tmp14154;
  wire tmp14155;
  wire tmp14156;
  wire tmp14157;
  wire tmp14158;
  wire tmp14159;
  wire tmp14160;
  wire tmp14161;
  wire tmp14162;
  wire tmp14163;
  wire tmp14164;
  wire tmp14165;
  wire tmp14166;
  wire tmp14167;
  wire tmp14168;
  wire tmp14169;
  wire tmp14170;
  wire tmp14171;
  wire tmp14172;
  wire tmp14173;
  wire tmp14174;
  wire tmp14175;
  wire tmp14176;
  wire tmp14177;
  wire tmp14178;
  wire tmp14179;
  wire tmp14180;
  wire tmp14181;
  wire tmp14182;
  wire tmp14183;
  wire tmp14184;
  wire tmp14185;
  wire tmp14186;
  wire tmp14187;
  wire tmp14188;
  wire tmp14189;
  wire tmp14190;
  wire tmp14191;
  wire tmp14192;
  wire tmp14193;
  wire tmp14194;
  wire tmp14195;
  wire tmp14196;
  wire tmp14197;
  wire tmp14198;
  wire tmp14199;
  wire tmp14200;
  wire tmp14201;
  wire tmp14202;
  wire tmp14203;
  wire tmp14204;
  wire tmp14205;
  wire tmp14206;
  wire tmp14207;
  wire tmp14208;
  wire tmp14209;
  wire tmp14210;
  wire tmp14211;
  wire tmp14212;
  wire tmp14213;
  wire tmp14214;
  wire tmp14215;
  wire tmp14216;
  wire tmp14217;
  wire tmp14218;
  wire tmp14219;
  wire tmp14220;
  wire tmp14221;
  wire tmp14222;
  wire tmp14223;
  wire tmp14224;
  wire tmp14225;
  wire tmp14226;
  wire tmp14227;
  wire tmp14228;
  wire tmp14229;
  wire tmp14230;
  wire tmp14231;
  wire tmp14232;
  wire tmp14233;
  wire tmp14234;
  wire tmp14235;
  wire tmp14236;
  wire tmp14237;
  wire tmp14238;
  wire tmp14239;
  wire tmp14240;
  wire tmp14241;
  wire tmp14242;
  wire tmp14243;
  wire tmp14244;
  wire tmp14245;
  wire tmp14246;
  wire tmp14247;
  wire tmp14248;
  wire tmp14249;
  wire tmp14250;
  wire tmp14251;
  wire tmp14252;
  wire tmp14253;
  wire tmp14254;
  wire tmp14255;
  wire tmp14256;
  wire tmp14257;
  wire tmp14258;
  wire tmp14259;
  wire tmp14260;
  wire tmp14261;
  wire tmp14262;
  wire tmp14263;
  wire tmp14264;
  wire tmp14265;
  wire tmp14266;
  wire tmp14267;
  wire tmp14268;
  wire tmp14269;
  wire tmp14270;
  wire tmp14271;
  wire tmp14272;
  wire tmp14273;
  wire tmp14274;
  wire tmp14275;
  wire tmp14276;
  wire tmp14277;
  wire tmp14278;
  wire tmp14279;
  wire tmp14280;
  wire tmp14281;
  wire tmp14282;
  wire tmp14283;
  wire tmp14284;
  wire tmp14285;
  wire tmp14286;
  wire tmp14287;
  wire tmp14288;
  wire tmp14289;
  wire tmp14290;
  wire tmp14291;
  wire tmp14292;
  wire tmp14293;
  wire tmp14294;
  wire tmp14295;
  wire tmp14296;
  wire tmp14297;
  wire tmp14298;
  wire tmp14299;
  wire tmp14300;
  wire tmp14301;
  wire tmp14302;
  wire tmp14303;
  wire tmp14304;
  wire tmp14305;
  wire tmp14306;
  wire tmp14307;
  wire tmp14308;
  wire tmp14309;
  wire tmp14310;
  wire tmp14311;
  wire tmp14312;
  wire tmp14313;
  wire tmp14314;
  wire tmp14315;
  wire tmp14316;
  wire tmp14317;
  wire tmp14318;
  wire tmp14319;
  wire tmp14320;
  wire tmp14321;
  wire tmp14322;
  wire tmp14323;
  wire tmp14324;
  wire tmp14325;
  wire tmp14326;
  wire tmp14327;
  wire tmp14328;
  wire tmp14329;
  wire tmp14330;
  wire tmp14331;
  wire tmp14332;
  wire tmp14333;
  wire tmp14334;
  wire tmp14335;
  wire tmp14336;
  wire tmp14337;
  wire tmp14338;
  wire tmp14339;
  wire tmp14340;
  wire tmp14341;
  wire tmp14342;
  wire tmp14343;
  wire tmp14344;
  wire tmp14345;
  wire tmp14346;
  wire tmp14347;
  wire tmp14348;
  wire tmp14349;
  wire tmp14350;
  wire tmp14351;
  wire tmp14352;
  wire tmp14353;
  wire tmp14354;
  wire tmp14355;
  wire tmp14356;
  wire tmp14357;
  wire tmp14358;
  wire tmp14359;
  wire tmp14360;
  wire tmp14361;
  wire tmp14362;
  wire tmp14363;
  wire tmp14364;
  wire tmp14365;
  wire tmp14366;
  wire tmp14367;
  wire tmp14368;
  wire tmp14369;
  wire tmp14370;
  wire tmp14371;
  wire tmp14372;
  wire tmp14373;
  wire tmp14374;
  wire tmp14375;
  wire tmp14376;
  wire tmp14377;
  wire tmp14378;
  wire tmp14379;
  wire tmp14380;
  wire tmp14381;
  wire tmp14382;
  wire tmp14383;
  wire tmp14384;
  wire tmp14385;
  wire tmp14386;
  wire tmp14387;
  wire tmp14388;
  wire tmp14389;
  wire tmp14390;
  wire tmp14391;
  wire tmp14392;
  wire tmp14393;
  wire tmp14394;
  wire tmp14395;
  wire tmp14396;
  wire tmp14397;
  wire tmp14398;
  wire tmp14399;
  wire tmp14400;
  wire tmp14401;
  wire tmp14402;
  wire tmp14403;
  wire tmp14404;
  wire tmp14405;
  wire tmp14406;
  wire tmp14407;
  wire tmp14408;
  wire tmp14409;
  wire tmp14410;
  wire tmp14411;
  wire tmp14412;
  wire tmp14413;
  wire tmp14414;
  wire tmp14415;
  wire tmp14416;
  wire tmp14417;
  wire tmp14418;
  wire tmp14419;
  wire tmp14420;
  wire tmp14421;
  wire tmp14422;
  wire tmp14423;
  wire tmp14424;
  wire tmp14425;
  wire tmp14426;
  wire tmp14427;
  wire tmp14428;
  wire tmp14429;
  wire tmp14430;
  wire tmp14431;
  wire tmp14432;
  wire tmp14433;
  wire tmp14434;
  wire tmp14435;
  wire tmp14436;
  wire tmp14437;
  wire tmp14438;
  wire tmp14439;
  wire tmp14440;
  wire tmp14441;
  wire tmp14442;
  wire tmp14443;
  wire tmp14444;
  wire tmp14445;
  wire tmp14446;
  wire tmp14447;
  wire tmp14448;
  wire tmp14449;
  wire tmp14450;
  wire tmp14451;
  wire tmp14452;
  wire tmp14453;
  wire tmp14454;
  wire tmp14455;
  wire tmp14456;
  wire tmp14457;
  wire tmp14458;
  wire tmp14459;
  wire tmp14460;
  wire tmp14461;
  wire tmp14462;
  wire tmp14463;
  wire tmp14464;
  wire tmp14465;
  wire tmp14466;
  wire tmp14467;
  wire tmp14468;
  wire tmp14469;
  wire tmp14470;
  wire tmp14471;
  wire tmp14472;
  wire tmp14473;
  wire tmp14474;
  wire tmp14475;
  wire tmp14476;
  wire tmp14477;
  wire tmp14478;
  wire tmp14479;
  wire tmp14480;
  wire tmp14481;
  wire tmp14482;
  wire tmp14483;
  wire tmp14484;
  wire tmp14485;
  wire tmp14486;
  wire tmp14487;
  wire tmp14488;
  wire tmp14489;
  wire tmp14490;
  wire tmp14491;
  wire tmp14492;
  wire tmp14493;
  wire tmp14494;
  wire tmp14495;
  wire tmp14496;
  wire tmp14497;
  wire tmp14498;
  wire tmp14499;
  wire tmp14500;
  wire tmp14501;
  wire tmp14502;
  wire tmp14503;
  wire tmp14504;
  wire tmp14505;
  wire tmp14506;
  wire tmp14507;
  wire tmp14508;
  wire tmp14509;
  wire tmp14510;
  wire tmp14511;
  wire tmp14512;
  wire tmp14513;
  wire tmp14514;
  wire tmp14515;
  wire tmp14516;
  wire tmp14517;
  wire tmp14518;
  wire tmp14519;
  wire tmp14520;
  wire tmp14521;
  wire tmp14522;
  wire tmp14523;
  wire tmp14524;
  wire tmp14525;
  wire tmp14526;
  wire tmp14527;
  wire tmp14528;
  wire tmp14529;
  wire tmp14530;
  wire tmp14531;
  wire tmp14532;
  wire tmp14533;
  wire tmp14534;
  wire tmp14535;
  wire tmp14536;
  wire tmp14537;
  wire tmp14538;
  wire tmp14539;
  wire tmp14540;
  wire tmp14541;
  wire tmp14542;
  wire tmp14543;
  wire tmp14544;
  wire tmp14545;
  wire tmp14546;
  wire tmp14547;
  wire tmp14548;
  wire tmp14549;
  wire tmp14550;
  wire tmp14551;
  wire tmp14552;
  wire tmp14553;
  wire tmp14554;
  wire tmp14555;
  wire tmp14556;
  wire tmp14557;
  wire tmp14558;
  wire tmp14559;
  wire tmp14560;
  wire tmp14561;
  wire tmp14562;
  wire tmp14563;
  wire tmp14564;
  wire tmp14565;
  wire tmp14566;
  wire tmp14567;
  wire tmp14568;
  wire tmp14569;
  wire tmp14570;
  wire tmp14571;
  wire tmp14572;
  wire tmp14573;
  wire tmp14574;
  wire tmp14575;
  wire tmp14576;
  wire tmp14577;
  wire tmp14578;
  wire tmp14579;
  wire tmp14580;
  wire tmp14581;
  wire tmp14582;
  wire tmp14583;
  wire tmp14584;
  wire tmp14585;
  wire tmp14586;
  wire tmp14587;
  wire tmp14588;
  wire tmp14589;
  wire tmp14590;
  wire tmp14591;
  wire tmp14592;
  wire tmp14593;
  wire tmp14594;
  wire tmp14595;
  wire tmp14596;
  wire tmp14597;
  wire tmp14598;
  wire tmp14599;
  wire tmp14600;
  wire tmp14601;
  wire tmp14602;
  wire tmp14603;
  wire tmp14604;
  wire tmp14605;
  wire tmp14606;
  wire tmp14607;
  wire tmp14608;
  wire tmp14609;
  wire tmp14610;
  wire tmp14611;
  wire tmp14612;
  wire tmp14613;
  wire tmp14614;
  wire tmp14615;
  wire tmp14616;
  wire tmp14617;
  wire tmp14618;
  wire tmp14619;
  wire tmp14620;
  wire tmp14621;
  wire tmp14622;
  wire tmp14623;
  wire tmp14624;
  wire tmp14625;
  wire tmp14626;
  wire tmp14627;
  wire tmp14628;
  wire tmp14629;
  wire tmp14630;
  wire tmp14631;
  wire tmp14632;
  wire tmp14633;
  wire tmp14634;
  wire tmp14635;
  wire tmp14636;
  wire tmp14637;
  wire tmp14638;
  wire tmp14639;
  wire tmp14640;
  wire tmp14641;
  wire tmp14642;
  wire tmp14643;
  wire tmp14644;
  wire tmp14645;
  wire tmp14646;
  wire tmp14647;
  wire tmp14648;
  wire tmp14649;
  wire tmp14650;
  wire tmp14651;
  wire tmp14652;
  wire tmp14653;
  wire tmp14654;
  wire tmp14655;
  wire tmp14656;
  wire tmp14657;
  wire tmp14658;
  wire tmp14659;
  wire tmp14660;
  wire tmp14661;
  wire tmp14662;
  wire tmp14663;
  wire tmp14664;
  wire tmp14665;
  wire tmp14666;
  wire tmp14667;
  wire tmp14668;
  wire tmp14669;
  wire tmp14670;
  wire tmp14671;
  wire tmp14672;
  wire tmp14673;
  wire tmp14674;
  wire tmp14675;
  wire tmp14676;
  wire tmp14677;
  wire tmp14678;
  wire tmp14679;
  wire tmp14680;
  wire tmp14681;
  wire tmp14682;
  wire tmp14683;
  wire tmp14684;
  wire tmp14685;
  wire tmp14686;
  wire tmp14687;
  wire tmp14688;
  wire tmp14689;
  wire tmp14690;
  wire tmp14691;
  wire tmp14692;
  wire tmp14693;
  wire tmp14694;
  wire tmp14695;
  wire tmp14696;
  wire tmp14697;
  wire tmp14698;
  wire tmp14699;
  wire tmp14700;
  wire tmp14701;
  wire tmp14702;
  wire tmp14703;
  wire tmp14704;
  wire tmp14705;
  wire tmp14706;
  wire tmp14707;
  wire tmp14708;
  wire tmp14709;
  wire tmp14710;
  wire tmp14711;
  wire tmp14712;
  wire tmp14713;
  wire tmp14714;
  wire tmp14715;
  wire tmp14716;
  wire tmp14717;
  wire tmp14718;
  wire tmp14719;
  wire tmp14720;
  wire tmp14721;
  wire tmp14722;
  wire tmp14723;
  wire tmp14724;
  wire tmp14725;
  wire tmp14726;
  wire tmp14727;
  wire tmp14728;
  wire tmp14729;
  wire tmp14730;
  wire tmp14731;
  wire tmp14732;
  wire tmp14733;
  wire tmp14734;
  wire tmp14735;
  wire tmp14736;
  wire tmp14737;
  wire tmp14738;
  wire tmp14739;
  wire tmp14740;
  wire tmp14741;
  wire tmp14742;
  wire tmp14743;
  wire tmp14744;
  wire tmp14745;
  wire tmp14746;
  wire tmp14747;
  wire tmp14748;
  wire tmp14749;
  wire tmp14750;
  wire tmp14751;
  wire tmp14752;
  wire tmp14753;
  wire tmp14754;
  wire tmp14755;
  wire tmp14756;
  wire tmp14757;
  wire tmp14758;
  wire tmp14759;
  wire tmp14760;
  wire tmp14761;
  wire tmp14762;
  wire tmp14763;
  wire tmp14764;
  wire tmp14765;
  wire tmp14766;
  wire tmp14767;
  wire tmp14768;
  wire tmp14769;
  wire tmp14770;
  wire tmp14771;
  wire tmp14772;
  wire tmp14773;
  wire tmp14774;
  wire tmp14775;
  wire tmp14776;
  wire tmp14777;
  wire tmp14778;
  wire tmp14779;
  wire tmp14780;
  wire tmp14781;
  wire tmp14782;
  wire tmp14783;
  wire tmp14784;
  wire tmp14785;
  wire tmp14786;
  wire tmp14787;
  wire tmp14788;
  wire tmp14789;
  wire tmp14790;
  wire tmp14791;
  wire tmp14792;
  wire tmp14793;
  wire tmp14794;
  wire tmp14795;
  wire tmp14796;
  wire tmp14797;
  wire tmp14798;
  wire tmp14799;
  wire tmp14800;
  wire tmp14801;
  wire tmp14802;
  wire tmp14803;
  wire tmp14804;
  wire tmp14805;
  wire tmp14806;
  wire tmp14807;
  wire tmp14808;
  wire tmp14809;
  wire tmp14810;
  wire tmp14811;
  wire tmp14812;
  wire tmp14813;
  wire tmp14814;
  wire tmp14815;
  wire tmp14816;
  wire tmp14817;
  wire tmp14818;
  wire tmp14819;
  wire tmp14820;
  wire tmp14821;
  wire tmp14822;
  wire tmp14823;
  wire tmp14824;
  wire tmp14825;
  wire tmp14826;
  wire tmp14827;
  wire tmp14828;
  wire tmp14829;
  wire tmp14830;
  wire tmp14831;
  wire tmp14832;
  wire tmp14833;
  wire tmp14834;
  wire tmp14835;
  wire tmp14836;
  wire tmp14837;
  wire tmp14838;
  wire tmp14839;
  wire tmp14840;
  wire tmp14841;
  wire tmp14842;
  wire tmp14843;
  wire tmp14844;
  wire tmp14845;
  wire tmp14846;
  wire tmp14847;
  wire tmp14848;
  wire tmp14849;
  wire tmp14850;
  wire tmp14851;
  wire tmp14852;
  wire tmp14853;
  wire tmp14854;
  wire tmp14855;
  wire tmp14856;
  wire tmp14857;
  wire tmp14858;
  wire tmp14859;
  wire tmp14860;
  wire tmp14861;
  wire tmp14862;
  wire tmp14863;
  wire tmp14864;
  wire tmp14865;
  wire tmp14866;
  wire tmp14867;
  wire tmp14868;
  wire tmp14869;
  wire tmp14870;
  wire tmp14871;
  wire tmp14872;
  wire tmp14873;
  wire tmp14874;
  wire tmp14875;
  wire tmp14876;
  wire tmp14877;
  wire tmp14878;
  wire tmp14879;
  wire tmp14880;
  wire tmp14881;
  wire tmp14882;
  wire tmp14883;
  wire tmp14884;
  wire tmp14885;
  wire tmp14886;
  wire tmp14887;
  wire tmp14888;
  wire tmp14889;
  wire tmp14890;
  wire tmp14891;
  wire tmp14892;
  wire tmp14893;
  wire tmp14894;
  wire tmp14895;
  wire tmp14896;
  wire tmp14897;
  wire tmp14898;
  wire tmp14899;
  wire tmp14900;
  wire tmp14901;
  wire tmp14902;
  wire tmp14903;
  wire tmp14904;
  wire tmp14905;
  wire tmp14906;
  wire tmp14907;
  wire tmp14908;
  wire tmp14909;
  wire tmp14910;
  wire tmp14911;
  wire tmp14912;
  wire tmp14913;
  wire tmp14914;
  wire tmp14915;
  wire tmp14916;
  wire tmp14917;
  wire tmp14918;
  wire tmp14919;
  wire tmp14920;
  wire tmp14921;
  wire tmp14922;
  wire tmp14923;
  wire tmp14924;
  wire tmp14925;
  wire tmp14926;
  wire tmp14927;
  wire tmp14928;
  wire tmp14929;
  wire tmp14930;
  wire tmp14931;
  wire tmp14932;
  wire tmp14933;
  wire tmp14934;
  wire tmp14935;
  wire tmp14936;
  wire tmp14937;
  wire tmp14938;
  wire tmp14939;
  wire tmp14940;
  wire tmp14941;
  wire tmp14942;
  wire tmp14943;
  wire tmp14944;
  wire tmp14945;
  wire tmp14946;
  wire tmp14947;
  wire tmp14948;
  wire tmp14949;
  wire tmp14950;
  wire tmp14951;
  wire tmp14952;
  wire tmp14953;
  wire tmp14954;
  wire tmp14955;
  wire tmp14956;
  wire tmp14957;
  wire tmp14958;
  wire tmp14959;
  wire tmp14960;
  wire tmp14961;
  wire tmp14962;
  wire tmp14963;
  wire tmp14964;
  wire tmp14965;
  wire tmp14966;
  wire tmp14967;
  wire tmp14968;
  wire tmp14969;
  wire tmp14970;
  wire tmp14971;
  wire tmp14972;
  wire tmp14973;
  wire tmp14974;
  wire tmp14975;
  wire tmp14976;
  wire tmp14977;
  wire tmp14978;
  wire tmp14979;
  wire tmp14980;
  wire tmp14981;
  wire tmp14982;
  wire tmp14983;
  wire tmp14984;
  wire tmp14985;
  wire tmp14986;
  wire tmp14987;
  wire tmp14988;
  wire tmp14989;
  wire tmp14990;
  wire tmp14991;
  wire tmp14992;
  wire tmp14993;
  wire tmp14994;
  wire tmp14995;
  wire tmp14996;
  wire tmp14997;
  wire tmp14998;
  wire tmp14999;
  wire tmp15000;
  wire tmp15001;
  wire tmp15002;
  wire tmp15003;
  wire tmp15004;
  wire tmp15005;
  wire tmp15006;
  wire tmp15007;
  wire tmp15008;
  wire tmp15009;
  wire tmp15010;
  wire tmp15011;
  wire tmp15012;
  wire tmp15013;
  wire tmp15014;
  wire tmp15015;
  wire tmp15016;
  wire tmp15017;
  wire tmp15018;
  wire tmp15019;
  wire tmp15020;
  wire tmp15021;
  wire tmp15022;
  wire tmp15023;
  wire tmp15024;
  wire tmp15025;
  wire tmp15026;
  wire tmp15027;
  wire tmp15028;
  wire tmp15029;
  wire tmp15030;
  wire tmp15031;
  wire tmp15032;
  wire tmp15033;
  wire tmp15034;
  wire tmp15035;
  wire tmp15036;
  wire tmp15037;
  wire tmp15038;
  wire tmp15039;
  wire tmp15040;
  wire tmp15041;
  wire tmp15042;
  wire tmp15043;
  wire tmp15044;
  wire tmp15045;
  wire tmp15046;
  wire tmp15047;
  wire tmp15048;
  wire tmp15049;
  wire tmp15050;
  wire tmp15051;
  wire tmp15052;
  wire tmp15053;
  wire tmp15054;
  wire tmp15055;
  wire tmp15056;
  wire tmp15057;
  wire tmp15058;
  wire tmp15059;
  wire tmp15060;
  wire tmp15061;
  wire tmp15062;
  wire tmp15063;
  wire tmp15064;
  wire tmp15065;
  wire tmp15066;
  wire tmp15067;
  wire tmp15068;
  wire tmp15069;
  wire tmp15070;
  wire tmp15071;
  wire tmp15072;
  wire tmp15073;
  wire tmp15074;
  wire tmp15075;
  wire tmp15076;
  wire tmp15077;
  wire tmp15078;
  wire tmp15079;
  wire tmp15080;
  wire tmp15081;
  wire tmp15082;
  wire tmp15083;
  wire tmp15084;
  wire tmp15085;
  wire tmp15086;
  wire tmp15087;
  wire tmp15088;
  wire tmp15089;
  wire tmp15090;
  wire tmp15091;
  wire tmp15092;
  wire tmp15093;
  wire tmp15094;
  wire tmp15095;
  wire tmp15096;
  wire tmp15097;
  wire tmp15098;
  wire tmp15099;
  wire tmp15100;
  wire tmp15101;
  wire tmp15102;
  wire tmp15103;
  wire tmp15104;
  wire tmp15105;
  wire tmp15106;
  wire tmp15107;
  wire tmp15108;
  wire tmp15109;
  wire tmp15110;
  wire tmp15111;
  wire tmp15112;
  wire tmp15113;
  wire tmp15114;
  wire tmp15115;
  wire tmp15116;
  wire tmp15117;
  wire tmp15118;
  wire tmp15119;
  wire tmp15120;
  wire tmp15121;
  wire tmp15122;
  wire tmp15123;
  wire tmp15124;
  wire tmp15125;
  wire tmp15126;
  wire tmp15127;
  wire tmp15128;
  wire tmp15129;
  wire tmp15130;
  wire tmp15131;
  wire tmp15132;
  wire tmp15133;
  wire tmp15134;
  wire tmp15135;
  wire tmp15136;
  wire tmp15137;
  wire tmp15138;
  wire tmp15139;
  wire tmp15140;
  wire tmp15141;
  wire tmp15142;
  wire tmp15143;
  wire tmp15144;
  wire tmp15145;
  wire tmp15146;
  wire tmp15147;
  wire tmp15148;
  wire tmp15149;
  wire tmp15150;
  wire tmp15151;
  wire tmp15152;
  wire tmp15153;
  wire tmp15154;
  wire tmp15155;
  wire tmp15156;
  wire tmp15157;
  wire tmp15158;
  wire tmp15159;
  wire tmp15160;
  wire tmp15161;
  wire tmp15162;
  wire tmp15163;
  wire tmp15164;
  wire tmp15165;
  wire tmp15166;
  wire tmp15167;
  wire tmp15168;
  wire tmp15169;
  wire tmp15170;
  wire tmp15171;
  wire tmp15172;
  wire tmp15173;
  wire tmp15174;
  wire tmp15175;
  wire tmp15176;
  wire tmp15177;
  wire tmp15178;
  wire tmp15179;
  wire tmp15180;
  wire tmp15181;
  wire tmp15182;
  wire tmp15183;
  wire tmp15184;
  wire tmp15185;
  wire tmp15186;
  wire tmp15187;
  wire tmp15188;
  wire tmp15189;
  wire tmp15190;
  wire tmp15191;
  wire tmp15192;
  wire tmp15193;
  wire tmp15194;
  wire tmp15195;
  wire tmp15196;
  wire tmp15197;
  wire tmp15198;
  wire tmp15199;
  wire tmp15200;
  wire tmp15201;
  wire tmp15202;
  wire tmp15203;
  wire tmp15204;
  wire tmp15205;
  wire tmp15206;
  wire tmp15207;
  wire tmp15208;
  wire tmp15209;
  wire tmp15210;
  wire tmp15211;
  wire tmp15212;
  wire tmp15213;
  wire tmp15214;
  wire tmp15215;
  wire tmp15216;
  wire tmp15217;
  wire tmp15218;
  wire tmp15219;
  wire tmp15220;
  wire tmp15221;
  wire tmp15222;
  wire tmp15223;
  wire tmp15224;
  wire tmp15225;
  wire tmp15226;
  wire tmp15227;
  wire tmp15228;
  wire tmp15229;
  wire tmp15230;
  wire tmp15231;
  wire tmp15232;
  wire tmp15233;
  wire tmp15234;
  wire tmp15235;
  wire tmp15236;
  wire tmp15237;
  wire tmp15238;
  wire tmp15239;
  wire tmp15240;
  wire tmp15241;
  wire tmp15242;
  wire tmp15243;
  wire tmp15244;
  wire tmp15245;
  wire tmp15246;
  wire tmp15247;
  wire tmp15248;
  wire tmp15249;
  wire tmp15250;
  wire tmp15251;
  wire tmp15252;
  wire tmp15253;
  wire tmp15254;
  wire tmp15255;
  wire tmp15256;
  wire tmp15257;
  wire tmp15258;
  wire tmp15259;
  wire tmp15260;
  wire tmp15261;
  wire tmp15262;
  wire tmp15263;
  wire tmp15264;
  wire tmp15265;
  wire tmp15266;
  wire tmp15267;
  wire tmp15268;
  wire tmp15269;
  wire tmp15270;
  wire tmp15271;
  wire tmp15272;
  wire tmp15273;
  wire tmp15274;
  wire tmp15275;
  wire tmp15276;
  wire tmp15277;
  wire tmp15278;
  wire tmp15279;
  wire tmp15280;
  wire tmp15281;
  wire tmp15282;
  wire tmp15283;
  wire tmp15284;
  wire tmp15285;
  wire tmp15286;
  wire tmp15287;
  wire tmp15288;
  wire tmp15289;
  wire tmp15290;
  wire tmp15291;
  wire tmp15292;
  wire tmp15293;
  wire tmp15294;
  wire tmp15295;
  wire tmp15296;
  wire tmp15297;
  wire tmp15298;
  wire tmp15299;
  wire tmp15300;
  wire tmp15301;
  wire tmp15302;
  wire tmp15303;
  wire tmp15304;
  wire tmp15305;
  wire tmp15306;
  wire tmp15307;
  wire tmp15308;
  wire tmp15309;
  wire tmp15310;
  wire tmp15311;
  wire tmp15312;
  wire tmp15313;
  wire tmp15314;
  wire tmp15315;
  wire tmp15316;
  wire tmp15317;
  wire tmp15318;
  wire tmp15319;
  wire tmp15320;
  wire tmp15321;
  wire tmp15322;
  wire tmp15323;
  wire tmp15324;
  wire tmp15325;
  wire tmp15326;
  wire tmp15327;
  wire tmp15328;
  wire tmp15329;
  wire tmp15330;
  wire tmp15331;
  wire tmp15332;
  wire tmp15333;
  wire tmp15334;
  wire tmp15335;
  wire tmp15336;
  wire tmp15337;
  wire tmp15338;
  wire tmp15339;
  wire tmp15340;
  wire tmp15341;
  wire tmp15342;
  wire tmp15343;
  wire tmp15344;
  wire tmp15345;
  wire tmp15346;
  wire tmp15347;
  wire tmp15348;
  wire tmp15349;
  wire tmp15350;
  wire tmp15351;
  wire tmp15352;
  wire tmp15353;
  wire tmp15354;
  wire tmp15355;
  wire tmp15356;
  wire tmp15357;
  wire tmp15358;
  wire tmp15359;
  wire tmp15360;
  wire tmp15361;
  wire tmp15362;
  wire tmp15363;
  wire tmp15364;
  wire tmp15365;
  wire tmp15366;
  wire tmp15367;
  wire tmp15368;
  wire tmp15369;
  wire tmp15370;
  wire tmp15371;
  wire tmp15372;
  wire tmp15373;
  wire tmp15374;
  wire tmp15375;
  wire tmp15376;
  wire tmp15377;
  wire tmp15378;
  wire tmp15379;
  wire tmp15380;
  wire tmp15381;
  wire tmp15382;
  wire tmp15383;
  wire tmp15384;
  wire tmp15385;
  wire tmp15386;
  wire tmp15387;
  wire tmp15388;
  wire tmp15389;
  wire tmp15390;
  wire tmp15391;
  wire tmp15392;
  wire tmp15393;
  wire tmp15394;
  wire tmp15395;
  wire tmp15396;
  wire tmp15397;
  wire tmp15398;
  wire tmp15399;
  wire tmp15400;
  wire tmp15401;
  wire tmp15402;
  wire tmp15403;
  wire tmp15404;
  wire tmp15405;
  wire tmp15406;
  wire tmp15407;
  wire tmp15408;
  wire tmp15409;
  wire tmp15410;
  wire tmp15411;
  wire tmp15412;
  wire tmp15413;
  wire tmp15414;
  wire tmp15415;
  wire tmp15416;
  wire tmp15417;
  wire tmp15418;
  wire tmp15419;
  wire tmp15420;
  wire tmp15421;
  wire tmp15422;
  wire tmp15423;
  wire tmp15424;
  wire tmp15425;
  wire tmp15426;
  wire tmp15427;
  wire tmp15428;
  wire tmp15429;
  wire tmp15430;
  wire tmp15431;
  wire tmp15432;
  wire tmp15433;
  wire tmp15434;
  wire tmp15435;
  wire tmp15436;
  wire tmp15437;
  wire tmp15438;
  wire tmp15439;
  wire tmp15440;
  wire tmp15441;
  wire tmp15442;
  wire tmp15443;
  wire tmp15444;
  wire tmp15445;
  wire tmp15446;
  wire tmp15447;
  wire tmp15448;
  wire tmp15449;
  wire tmp15450;
  wire tmp15451;
  wire tmp15452;
  wire tmp15453;
  wire tmp15454;
  wire tmp15455;
  wire tmp15456;
  wire tmp15457;
  wire tmp15458;
  wire tmp15459;
  wire tmp15460;
  wire tmp15461;
  wire tmp15462;
  wire tmp15463;
  wire tmp15464;
  wire tmp15465;
  wire tmp15466;
  wire tmp15467;
  wire tmp15468;
  wire tmp15469;
  wire tmp15470;
  wire tmp15471;
  wire tmp15472;
  wire tmp15473;
  wire tmp15474;
  wire tmp15475;
  wire tmp15476;
  wire tmp15477;
  wire tmp15478;
  wire tmp15479;
  wire tmp15480;
  wire tmp15481;
  wire tmp15482;
  wire tmp15483;
  wire tmp15484;
  wire tmp15485;
  wire tmp15486;
  wire tmp15487;
  wire tmp15488;
  wire tmp15489;
  wire tmp15490;
  wire tmp15491;
  wire tmp15492;
  wire tmp15493;
  wire tmp15494;
  wire tmp15495;
  wire tmp15496;
  wire tmp15497;
  wire tmp15498;
  wire tmp15499;
  wire tmp15500;
  wire tmp15501;
  wire tmp15502;
  wire tmp15503;
  wire tmp15504;
  wire tmp15505;
  wire tmp15506;
  wire tmp15507;
  wire tmp15508;
  wire tmp15509;
  wire tmp15510;
  wire tmp15511;
  wire tmp15512;
  wire tmp15513;
  wire tmp15514;
  wire tmp15515;
  wire tmp15516;
  wire tmp15517;
  wire tmp15518;
  wire tmp15519;
  wire tmp15520;
  wire tmp15521;
  wire tmp15522;
  wire tmp15523;
  wire tmp15524;
  wire tmp15525;
  wire tmp15526;
  wire tmp15527;
  wire tmp15528;
  wire tmp15529;
  wire tmp15530;
  wire tmp15531;
  wire tmp15532;
  wire tmp15533;
  wire tmp15534;
  wire tmp15535;
  wire tmp15536;
  wire tmp15537;
  wire tmp15538;
  wire tmp15539;
  wire tmp15540;
  wire tmp15541;
  wire tmp15542;
  wire tmp15543;
  wire tmp15544;
  wire tmp15545;
  wire tmp15546;
  wire tmp15547;
  wire tmp15548;
  wire tmp15549;
  wire tmp15550;
  wire tmp15551;
  wire tmp15552;
  wire tmp15553;
  wire tmp15554;
  wire tmp15555;
  wire tmp15556;
  wire tmp15557;
  wire tmp15558;
  wire tmp15559;
  wire tmp15560;
  wire tmp15561;
  wire tmp15562;
  wire tmp15563;
  wire tmp15564;
  wire tmp15565;
  wire tmp15566;
  wire tmp15567;
  wire tmp15568;
  wire tmp15569;
  wire tmp15570;
  wire tmp15571;
  wire tmp15572;
  wire tmp15573;
  wire tmp15574;
  wire tmp15575;
  wire tmp15576;
  wire tmp15577;
  wire tmp15578;
  wire tmp15579;
  wire tmp15580;
  wire tmp15581;
  wire tmp15582;
  wire tmp15583;
  wire tmp15584;
  wire tmp15585;
  wire tmp15586;
  wire tmp15587;
  wire tmp15588;
  wire tmp15589;
  wire tmp15590;
  wire tmp15591;
  wire tmp15592;
  wire tmp15593;
  wire tmp15594;
  wire tmp15595;
  wire tmp15596;
  wire tmp15597;
  wire tmp15598;
  wire tmp15599;
  wire tmp15600;
  wire tmp15601;
  wire tmp15602;
  wire tmp15603;
  wire tmp15604;
  wire tmp15605;
  wire tmp15606;
  wire tmp15607;
  wire tmp15608;
  wire tmp15609;
  wire tmp15610;
  wire tmp15611;
  wire tmp15612;
  wire tmp15613;
  wire tmp15614;
  wire tmp15615;
  wire tmp15616;
  wire tmp15617;
  wire tmp15618;
  wire tmp15619;
  wire tmp15620;
  wire tmp15621;
  wire tmp15622;
  wire tmp15623;
  wire tmp15624;
  wire tmp15625;
  wire tmp15626;
  wire tmp15627;
  wire tmp15628;
  wire tmp15629;
  wire tmp15630;
  wire tmp15631;
  wire tmp15632;
  wire tmp15633;
  wire tmp15634;
  wire tmp15635;
  wire tmp15636;
  wire tmp15637;
  wire tmp15638;
  wire tmp15639;
  wire tmp15640;
  wire tmp15641;
  wire tmp15642;
  wire tmp15643;
  wire tmp15644;
  wire tmp15645;
  wire tmp15646;
  wire tmp15647;
  wire tmp15648;
  wire tmp15649;
  wire tmp15650;
  wire tmp15651;
  wire tmp15652;
  wire tmp15653;
  wire tmp15654;
  wire tmp15655;
  wire tmp15656;
  wire tmp15657;
  wire tmp15658;
  wire tmp15659;
  wire tmp15660;
  wire tmp15661;
  wire tmp15662;
  wire tmp15663;
  wire tmp15664;
  wire tmp15665;
  wire tmp15666;
  wire tmp15667;
  wire tmp15668;
  wire tmp15669;
  wire tmp15670;
  wire tmp15671;
  wire tmp15672;
  wire tmp15673;
  wire tmp15674;
  wire tmp15675;
  wire tmp15676;
  wire tmp15677;
  wire tmp15678;
  wire tmp15679;
  wire tmp15680;
  wire tmp15681;
  wire tmp15682;
  wire tmp15683;
  wire tmp15684;
  wire tmp15685;
  wire tmp15686;
  wire tmp15687;
  wire tmp15688;
  wire tmp15689;
  wire tmp15690;
  wire tmp15691;
  wire tmp15692;
  wire tmp15693;
  wire tmp15694;
  wire tmp15695;
  wire tmp15696;
  wire tmp15697;
  wire tmp15698;
  wire tmp15699;
  wire tmp15700;
  wire tmp15701;
  wire tmp15702;
  wire tmp15703;
  wire tmp15704;
  wire tmp15705;
  wire tmp15706;
  wire tmp15707;
  wire tmp15708;
  wire tmp15709;
  wire tmp15710;
  wire tmp15711;
  wire tmp15712;
  wire tmp15713;
  wire tmp15714;
  wire tmp15715;
  wire tmp15716;
  wire tmp15717;
  wire tmp15718;
  wire tmp15719;
  wire tmp15720;
  wire tmp15721;
  wire tmp15722;
  wire tmp15723;
  wire tmp15724;
  wire tmp15725;
  wire tmp15726;
  wire tmp15727;
  wire tmp15728;
  wire tmp15729;
  wire tmp15730;
  wire tmp15731;
  wire tmp15732;
  wire tmp15733;
  wire tmp15734;
  wire tmp15735;
  wire tmp15736;
  wire tmp15737;
  wire tmp15738;
  wire tmp15739;
  wire tmp15740;
  wire tmp15741;
  wire tmp15742;
  wire tmp15743;
  wire tmp15744;
  wire tmp15745;
  wire tmp15746;
  wire tmp15747;
  wire tmp15748;
  wire tmp15749;
  wire tmp15750;
  wire tmp15751;
  wire tmp15752;
  wire tmp15753;
  wire tmp15754;
  wire tmp15755;
  wire tmp15756;
  wire tmp15757;
  wire tmp15758;
  wire tmp15759;
  wire tmp15760;
  wire tmp15761;
  wire tmp15762;
  wire tmp15763;
  wire tmp15764;
  wire tmp15765;
  wire tmp15766;
  wire tmp15767;
  wire tmp15768;
  wire tmp15769;
  wire tmp15770;
  wire tmp15771;
  wire tmp15772;
  wire tmp15773;
  wire tmp15774;
  wire tmp15775;
  wire tmp15776;
  wire tmp15777;
  wire tmp15778;
  wire tmp15779;
  wire tmp15780;
  wire tmp15781;
  wire tmp15782;
  wire tmp15783;
  wire tmp15784;
  wire tmp15785;
  wire tmp15786;
  wire tmp15787;
  wire tmp15788;
  wire tmp15789;
  wire tmp15790;
  wire tmp15791;
  wire tmp15792;
  wire tmp15793;
  wire tmp15794;
  wire tmp15795;
  wire tmp15796;
  wire tmp15797;
  wire tmp15798;
  wire tmp15799;
  wire tmp15800;
  wire tmp15801;
  wire tmp15802;
  wire tmp15803;
  wire tmp15804;
  wire tmp15805;
  wire tmp15806;
  wire tmp15807;
  wire tmp15808;
  wire tmp15809;
  wire tmp15810;
  wire tmp15811;
  wire tmp15812;
  wire tmp15813;
  wire tmp15814;
  wire tmp15815;
  wire tmp15816;
  wire tmp15817;
  wire tmp15818;
  wire tmp15819;
  wire tmp15820;
  wire tmp15821;
  wire tmp15822;
  wire tmp15823;
  wire tmp15824;
  wire tmp15825;
  wire tmp15826;
  wire tmp15827;
  wire tmp15828;
  wire tmp15829;
  wire tmp15830;
  wire tmp15831;
  wire tmp15832;
  wire tmp15833;
  wire tmp15834;
  wire tmp15835;
  wire tmp15836;
  wire tmp15837;
  wire tmp15838;
  wire tmp15839;
  wire tmp15840;
  wire tmp15841;
  wire tmp15842;
  wire tmp15843;
  wire tmp15844;
  wire tmp15845;
  wire tmp15846;
  wire tmp15847;
  wire tmp15848;
  wire tmp15849;
  wire tmp15850;
  wire tmp15851;
  wire tmp15852;
  wire tmp15853;
  wire tmp15854;
  wire tmp15855;
  wire tmp15856;
  wire tmp15857;
  wire tmp15858;
  wire tmp15859;
  wire tmp15860;
  wire tmp15861;
  wire tmp15862;
  wire tmp15863;
  wire tmp15864;
  wire tmp15865;
  wire tmp15866;
  wire tmp15867;
  wire tmp15868;
  wire tmp15869;
  wire tmp15870;
  wire tmp15871;
  wire tmp15872;
  wire tmp15873;
  wire tmp15874;
  wire tmp15875;
  wire tmp15876;
  wire tmp15877;
  wire tmp15878;
  wire tmp15879;
  wire tmp15880;
  wire tmp15881;
  wire tmp15882;
  wire tmp15883;
  wire tmp15884;
  wire tmp15885;
  wire tmp15886;
  wire tmp15887;
  wire tmp15888;
  wire tmp15889;
  wire tmp15890;
  wire tmp15891;
  wire tmp15892;
  wire tmp15893;
  wire tmp15894;
  wire tmp15895;
  wire tmp15896;
  wire tmp15897;
  wire tmp15898;
  wire tmp15899;
  wire tmp15900;
  wire tmp15901;
  wire tmp15902;
  wire tmp15903;
  wire tmp15904;
  wire tmp15905;
  wire tmp15906;
  wire tmp15907;
  wire tmp15908;
  wire tmp15909;
  wire tmp15910;
  wire tmp15911;
  wire tmp15912;
  wire tmp15913;
  wire tmp15914;
  wire tmp15915;
  wire tmp15916;
  wire tmp15917;
  wire tmp15918;
  wire tmp15919;
  wire tmp15920;
  wire tmp15921;
  wire tmp15922;
  wire tmp15923;
  wire tmp15924;
  wire tmp15925;
  wire tmp15926;
  wire tmp15927;
  wire tmp15928;
  wire tmp15929;
  wire tmp15930;
  wire tmp15931;
  wire tmp15932;
  wire tmp15933;
  wire tmp15934;
  wire tmp15935;
  wire tmp15936;
  wire tmp15937;
  wire tmp15938;
  wire tmp15939;
  wire tmp15940;
  wire tmp15941;
  wire tmp15942;
  wire tmp15943;
  wire tmp15944;
  wire tmp15945;
  wire tmp15946;
  wire tmp15947;
  wire tmp15948;
  wire tmp15949;
  wire tmp15950;
  wire tmp15951;
  wire tmp15952;
  wire tmp15953;
  wire tmp15954;
  wire tmp15955;
  wire tmp15956;
  wire tmp15957;
  wire tmp15958;
  wire tmp15959;
  wire tmp15960;
  wire tmp15961;
  wire tmp15962;
  wire tmp15963;
  wire tmp15964;
  wire tmp15965;
  wire tmp15966;
  wire tmp15967;
  wire tmp15968;
  wire tmp15969;
  wire tmp15970;
  wire tmp15971;
  wire tmp15972;
  wire tmp15973;
  wire tmp15974;
  wire tmp15975;
  wire tmp15976;
  wire tmp15977;
  wire tmp15978;
  wire tmp15979;
  wire tmp15980;
  wire tmp15981;
  wire tmp15982;
  wire tmp15983;
  wire tmp15984;
  wire tmp15985;
  wire tmp15986;
  wire tmp15987;
  wire tmp15988;
  wire tmp15989;
  wire tmp15990;
  wire tmp15991;
  wire tmp15992;
  wire tmp15993;
  wire tmp15994;
  wire tmp15995;
  wire tmp15996;
  wire tmp15997;
  wire tmp15998;
  wire tmp15999;
  wire tmp16000;
  wire tmp16001;
  wire tmp16002;
  wire tmp16003;
  wire tmp16004;
  wire tmp16005;
  wire tmp16006;
  wire tmp16007;
  wire tmp16008;
  wire tmp16009;
  wire tmp16010;
  wire tmp16011;
  wire tmp16012;
  wire tmp16013;
  wire tmp16014;
  wire tmp16015;
  wire tmp16016;
  wire tmp16017;
  wire tmp16018;
  wire tmp16019;
  wire tmp16020;
  wire tmp16021;
  wire tmp16022;
  wire tmp16023;
  wire tmp16024;
  wire tmp16025;
  wire tmp16026;
  wire tmp16027;
  wire tmp16028;
  wire tmp16029;
  wire tmp16030;
  wire tmp16031;
  wire tmp16032;
  wire tmp16033;
  wire tmp16034;
  wire tmp16035;
  wire tmp16036;
  wire tmp16037;
  wire tmp16038;
  wire tmp16039;
  wire tmp16040;
  wire tmp16041;
  wire tmp16042;
  wire tmp16043;
  wire tmp16044;
  wire tmp16045;
  wire tmp16046;
  wire tmp16047;
  wire tmp16048;
  wire tmp16049;
  wire tmp16050;
  wire tmp16051;
  wire tmp16052;
  wire tmp16053;
  wire tmp16054;
  wire tmp16055;
  wire tmp16056;
  wire tmp16057;
  wire tmp16058;
  wire tmp16059;
  wire tmp16060;
  wire tmp16061;
  wire tmp16062;
  wire tmp16063;
  wire tmp16064;
  wire tmp16065;
  wire tmp16066;
  wire tmp16067;
  wire tmp16068;
  wire tmp16069;
  wire tmp16070;
  wire tmp16071;
  wire tmp16072;
  wire tmp16073;
  wire tmp16074;
  wire tmp16075;
  wire tmp16076;
  wire tmp16077;
  wire tmp16078;
  wire tmp16079;
  wire tmp16080;
  wire tmp16081;
  wire tmp16082;
  wire tmp16083;
  wire tmp16084;
  wire tmp16085;
  wire tmp16086;
  wire tmp16087;
  wire tmp16088;
  wire tmp16089;
  wire tmp16090;
  wire tmp16091;
  wire tmp16092;
  wire tmp16093;
  wire tmp16094;
  wire tmp16095;
  wire tmp16096;
  wire tmp16097;
  wire tmp16098;
  wire tmp16099;
  wire tmp16100;
  wire tmp16101;
  wire tmp16102;
  wire tmp16103;
  wire tmp16104;
  wire tmp16105;
  wire tmp16106;
  wire tmp16107;
  wire tmp16108;
  wire tmp16109;
  wire tmp16110;
  wire tmp16111;
  wire tmp16112;
  wire tmp16113;
  wire tmp16114;
  wire tmp16115;
  wire tmp16116;
  wire tmp16117;
  wire tmp16118;
  wire tmp16119;
  wire tmp16120;
  wire tmp16121;
  wire tmp16122;
  wire tmp16123;
  wire tmp16124;
  wire tmp16125;
  wire tmp16126;
  wire tmp16127;
  wire tmp16128;
  wire tmp16129;
  wire tmp16130;
  wire tmp16131;
  wire tmp16132;
  wire tmp16133;
  wire tmp16134;
  wire tmp16135;
  wire tmp16136;
  wire tmp16137;
  wire tmp16138;
  wire tmp16139;
  wire tmp16140;
  wire tmp16141;
  wire tmp16142;
  wire tmp16143;
  wire tmp16144;
  wire tmp16145;
  wire tmp16146;
  wire tmp16147;
  wire tmp16148;
  wire tmp16149;
  wire tmp16150;
  wire tmp16151;
  wire tmp16152;
  wire tmp16153;
  wire tmp16154;
  wire tmp16155;
  wire tmp16156;
  wire tmp16157;
  wire tmp16158;
  wire tmp16159;
  wire tmp16160;
  wire tmp16161;
  wire tmp16162;
  wire tmp16163;
  wire tmp16164;
  wire tmp16165;
  wire tmp16166;
  wire tmp16167;
  wire tmp16168;
  wire tmp16169;
  wire tmp16170;
  wire tmp16171;
  wire tmp16172;
  wire tmp16173;
  wire tmp16174;
  wire tmp16175;
  wire tmp16176;
  wire tmp16177;
  wire tmp16178;
  wire tmp16179;
  wire tmp16180;
  wire tmp16181;
  wire tmp16182;
  wire tmp16183;
  wire tmp16184;
  wire tmp16185;
  wire tmp16186;
  wire tmp16187;
  wire tmp16188;
  wire tmp16189;
  wire tmp16190;
  wire tmp16191;
  wire tmp16192;
  wire tmp16193;
  wire tmp16194;
  wire tmp16195;
  wire tmp16196;
  wire tmp16197;
  wire tmp16198;
  wire tmp16199;
  wire tmp16200;
  wire tmp16201;
  wire tmp16202;
  wire tmp16203;
  wire tmp16204;
  wire tmp16205;
  wire tmp16206;
  wire tmp16207;
  wire tmp16208;
  wire tmp16209;
  wire tmp16210;
  wire tmp16211;
  wire tmp16212;
  wire tmp16213;
  wire tmp16214;
  wire tmp16215;
  wire tmp16216;
  wire tmp16217;
  wire tmp16218;
  wire tmp16219;
  wire tmp16220;
  wire tmp16221;
  wire tmp16222;
  wire tmp16223;
  wire tmp16224;
  wire tmp16225;
  wire tmp16226;
  wire tmp16227;
  wire tmp16228;
  wire tmp16229;
  wire tmp16230;
  wire tmp16231;
  wire tmp16232;
  wire tmp16233;
  wire tmp16234;
  wire tmp16235;
  wire tmp16236;
  wire tmp16237;
  wire tmp16238;
  wire tmp16239;
  wire tmp16240;
  wire tmp16241;
  wire tmp16242;
  wire tmp16243;
  wire tmp16244;
  wire tmp16245;
  wire tmp16246;
  wire tmp16247;
  wire tmp16248;
  wire tmp16249;
  wire tmp16250;
  wire tmp16251;
  wire tmp16252;
  wire tmp16253;
  wire tmp16254;
  wire tmp16255;
  wire tmp16256;
  wire tmp16257;
  wire tmp16258;
  wire tmp16259;
  wire tmp16260;
  wire tmp16261;
  wire tmp16262;
  wire tmp16263;
  wire tmp16264;
  wire tmp16265;
  wire tmp16266;
  wire tmp16267;
  wire tmp16268;
  wire tmp16269;
  wire tmp16270;
  wire tmp16271;
  wire tmp16272;
  wire tmp16273;
  wire tmp16274;
  wire tmp16275;
  wire tmp16276;
  wire tmp16277;
  wire tmp16278;
  wire tmp16279;
  wire tmp16280;
  wire tmp16281;
  wire tmp16282;
  wire tmp16283;
  wire tmp16284;
  wire tmp16285;
  wire tmp16286;
  wire tmp16287;
  wire tmp16288;
  wire tmp16289;
  wire tmp16290;
  wire tmp16291;
  wire tmp16292;
  wire tmp16293;
  wire tmp16294;
  wire tmp16295;
  wire tmp16296;
  wire tmp16297;
  wire tmp16298;
  wire tmp16299;
  wire tmp16300;
  wire tmp16301;
  wire tmp16302;
  wire tmp16303;
  wire tmp16304;
  wire tmp16305;
  wire tmp16306;
  wire tmp16307;
  wire tmp16308;
  wire tmp16309;
  wire tmp16310;
  wire tmp16311;
  wire tmp16312;
  wire tmp16313;
  wire tmp16314;
  wire tmp16315;
  wire tmp16316;
  wire tmp16317;
  wire tmp16318;
  wire tmp16319;
  wire tmp16320;
  wire tmp16321;
  wire tmp16322;
  wire tmp16323;
  wire tmp16324;
  wire tmp16325;
  wire tmp16326;
  wire tmp16327;
  wire tmp16328;
  wire tmp16329;
  wire tmp16330;
  wire tmp16331;
  wire tmp16332;
  wire tmp16333;
  wire tmp16334;
  wire tmp16335;
  wire tmp16336;
  wire tmp16337;
  wire tmp16338;
  wire tmp16339;
  wire tmp16340;
  wire tmp16341;
  wire tmp16342;
  wire tmp16343;
  wire tmp16344;
  wire tmp16345;
  wire tmp16346;
  wire tmp16347;
  wire tmp16348;
  wire tmp16349;
  wire tmp16350;
  wire tmp16351;
  wire tmp16352;
  wire tmp16353;
  wire tmp16354;
  wire tmp16355;
  wire tmp16356;
  wire tmp16357;
  wire tmp16358;
  wire tmp16359;
  wire tmp16360;
  wire tmp16361;
  wire tmp16362;
  wire tmp16363;
  wire tmp16364;
  wire tmp16365;
  wire tmp16366;
  wire tmp16367;
  wire tmp16368;
  wire tmp16369;
  wire tmp16370;
  wire tmp16371;
  wire tmp16372;
  wire tmp16373;
  wire tmp16374;
  wire tmp16375;
  wire tmp16376;
  wire tmp16377;
  wire tmp16378;
  wire tmp16379;
  wire tmp16380;
  wire tmp16381;
  wire tmp16382;
  wire tmp16383;
  wire tmp16384;
  wire tmp16385;
  wire tmp16386;
  wire tmp16387;
  wire tmp16388;
  wire tmp16389;
  wire tmp16390;
  wire tmp16391;
  wire tmp16392;
  wire tmp16393;
  wire tmp16394;
  wire tmp16395;
  wire tmp16396;
  wire tmp16397;
  wire tmp16398;
  wire tmp16399;
  wire tmp16400;
  wire tmp16401;
  wire tmp16402;
  wire tmp16403;
  wire tmp16404;
  wire tmp16405;
  wire tmp16406;
  wire tmp16407;
  wire tmp16408;
  wire tmp16409;
  wire tmp16410;
  wire tmp16411;
  wire tmp16412;
  wire tmp16413;
  wire tmp16414;
  wire tmp16415;
  wire tmp16416;
  wire tmp16417;
  wire tmp16418;
  wire tmp16419;
  wire tmp16420;
  wire tmp16421;
  wire tmp16422;
  wire tmp16423;
  wire tmp16424;
  wire tmp16425;
  wire tmp16426;
  wire tmp16427;
  wire tmp16428;
  wire tmp16429;
  wire tmp16430;
  wire tmp16431;
  wire tmp16432;
  wire tmp16433;
  wire tmp16434;
  wire tmp16435;
  wire tmp16436;
  wire tmp16437;
  wire tmp16438;
  wire tmp16439;
  wire tmp16440;
  wire tmp16441;
  wire tmp16442;
  wire tmp16443;
  wire tmp16444;
  wire tmp16445;
  wire tmp16446;
  wire tmp16447;
  wire tmp16448;
  wire tmp16449;
  wire tmp16450;
  wire tmp16451;
  wire tmp16452;
  wire tmp16453;
  wire tmp16454;
  wire tmp16455;
  wire tmp16456;
  wire tmp16457;
  wire tmp16458;
  wire tmp16459;
  wire tmp16460;
  wire tmp16461;
  wire tmp16462;
  wire tmp16463;
  wire tmp16464;
  wire tmp16465;
  wire tmp16466;
  wire tmp16467;
  wire tmp16468;
  wire tmp16469;
  wire tmp16470;
  wire tmp16471;
  wire tmp16472;
  wire tmp16473;
  wire tmp16474;
  wire tmp16475;
  wire tmp16476;
  wire tmp16477;
  wire tmp16478;
  wire tmp16479;
  wire tmp16480;
  wire tmp16481;
  wire tmp16482;
  wire tmp16483;
  wire tmp16484;
  wire tmp16485;
  wire tmp16486;
  wire tmp16487;
  wire tmp16488;
  wire tmp16489;
  wire tmp16490;
  wire tmp16491;
  wire tmp16492;
  wire tmp16493;
  wire tmp16494;
  wire tmp16495;
  wire tmp16496;
  wire tmp16497;
  wire tmp16498;
  wire tmp16499;
  wire tmp16500;
  wire tmp16501;
  wire tmp16502;
  wire tmp16503;
  wire tmp16504;
  wire tmp16505;
  wire tmp16506;
  wire tmp16507;
  wire tmp16508;
  wire tmp16509;
  wire tmp16510;
  wire tmp16511;
  wire tmp16512;
  wire tmp16513;
  wire tmp16514;
  wire tmp16515;
  wire tmp16516;
  wire tmp16517;
  wire tmp16518;
  wire tmp16519;
  wire tmp16520;
  wire tmp16521;
  wire tmp16522;
  wire tmp16523;
  wire tmp16524;
  wire tmp16525;
  wire tmp16526;
  wire tmp16527;
  wire tmp16528;
  wire tmp16529;
  wire tmp16530;
  wire tmp16531;
  wire tmp16532;
  wire tmp16533;
  wire tmp16534;
  wire tmp16535;
  wire tmp16536;
  wire tmp16537;
  wire tmp16538;
  wire tmp16539;
  wire tmp16540;
  wire tmp16541;
  wire tmp16542;
  wire tmp16543;
  wire tmp16544;
  wire tmp16545;
  wire tmp16546;
  wire tmp16547;
  wire tmp16548;
  wire tmp16549;
  wire tmp16550;
  wire tmp16551;
  wire tmp16552;
  wire tmp16553;
  wire tmp16554;
  wire tmp16555;
  wire tmp16556;
  wire tmp16557;
  wire tmp16558;
  wire tmp16559;
  wire tmp16560;
  wire tmp16561;
  wire tmp16562;
  wire tmp16563;
  wire tmp16564;
  wire tmp16565;
  wire tmp16566;
  wire tmp16567;
  wire tmp16568;
  wire tmp16569;
  wire tmp16570;
  wire tmp16571;
  wire tmp16572;
  wire tmp16573;
  wire tmp16574;
  wire tmp16575;
  wire tmp16576;
  wire tmp16577;
  wire tmp16578;
  wire tmp16579;
  wire tmp16580;
  wire tmp16581;
  wire tmp16582;
  wire tmp16583;
  wire tmp16584;
  wire tmp16585;
  wire tmp16586;
  wire tmp16587;
  wire tmp16588;
  wire tmp16589;
  wire tmp16590;
  wire tmp16591;
  wire tmp16592;
  wire tmp16593;
  wire tmp16594;
  wire tmp16595;
  wire tmp16596;
  wire tmp16597;
  wire tmp16598;
  wire tmp16599;
  wire tmp16600;
  wire tmp16601;
  wire tmp16602;
  wire tmp16603;
  wire tmp16604;
  wire tmp16605;
  wire tmp16606;
  wire tmp16607;
  wire tmp16608;
  wire tmp16609;
  wire tmp16610;
  wire tmp16611;
  wire tmp16612;
  wire tmp16613;
  wire tmp16614;
  wire tmp16615;
  wire tmp16616;
  wire tmp16617;
  wire tmp16618;
  wire tmp16619;
  wire tmp16620;
  wire tmp16621;
  wire tmp16622;
  wire tmp16623;
  wire tmp16624;
  wire tmp16625;
  wire tmp16626;
  wire tmp16627;
  wire tmp16628;
  wire tmp16629;
  wire tmp16630;
  wire tmp16631;
  wire tmp16632;
  wire tmp16633;
  wire tmp16634;
  wire tmp16635;
  wire tmp16636;
  wire tmp16637;
  wire tmp16638;
  wire tmp16639;
  wire tmp16640;
  wire tmp16641;
  wire tmp16642;
  wire tmp16643;
  wire tmp16644;
  wire tmp16645;
  wire tmp16646;
  wire tmp16647;
  wire tmp16648;
  wire tmp16649;
  wire tmp16650;
  wire tmp16651;
  wire tmp16652;
  wire tmp16653;
  wire tmp16654;
  wire tmp16655;
  wire tmp16656;
  wire tmp16657;
  wire tmp16658;
  wire tmp16659;
  wire tmp16660;
  wire tmp16661;
  wire tmp16662;
  wire tmp16663;
  wire tmp16664;
  wire tmp16665;
  wire tmp16666;
  wire tmp16667;
  wire tmp16668;
  wire tmp16669;
  wire tmp16670;
  wire tmp16671;
  wire tmp16672;
  wire tmp16673;
  wire tmp16674;
  wire tmp16675;
  wire tmp16676;
  wire tmp16677;
  wire tmp16678;
  wire tmp16679;
  wire tmp16680;
  wire tmp16681;
  wire tmp16682;
  wire tmp16683;
  wire tmp16684;
  wire tmp16685;
  wire tmp16686;
  wire tmp16687;
  wire tmp16688;
  wire tmp16689;
  wire tmp16690;
  wire tmp16691;
  wire tmp16692;
  wire tmp16693;
  wire tmp16694;
  wire tmp16695;
  wire tmp16696;
  wire tmp16697;
  wire tmp16698;
  wire tmp16699;
  wire tmp16700;
  wire tmp16701;
  wire tmp16702;
  wire tmp16703;
  wire tmp16704;
  wire tmp16705;
  wire tmp16706;
  wire tmp16707;
  wire tmp16708;
  wire tmp16709;
  wire tmp16710;
  wire tmp16711;
  wire tmp16712;
  wire tmp16713;
  wire tmp16714;
  wire tmp16715;
  wire tmp16716;
  wire tmp16717;
  wire tmp16718;
  wire tmp16719;
  wire tmp16720;
  wire tmp16721;
  wire tmp16722;
  wire tmp16723;
  wire tmp16724;
  wire tmp16725;
  wire tmp16726;
  wire tmp16727;
  wire tmp16728;
  wire tmp16729;
  wire tmp16730;
  wire tmp16731;
  wire tmp16732;
  wire tmp16733;
  wire tmp16734;
  wire tmp16735;
  wire tmp16736;
  wire tmp16737;
  wire tmp16738;
  wire tmp16739;
  wire tmp16740;
  wire tmp16741;
  wire tmp16742;
  wire tmp16743;
  wire tmp16744;
  wire tmp16745;
  wire tmp16746;
  wire tmp16747;
  wire tmp16748;
  wire tmp16749;
  wire tmp16750;
  wire tmp16751;
  wire tmp16752;
  wire tmp16753;
  wire tmp16754;
  wire tmp16755;
  wire tmp16756;
  wire tmp16757;
  wire tmp16758;
  wire tmp16759;
  wire tmp16760;
  wire tmp16761;
  wire tmp16762;
  wire tmp16763;
  wire tmp16764;
  wire tmp16765;
  wire tmp16766;
  wire tmp16767;
  wire tmp16768;
  wire tmp16769;
  wire tmp16770;
  wire tmp16771;
  wire tmp16772;
  wire tmp16773;
  wire tmp16774;
  wire tmp16775;
  wire tmp16776;
  wire tmp16777;
  wire tmp16778;
  wire tmp16779;
  wire tmp16780;
  wire tmp16781;
  wire tmp16782;
  wire tmp16783;
  wire tmp16784;
  wire tmp16785;
  wire tmp16786;
  wire tmp16787;
  wire tmp16788;
  wire tmp16789;
  wire tmp16790;
  wire tmp16791;
  wire tmp16792;
  wire tmp16793;
  wire tmp16794;
  wire tmp16795;
  wire tmp16796;
  wire tmp16797;
  wire tmp16798;
  wire tmp16799;
  wire tmp16800;
  wire tmp16801;
  wire tmp16802;
  wire tmp16803;
  wire tmp16804;
  wire tmp16805;
  wire tmp16806;
  wire tmp16807;
  wire tmp16808;
  wire tmp16809;
  wire tmp16810;
  wire tmp16811;
  wire tmp16812;
  wire tmp16813;
  wire tmp16814;
  wire tmp16815;
  wire tmp16816;
  wire tmp16817;
  wire tmp16818;
  wire tmp16819;
  wire tmp16820;
  wire tmp16821;
  wire tmp16822;
  wire tmp16823;
  wire tmp16824;
  wire tmp16825;
  wire tmp16826;
  wire tmp16827;
  wire tmp16828;
  wire tmp16829;
  wire tmp16830;
  wire tmp16831;
  wire tmp16832;
  wire tmp16833;
  wire tmp16834;
  wire tmp16835;
  wire tmp16836;
  wire tmp16837;
  wire tmp16838;
  wire tmp16839;
  wire tmp16840;
  wire tmp16841;
  wire tmp16842;
  wire tmp16843;
  wire tmp16844;
  wire tmp16845;
  wire tmp16846;
  wire tmp16847;
  wire tmp16848;
  wire tmp16849;
  wire tmp16850;
  wire tmp16851;
  wire tmp16852;
  wire tmp16853;
  wire tmp16854;
  wire tmp16855;
  wire tmp16856;
  wire tmp16857;
  wire tmp16858;
  wire tmp16859;
  wire tmp16860;
  wire tmp16861;
  wire tmp16862;
  wire tmp16863;
  wire tmp16864;
  wire tmp16865;
  wire tmp16866;
  wire tmp16867;
  wire tmp16868;
  wire tmp16869;
  wire tmp16870;
  wire tmp16871;
  wire tmp16872;
  wire tmp16873;
  wire tmp16874;
  wire tmp16875;
  wire tmp16876;
  wire tmp16877;
  wire tmp16878;
  wire tmp16879;
  wire tmp16880;
  wire tmp16881;
  wire tmp16882;
  wire tmp16883;
  wire tmp16884;
  wire tmp16885;
  wire tmp16886;
  wire tmp16887;
  wire tmp16888;
  wire tmp16889;
  wire tmp16890;
  wire tmp16891;
  wire tmp16892;
  wire tmp16893;
  wire tmp16894;
  wire tmp16895;
  wire tmp16896;
  wire tmp16897;
  wire tmp16898;
  wire tmp16899;
  wire tmp16900;
  wire tmp16901;
  wire tmp16902;
  wire tmp16903;
  wire tmp16904;
  wire tmp16905;
  wire tmp16906;
  wire tmp16907;
  wire tmp16908;
  wire tmp16909;
  wire tmp16910;
  wire tmp16911;
  wire tmp16912;
  wire tmp16913;
  wire tmp16914;
  wire tmp16915;
  wire tmp16916;
  wire tmp16917;
  wire tmp16918;
  wire tmp16919;
  wire tmp16920;
  wire tmp16921;
  wire tmp16922;
  wire tmp16923;
  wire tmp16924;
  wire tmp16925;
  wire tmp16926;
  wire tmp16927;
  wire tmp16928;
  wire tmp16929;
  wire tmp16930;
  wire tmp16931;
  wire tmp16932;
  wire tmp16933;
  wire tmp16934;
  wire tmp16935;
  wire tmp16936;
  wire tmp16937;
  wire tmp16938;
  wire tmp16939;
  wire tmp16940;
  wire tmp16941;
  wire tmp16942;
  wire tmp16943;
  wire tmp16944;
  wire tmp16945;
  wire tmp16946;
  wire tmp16947;
  wire tmp16948;
  wire tmp16949;
  wire tmp16950;
  wire tmp16951;
  wire tmp16952;
  wire tmp16953;
  wire tmp16954;
  wire tmp16955;
  wire tmp16956;
  wire tmp16957;
  wire tmp16958;
  wire tmp16959;
  wire tmp16960;
  wire tmp16961;
  wire tmp16962;
  wire tmp16963;
  wire tmp16964;
  wire tmp16965;
  wire tmp16966;
  wire tmp16967;
  wire tmp16968;
  wire tmp16969;
  wire tmp16970;
  wire tmp16971;
  wire tmp16972;
  wire tmp16973;
  wire tmp16974;
  wire tmp16975;
  wire tmp16976;
  wire tmp16977;
  wire tmp16978;
  wire tmp16979;
  wire tmp16980;
  wire tmp16981;
  wire tmp16982;
  wire tmp16983;
  wire tmp16984;
  wire tmp16985;
  wire tmp16986;
  wire tmp16987;
  wire tmp16988;
  wire tmp16989;
  wire tmp16990;
  wire tmp16991;
  wire tmp16992;
  wire tmp16993;
  wire tmp16994;
  wire tmp16995;
  wire tmp16996;
  wire tmp16997;
  wire tmp16998;
  wire tmp16999;
  wire tmp17000;
  wire tmp17001;
  wire tmp17002;
  wire tmp17003;
  wire tmp17004;
  wire tmp17005;
  wire tmp17006;
  wire tmp17007;
  wire tmp17008;
  wire tmp17009;
  wire tmp17010;
  wire tmp17011;
  wire tmp17012;
  wire tmp17013;
  wire tmp17014;
  wire tmp17015;
  wire tmp17016;
  wire tmp17017;
  wire tmp17018;
  wire tmp17019;
  wire tmp17020;
  wire tmp17021;
  wire tmp17022;
  wire tmp17023;
  wire tmp17024;
  wire tmp17025;
  wire tmp17026;
  wire tmp17027;
  wire tmp17028;
  wire tmp17029;
  wire tmp17030;
  wire tmp17031;
  wire tmp17032;
  wire tmp17033;
  wire tmp17034;
  wire tmp17035;
  wire tmp17036;
  wire tmp17037;
  wire tmp17038;
  wire tmp17039;
  wire tmp17040;
  wire tmp17041;
  wire tmp17042;
  wire tmp17043;
  wire tmp17044;
  wire tmp17045;
  wire tmp17046;
  wire tmp17047;
  wire tmp17048;
  wire tmp17049;
  wire tmp17050;
  wire tmp17051;
  wire tmp17052;
  wire tmp17053;
  wire tmp17054;
  wire tmp17055;
  wire tmp17056;
  wire tmp17057;
  wire tmp17058;
  wire tmp17059;
  wire tmp17060;
  wire tmp17061;
  wire tmp17062;
  wire tmp17063;
  wire tmp17064;
  wire tmp17065;
  wire tmp17066;
  wire tmp17067;
  wire tmp17068;
  wire tmp17069;
  wire tmp17070;
  wire tmp17071;
  wire tmp17072;
  wire tmp17073;
  wire tmp17074;
  wire tmp17075;
  wire tmp17076;
  wire tmp17077;
  wire tmp17078;
  wire tmp17079;
  wire tmp17080;
  wire tmp17081;
  wire tmp17082;
  wire tmp17083;
  wire tmp17084;
  wire tmp17085;
  wire tmp17086;
  wire tmp17087;
  wire tmp17088;
  wire tmp17089;
  wire tmp17090;
  wire tmp17091;
  wire tmp17092;
  wire tmp17093;
  wire tmp17094;
  wire tmp17095;
  wire tmp17096;
  wire tmp17097;
  wire tmp17098;
  wire tmp17099;
  wire tmp17100;
  wire tmp17101;
  wire tmp17102;
  wire tmp17103;
  wire tmp17104;
  wire tmp17105;
  wire tmp17106;
  wire tmp17107;
  wire tmp17108;
  wire tmp17109;
  wire tmp17110;
  wire tmp17111;
  wire tmp17112;
  wire tmp17113;
  wire tmp17114;
  wire tmp17115;
  wire tmp17116;
  wire tmp17117;
  wire tmp17118;
  wire tmp17119;
  wire tmp17120;
  wire tmp17121;
  wire tmp17122;
  wire tmp17123;
  wire tmp17124;
  wire tmp17125;
  wire tmp17126;
  wire tmp17127;
  wire tmp17128;
  wire tmp17129;
  wire tmp17130;
  wire tmp17131;
  wire tmp17132;
  wire tmp17133;
  wire tmp17134;
  wire tmp17135;
  wire tmp17136;
  wire tmp17137;
  wire tmp17138;
  wire tmp17139;
  wire tmp17140;
  wire tmp17141;
  wire tmp17142;
  wire tmp17143;
  wire tmp17144;
  wire tmp17145;
  wire tmp17146;
  wire tmp17147;
  wire tmp17148;
  wire tmp17149;
  wire tmp17150;
  wire tmp17151;
  wire tmp17152;
  wire tmp17153;
  wire tmp17154;
  wire tmp17155;
  wire tmp17156;
  wire tmp17157;
  wire tmp17158;
  wire tmp17159;
  wire tmp17160;
  wire tmp17161;
  wire tmp17162;
  wire tmp17163;
  wire tmp17164;
  wire tmp17165;
  wire tmp17166;
  wire tmp17167;
  wire tmp17168;
  wire tmp17169;
  wire tmp17170;
  wire tmp17171;
  wire tmp17172;
  wire tmp17173;
  wire tmp17174;
  wire tmp17175;
  wire tmp17176;
  wire tmp17177;
  wire tmp17178;
  wire tmp17179;
  wire tmp17180;
  wire tmp17181;
  wire tmp17182;
  wire tmp17183;
  wire tmp17184;
  wire tmp17185;
  wire tmp17186;
  wire tmp17187;
  wire tmp17188;
  wire tmp17189;
  wire tmp17190;
  wire tmp17191;
  wire tmp17192;
  wire tmp17193;
  wire tmp17194;
  wire tmp17195;
  wire tmp17196;
  wire tmp17197;
  wire tmp17198;
  wire tmp17199;
  wire tmp17200;
  wire tmp17201;
  wire tmp17202;
  wire tmp17203;
  wire tmp17204;
  wire tmp17205;
  wire tmp17206;
  wire tmp17207;
  wire tmp17208;
  wire tmp17209;
  wire tmp17210;
  wire tmp17211;
  wire tmp17212;
  wire tmp17213;
  wire tmp17214;
  wire tmp17215;
  wire tmp17216;
  wire tmp17217;
  wire tmp17218;
  wire tmp17219;
  wire tmp17220;
  wire tmp17221;
  wire tmp17222;
  wire tmp17223;
  wire tmp17224;
  wire tmp17225;
  wire tmp17226;
  wire tmp17227;
  wire tmp17228;
  wire tmp17229;
  wire tmp17230;
  wire tmp17231;
  wire tmp17232;
  wire tmp17233;
  wire tmp17234;
  wire tmp17235;
  wire tmp17236;
  wire tmp17237;
  wire tmp17238;
  wire tmp17239;
  wire tmp17240;
  wire tmp17241;
  wire tmp17242;
  wire tmp17243;
  wire tmp17244;
  wire tmp17245;
  wire tmp17246;
  wire tmp17247;
  wire tmp17248;
  wire tmp17249;
  wire tmp17250;
  wire tmp17251;
  wire tmp17252;
  wire tmp17253;
  wire tmp17254;
  wire tmp17255;
  wire tmp17256;
  wire tmp17257;
  wire tmp17258;
  wire tmp17259;
  wire tmp17260;
  wire tmp17261;
  wire tmp17262;
  wire tmp17263;
  wire tmp17264;
  wire tmp17265;
  wire tmp17266;
  wire tmp17267;
  wire tmp17268;
  wire tmp17269;
  wire tmp17270;
  wire tmp17271;
  wire tmp17272;
  wire tmp17273;
  wire tmp17274;
  wire tmp17275;
  wire tmp17276;
  wire tmp17277;
  wire tmp17278;
  wire tmp17279;
  wire tmp17280;
  wire tmp17281;
  wire tmp17282;
  wire tmp17283;
  wire tmp17284;
  wire tmp17285;
  wire tmp17286;
  wire tmp17287;
  wire tmp17288;
  wire tmp17289;
  wire tmp17290;
  wire tmp17291;
  wire tmp17292;
  wire tmp17293;
  wire tmp17294;
  wire tmp17295;
  wire tmp17296;
  wire tmp17297;
  wire tmp17298;
  wire tmp17299;
  wire tmp17300;
  wire tmp17301;
  wire tmp17302;
  wire tmp17303;
  wire tmp17304;
  wire tmp17305;
  wire tmp17306;
  wire tmp17307;
  wire tmp17308;
  wire tmp17309;
  wire tmp17310;
  wire tmp17311;
  wire tmp17312;
  wire tmp17313;
  wire tmp17314;
  wire tmp17315;
  wire tmp17316;
  wire tmp17317;
  wire tmp17318;
  wire tmp17319;
  wire tmp17320;
  wire tmp17321;
  wire tmp17322;
  wire tmp17323;
  wire tmp17324;
  wire tmp17325;
  wire tmp17326;
  wire tmp17327;
  wire tmp17328;
  wire tmp17329;
  wire tmp17330;
  wire tmp17331;
  wire tmp17332;
  wire tmp17333;
  wire tmp17334;
  wire tmp17335;
  wire tmp17336;
  wire tmp17337;
  wire tmp17338;
  wire tmp17339;
  wire tmp17340;
  wire tmp17341;
  wire tmp17342;
  wire tmp17343;
  wire tmp17344;
  wire tmp17345;
  wire tmp17346;
  wire tmp17347;
  wire tmp17348;
  wire tmp17349;
  wire tmp17350;
  wire tmp17351;
  wire tmp17352;
  wire tmp17353;
  wire tmp17354;
  wire tmp17355;
  wire tmp17356;
  wire tmp17357;
  wire tmp17358;
  wire tmp17359;
  wire tmp17360;
  wire tmp17361;
  wire tmp17362;
  wire tmp17363;
  wire tmp17364;
  wire tmp17365;
  wire tmp17366;
  wire tmp17367;
  wire tmp17368;
  wire tmp17369;
  wire tmp17370;
  wire tmp17371;
  wire tmp17372;
  wire tmp17373;
  wire tmp17374;
  wire tmp17375;
  wire tmp17376;
  wire tmp17377;
  wire tmp17378;
  wire tmp17379;
  wire tmp17380;
  wire tmp17381;
  wire tmp17382;
  wire tmp17383;
  wire tmp17384;
  wire tmp17385;
  wire tmp17386;
  wire tmp17387;
  wire tmp17388;
  wire tmp17389;
  wire tmp17390;
  wire tmp17391;
  wire tmp17392;
  wire tmp17393;
  wire tmp17394;
  wire tmp17395;
  wire tmp17396;
  wire tmp17397;
  wire tmp17398;
  wire tmp17399;
  wire tmp17400;
  wire tmp17401;
  wire tmp17402;
  wire tmp17403;
  wire tmp17404;
  wire tmp17405;
  wire tmp17406;
  wire tmp17407;
  wire tmp17408;
  wire tmp17409;
  wire tmp17410;
  wire tmp17411;
  wire tmp17412;
  wire tmp17413;
  wire tmp17414;
  wire tmp17415;
  wire tmp17416;
  wire tmp17417;
  wire tmp17418;
  wire tmp17419;
  wire tmp17420;
  wire tmp17421;
  wire tmp17422;
  wire tmp17423;
  wire tmp17424;
  wire tmp17425;
  wire tmp17426;
  wire tmp17427;
  wire tmp17428;
  wire tmp17429;
  wire tmp17430;
  wire tmp17431;
  wire tmp17432;
  wire tmp17433;
  wire tmp17434;
  wire tmp17435;
  wire tmp17436;
  wire tmp17437;
  wire tmp17438;
  wire tmp17439;
  wire tmp17440;
  wire tmp17441;
  wire tmp17442;
  wire tmp17443;
  wire tmp17444;
  wire tmp17445;
  wire tmp17446;
  wire tmp17447;
  wire tmp17448;
  wire tmp17449;
  wire tmp17450;
  wire tmp17451;
  wire tmp17452;
  wire tmp17453;
  wire tmp17454;
  wire tmp17455;
  wire tmp17456;
  wire tmp17457;
  wire tmp17458;
  wire tmp17459;
  wire tmp17460;
  wire tmp17461;
  wire tmp17462;
  wire tmp17463;
  wire tmp17464;
  wire tmp17465;
  wire tmp17466;
  wire tmp17467;
  wire tmp17468;
  wire tmp17469;
  wire tmp17470;
  wire tmp17471;
  wire tmp17472;
  wire tmp17473;
  wire tmp17474;
  wire tmp17475;
  wire tmp17476;
  wire tmp17477;
  wire tmp17478;
  wire tmp17479;
  wire tmp17480;
  wire tmp17481;
  wire tmp17482;
  wire tmp17483;
  wire tmp17484;
  wire tmp17485;
  wire tmp17486;
  wire tmp17487;
  wire tmp17488;
  wire tmp17489;
  wire tmp17490;
  wire tmp17491;
  wire tmp17492;
  wire tmp17493;
  wire tmp17494;
  wire tmp17495;
  wire tmp17496;
  wire tmp17497;
  wire tmp17498;
  wire tmp17499;
  wire tmp17500;
  wire tmp17501;
  wire tmp17502;
  wire tmp17503;
  wire tmp17504;
  wire tmp17505;
  wire tmp17506;
  wire tmp17507;
  wire tmp17508;
  wire tmp17509;
  wire tmp17510;
  wire tmp17511;
  wire tmp17512;
  wire tmp17513;
  wire tmp17514;
  wire tmp17515;
  wire tmp17516;
  wire tmp17517;
  wire tmp17518;
  wire tmp17519;
  wire tmp17520;
  wire tmp17521;
  wire tmp17522;
  wire tmp17523;
  wire tmp17524;
  wire tmp17525;
  wire tmp17526;
  wire tmp17527;
  wire tmp17528;
  wire tmp17529;
  wire tmp17530;
  wire tmp17531;
  wire tmp17532;
  wire tmp17533;
  wire tmp17534;
  wire tmp17535;
  wire tmp17536;
  wire tmp17537;
  wire tmp17538;
  wire tmp17539;
  wire tmp17540;
  wire tmp17541;
  wire tmp17542;
  wire tmp17543;
  wire tmp17544;
  wire tmp17545;
  wire tmp17546;
  wire tmp17547;
  wire tmp17548;
  wire tmp17549;
  wire tmp17550;
  wire tmp17551;
  wire tmp17552;
  wire tmp17553;
  wire tmp17554;
  wire tmp17555;
  wire tmp17556;
  wire tmp17557;
  wire tmp17558;
  wire tmp17559;
  wire tmp17560;
  wire tmp17561;
  wire tmp17562;
  wire tmp17563;
  wire tmp17564;
  wire tmp17565;
  wire tmp17566;
  wire tmp17567;
  wire tmp17568;
  wire tmp17569;
  wire tmp17570;
  wire tmp17571;
  wire tmp17572;
  wire tmp17573;
  wire tmp17574;
  wire tmp17575;
  wire tmp17576;
  wire tmp17577;
  wire tmp17578;
  wire tmp17579;
  wire tmp17580;
  wire tmp17581;
  wire tmp17582;
  wire tmp17583;
  wire tmp17584;
  wire tmp17585;
  wire tmp17586;
  wire tmp17587;
  wire tmp17588;
  wire tmp17589;
  wire tmp17590;
  wire tmp17591;
  wire tmp17592;
  wire tmp17593;
  wire tmp17594;
  wire tmp17595;
  wire tmp17596;
  wire tmp17597;
  wire tmp17598;
  wire tmp17599;
  wire tmp17600;
  wire tmp17601;
  wire tmp17602;
  wire tmp17603;
  wire tmp17604;
  wire tmp17605;
  wire tmp17606;
  wire tmp17607;
  wire tmp17608;
  wire tmp17609;
  wire tmp17610;
  wire tmp17611;
  wire tmp17612;
  wire tmp17613;
  wire tmp17614;
  wire tmp17615;
  wire tmp17616;
  wire tmp17617;
  wire tmp17618;
  wire tmp17619;
  wire tmp17620;
  wire tmp17621;
  wire tmp17622;
  wire tmp17623;
  wire tmp17624;
  wire tmp17625;
  wire tmp17626;
  wire tmp17627;
  wire tmp17628;
  wire tmp17629;
  wire tmp17630;
  wire tmp17631;
  wire tmp17632;
  wire tmp17633;
  wire tmp17634;
  wire tmp17635;
  wire tmp17636;
  wire tmp17637;
  wire tmp17638;
  wire tmp17639;
  wire tmp17640;
  wire tmp17641;
  wire tmp17642;
  wire tmp17643;
  wire tmp17644;
  wire tmp17645;
  wire tmp17646;
  wire tmp17647;
  wire tmp17648;
  wire tmp17649;
  wire tmp17650;
  wire tmp17651;
  wire tmp17652;
  wire tmp17653;
  wire tmp17654;
  wire tmp17655;
  wire tmp17656;
  wire tmp17657;
  wire tmp17658;
  wire tmp17659;
  wire tmp17660;
  wire tmp17661;
  wire tmp17662;
  wire tmp17663;
  wire tmp17664;
  wire tmp17665;
  wire tmp17666;
  wire tmp17667;
  wire tmp17668;
  wire tmp17669;
  wire tmp17670;
  wire tmp17671;
  wire tmp17672;
  wire tmp17673;
  wire tmp17674;
  wire tmp17675;
  wire tmp17676;
  wire tmp17677;
  wire tmp17678;
  wire tmp17679;
  wire tmp17680;
  wire tmp17681;
  wire tmp17682;
  wire tmp17683;
  wire tmp17684;
  wire tmp17685;
  wire tmp17686;
  wire tmp17687;
  wire tmp17688;
  wire tmp17689;
  wire tmp17690;
  wire tmp17691;
  wire tmp17692;
  wire tmp17693;
  wire tmp17694;
  wire tmp17695;
  wire tmp17696;
  wire tmp17697;
  wire tmp17698;
  wire tmp17699;
  wire tmp17700;
  wire tmp17701;
  wire tmp17702;
  wire tmp17703;
  wire tmp17704;
  wire tmp17705;
  wire tmp17706;
  wire tmp17707;
  wire tmp17708;
  wire tmp17709;
  wire tmp17710;
  wire tmp17711;
  wire tmp17712;
  wire tmp17713;
  wire tmp17714;
  wire tmp17715;
  wire tmp17716;
  wire tmp17717;
  wire tmp17718;
  wire tmp17719;
  wire tmp17720;
  wire tmp17721;
  wire tmp17722;
  wire tmp17723;
  wire tmp17724;
  wire tmp17725;
  wire tmp17726;
  wire tmp17727;
  wire tmp17728;
  wire tmp17729;
  wire tmp17730;
  wire tmp17731;
  wire tmp17732;
  wire tmp17733;
  wire tmp17734;
  wire tmp17735;
  wire tmp17736;
  wire tmp17737;
  wire tmp17738;
  wire tmp17739;
  wire tmp17740;
  wire tmp17741;
  wire tmp17742;
  wire tmp17743;
  wire tmp17744;
  wire tmp17745;
  wire tmp17746;
  wire tmp17747;
  wire tmp17748;
  wire tmp17749;
  wire tmp17750;
  wire tmp17751;
  wire tmp17752;
  wire tmp17753;
  wire tmp17754;
  wire tmp17755;
  wire tmp17756;
  wire tmp17757;
  wire tmp17758;
  wire tmp17759;
  wire tmp17760;
  wire tmp17761;
  wire tmp17762;
  wire tmp17763;
  wire tmp17764;
  wire tmp17765;
  wire tmp17766;
  wire tmp17767;
  wire tmp17768;
  wire tmp17769;
  wire tmp17770;
  wire tmp17771;
  wire tmp17772;
  wire tmp17773;
  wire tmp17774;
  wire tmp17775;
  wire tmp17776;
  wire tmp17777;
  wire tmp17778;
  wire tmp17779;
  wire tmp17780;
  wire tmp17781;
  wire tmp17782;
  wire tmp17783;
  wire tmp17784;
  wire tmp17785;
  wire tmp17786;
  wire tmp17787;
  wire tmp17788;
  wire tmp17789;
  wire tmp17790;
  wire tmp17791;
  wire tmp17792;
  wire tmp17793;
  wire tmp17794;
  wire tmp17795;
  wire tmp17796;
  wire tmp17797;
  wire tmp17798;
  wire tmp17799;
  wire tmp17800;
  wire tmp17801;
  wire tmp17802;
  wire tmp17803;
  wire tmp17804;
  wire tmp17805;
  wire tmp17806;
  wire tmp17807;
  wire tmp17808;
  wire tmp17809;
  wire tmp17810;
  wire tmp17811;
  wire tmp17812;
  wire tmp17813;
  wire tmp17814;
  wire tmp17815;
  wire tmp17816;
  wire tmp17817;
  wire tmp17818;
  wire tmp17819;
  wire tmp17820;
  wire tmp17821;
  wire tmp17822;
  wire tmp17823;
  wire tmp17824;
  wire tmp17825;
  wire tmp17826;
  wire tmp17827;
  wire tmp17828;
  wire tmp17829;
  wire tmp17830;
  wire tmp17831;
  wire tmp17832;
  wire tmp17833;
  wire tmp17834;
  wire tmp17835;
  wire tmp17836;
  wire tmp17837;
  wire tmp17838;
  wire tmp17839;
  wire tmp17840;
  wire tmp17841;
  wire tmp17842;
  wire tmp17843;
  wire tmp17844;
  wire tmp17845;
  wire tmp17846;
  wire tmp17847;
  wire tmp17848;
  wire tmp17849;
  wire tmp17850;
  wire tmp17851;
  wire tmp17852;
  wire tmp17853;
  wire tmp17854;
  wire tmp17855;
  wire tmp17856;
  wire tmp17857;
  wire tmp17858;
  wire tmp17859;
  wire tmp17860;
  wire tmp17861;
  wire tmp17862;
  wire tmp17863;
  wire tmp17864;
  wire tmp17865;
  wire tmp17866;
  wire tmp17867;
  wire tmp17868;
  wire tmp17869;
  wire tmp17870;
  wire tmp17871;
  wire tmp17872;
  wire tmp17873;
  wire tmp17874;
  wire tmp17875;
  wire tmp17876;
  wire tmp17877;
  wire tmp17878;
  wire tmp17879;
  wire tmp17880;
  wire tmp17881;
  wire tmp17882;
  wire tmp17883;
  wire tmp17884;
  wire tmp17885;
  wire tmp17886;
  wire tmp17887;
  wire tmp17888;
  wire tmp17889;
  wire tmp17890;
  wire tmp17891;
  wire tmp17892;
  wire tmp17893;
  wire tmp17894;
  wire tmp17895;
  wire tmp17896;
  wire tmp17897;
  wire tmp17898;
  wire tmp17899;
  wire tmp17900;
  wire tmp17901;
  wire tmp17902;
  wire tmp17903;
  wire tmp17904;
  wire tmp17905;
  wire tmp17906;
  wire tmp17907;
  wire tmp17908;
  wire tmp17909;
  wire tmp17910;
  wire tmp17911;
  wire tmp17912;
  wire tmp17913;
  wire tmp17914;
  wire tmp17915;
  wire tmp17916;
  wire tmp17917;
  wire tmp17918;
  wire tmp17919;
  wire tmp17920;
  wire tmp17921;
  wire tmp17922;
  wire tmp17923;
  wire tmp17924;
  wire tmp17925;
  wire tmp17926;
  wire tmp17927;
  wire tmp17928;
  wire tmp17929;
  wire tmp17930;
  wire tmp17931;
  wire tmp17932;
  wire tmp17933;
  wire tmp17934;
  wire tmp17935;
  wire tmp17936;
  wire tmp17937;
  wire tmp17938;
  wire tmp17939;
  wire tmp17940;
  wire tmp17941;
  wire tmp17942;
  wire tmp17943;
  wire tmp17944;
  wire tmp17945;
  wire tmp17946;
  wire tmp17947;
  wire tmp17948;
  wire tmp17949;
  wire tmp17950;
  wire tmp17951;
  wire tmp17952;
  wire tmp17953;
  wire tmp17954;
  wire tmp17955;
  wire tmp17956;
  wire tmp17957;
  wire tmp17958;
  wire tmp17959;
  wire tmp17960;
  wire tmp17961;
  wire tmp17962;
  wire tmp17963;
  wire tmp17964;
  wire tmp17965;
  wire tmp17966;
  wire tmp17967;
  wire tmp17968;
  wire tmp17969;
  wire tmp17970;
  wire tmp17971;
  wire tmp17972;
  wire tmp17973;
  wire tmp17974;
  wire tmp17975;
  wire tmp17976;
  wire tmp17977;
  wire tmp17978;
  wire tmp17979;
  wire tmp17980;
  wire tmp17981;
  wire tmp17982;
  wire tmp17983;
  wire tmp17984;
  wire tmp17985;
  wire tmp17986;
  wire tmp17987;
  wire tmp17988;
  wire tmp17989;
  wire tmp17990;
  wire tmp17991;
  wire tmp17992;
  wire tmp17993;
  wire tmp17994;
  wire tmp17995;
  wire tmp17996;
  wire tmp17997;
  wire tmp17998;
  wire tmp17999;
  wire tmp18000;
  wire tmp18001;
  wire tmp18002;
  wire tmp18003;
  wire tmp18004;
  wire tmp18005;
  wire tmp18006;
  wire tmp18007;
  wire tmp18008;
  wire tmp18009;
  wire tmp18010;
  wire tmp18011;
  wire tmp18012;
  wire tmp18013;
  wire tmp18014;
  wire tmp18015;
  wire tmp18016;
  wire tmp18017;
  wire tmp18018;
  wire tmp18019;
  wire tmp18020;
  wire tmp18021;
  wire tmp18022;
  wire tmp18023;
  wire tmp18024;
  wire tmp18025;
  wire tmp18026;
  wire tmp18027;
  wire tmp18028;
  wire tmp18029;
  wire tmp18030;
  wire tmp18031;
  wire tmp18032;
  wire tmp18033;
  wire tmp18034;
  wire tmp18035;
  wire tmp18036;
  wire tmp18037;
  wire tmp18038;
  wire tmp18039;
  wire tmp18040;
  wire tmp18041;
  wire tmp18042;
  wire tmp18043;
  wire tmp18044;
  wire tmp18045;
  wire tmp18046;
  wire tmp18047;
  wire tmp18048;
  wire tmp18049;
  wire tmp18050;
  wire tmp18051;
  wire tmp18052;
  wire tmp18053;
  wire tmp18054;
  wire tmp18055;
  wire tmp18056;
  wire tmp18057;
  wire tmp18058;
  wire tmp18059;
  wire tmp18060;
  wire tmp18061;
  wire tmp18062;
  wire tmp18063;
  wire tmp18064;
  wire tmp18065;
  wire tmp18066;
  wire tmp18067;
  wire tmp18068;
  wire tmp18069;
  wire tmp18070;
  wire tmp18071;
  wire tmp18072;
  wire tmp18073;
  wire tmp18074;
  wire tmp18075;
  wire tmp18076;
  wire tmp18077;
  wire tmp18078;
  wire tmp18079;
  wire tmp18080;
  wire tmp18081;
  wire tmp18082;
  wire tmp18083;
  wire tmp18084;
  wire tmp18085;
  wire tmp18086;
  wire tmp18087;
  wire tmp18088;
  wire tmp18089;
  wire tmp18090;
  wire tmp18091;
  wire tmp18092;
  wire tmp18093;
  wire tmp18094;
  wire tmp18095;
  wire tmp18096;
  wire tmp18097;
  wire tmp18098;
  wire tmp18099;
  wire tmp18100;
  wire tmp18101;
  wire tmp18102;
  wire tmp18103;
  wire tmp18104;
  wire tmp18105;
  wire tmp18106;
  wire tmp18107;
  wire tmp18108;
  wire tmp18109;
  wire tmp18110;
  wire tmp18111;
  wire tmp18112;
  wire tmp18113;
  wire tmp18114;
  wire tmp18115;
  wire tmp18116;
  wire tmp18117;
  wire tmp18118;
  wire tmp18119;
  wire tmp18120;
  wire tmp18121;
  wire tmp18122;
  wire tmp18123;
  wire tmp18124;
  wire tmp18125;
  wire tmp18126;
  wire tmp18127;
  wire tmp18128;
  wire tmp18129;
  wire tmp18130;
  wire tmp18131;
  wire tmp18132;
  wire tmp18133;
  wire tmp18134;
  wire tmp18135;
  wire tmp18136;
  wire tmp18137;
  wire tmp18138;
  wire tmp18139;
  wire tmp18140;
  wire tmp18141;
  wire tmp18142;
  wire tmp18143;
  wire tmp18144;
  wire tmp18145;
  wire tmp18146;
  wire tmp18147;
  wire tmp18148;
  wire tmp18149;
  wire tmp18150;
  wire tmp18151;
  wire tmp18152;
  wire tmp18153;
  wire tmp18154;
  wire tmp18155;
  wire tmp18156;
  wire tmp18157;
  wire tmp18158;
  wire tmp18159;
  wire tmp18160;
  wire tmp18161;
  wire tmp18162;
  wire tmp18163;
  wire tmp18164;
  wire tmp18165;
  wire tmp18166;
  wire tmp18167;
  wire tmp18168;
  wire tmp18169;
  wire tmp18170;
  wire tmp18171;
  wire tmp18172;
  wire tmp18173;
  wire tmp18174;
  wire tmp18175;
  wire tmp18176;
  wire tmp18177;
  wire tmp18178;
  wire tmp18179;
  wire tmp18180;
  wire tmp18181;
  wire tmp18182;
  wire tmp18183;
  wire tmp18184;
  wire tmp18185;
  wire tmp18186;
  wire tmp18187;
  wire tmp18188;
  wire tmp18189;
  wire tmp18190;
  wire tmp18191;
  wire tmp18192;
  wire tmp18193;
  wire tmp18194;
  wire tmp18195;
  wire tmp18196;
  wire tmp18197;
  wire tmp18198;
  wire tmp18199;
  wire tmp18200;
  wire tmp18201;
  wire tmp18202;
  wire tmp18203;
  wire tmp18204;
  wire tmp18205;
  wire tmp18206;
  wire tmp18207;
  wire tmp18208;
  wire tmp18209;
  wire tmp18210;
  wire tmp18211;
  wire tmp18212;
  wire tmp18213;
  wire tmp18214;
  wire tmp18215;
  wire tmp18216;
  wire tmp18217;
  wire tmp18218;
  wire tmp18219;
  wire tmp18220;
  wire tmp18221;
  wire tmp18222;
  wire tmp18223;
  wire tmp18224;
  wire tmp18225;
  wire tmp18226;
  wire tmp18227;
  wire tmp18228;
  wire tmp18229;
  wire tmp18230;
  wire tmp18231;
  wire tmp18232;
  wire tmp18233;
  wire tmp18234;
  wire tmp18235;
  wire tmp18236;
  wire tmp18237;
  wire tmp18238;
  wire tmp18239;
  wire tmp18240;
  wire tmp18241;
  wire tmp18242;
  wire tmp18243;
  wire tmp18244;
  wire tmp18245;
  wire tmp18246;
  wire tmp18247;
  wire tmp18248;
  wire tmp18249;
  wire tmp18250;
  wire tmp18251;
  wire tmp18252;
  wire tmp18253;
  wire tmp18254;
  wire tmp18255;
  wire tmp18256;
  wire tmp18257;
  wire tmp18258;
  wire tmp18259;
  wire tmp18260;
  wire tmp18261;
  wire tmp18262;
  wire tmp18263;
  wire tmp18264;
  wire tmp18265;
  wire tmp18266;
  wire tmp18267;
  wire tmp18268;
  wire tmp18269;
  wire tmp18270;
  wire tmp18271;
  wire tmp18272;
  wire tmp18273;
  wire tmp18274;
  wire tmp18275;
  wire tmp18276;
  wire tmp18277;
  wire tmp18278;
  wire tmp18279;
  wire tmp18280;
  wire tmp18281;
  wire tmp18282;
  wire tmp18283;
  wire tmp18284;
  wire tmp18285;
  wire tmp18286;
  wire tmp18287;
  wire tmp18288;
  wire tmp18289;
  wire tmp18290;
  wire tmp18291;
  wire tmp18292;
  wire tmp18293;
  wire tmp18294;
  wire tmp18295;
  wire tmp18296;
  wire tmp18297;
  wire tmp18298;
  wire tmp18299;
  wire tmp18300;
  wire tmp18301;
  wire tmp18302;
  wire tmp18303;
  wire tmp18304;
  wire tmp18305;
  wire tmp18306;
  wire tmp18307;
  wire tmp18308;
  wire tmp18309;
  wire tmp18310;
  wire tmp18311;
  wire tmp18312;
  wire tmp18313;
  wire tmp18314;
  wire tmp18315;
  wire tmp18316;
  wire tmp18317;
  wire tmp18318;
  wire tmp18319;
  wire tmp18320;
  wire tmp18321;
  wire tmp18322;
  wire tmp18323;
  wire tmp18324;
  wire tmp18325;
  wire tmp18326;
  wire tmp18327;
  wire tmp18328;
  wire tmp18329;
  wire tmp18330;
  wire tmp18331;
  wire tmp18332;
  wire tmp18333;
  wire tmp18334;
  wire tmp18335;
  wire tmp18336;
  wire tmp18337;
  wire tmp18338;
  wire tmp18339;
  wire tmp18340;
  wire tmp18341;
  wire tmp18342;
  wire tmp18343;
  wire tmp18344;
  wire tmp18345;
  wire tmp18346;
  wire tmp18347;
  wire tmp18348;
  wire tmp18349;
  wire tmp18350;
  wire tmp18351;
  wire tmp18352;
  wire tmp18353;
  wire tmp18354;
  wire tmp18355;
  wire tmp18356;
  wire tmp18357;
  wire tmp18358;
  wire tmp18359;
  wire tmp18360;
  wire tmp18361;
  wire tmp18362;
  wire tmp18363;
  wire tmp18364;
  wire tmp18365;
  wire tmp18366;
  wire tmp18367;
  wire tmp18368;
  wire tmp18369;
  wire tmp18370;
  wire tmp18371;
  wire tmp18372;
  wire tmp18373;
  wire tmp18374;
  wire tmp18375;
  wire tmp18376;
  wire tmp18377;
  wire tmp18378;
  wire tmp18379;
  wire tmp18380;
  wire tmp18381;
  wire tmp18382;
  wire tmp18383;
  wire tmp18384;
  wire tmp18385;
  wire tmp18386;
  wire tmp18387;
  wire tmp18388;
  wire tmp18389;
  wire tmp18390;
  wire tmp18391;
  wire tmp18392;
  wire tmp18393;
  wire tmp18394;
  wire tmp18395;
  wire tmp18396;
  wire tmp18397;
  wire tmp18398;
  wire tmp18399;
  wire tmp18400;
  wire tmp18401;
  wire tmp18402;
  wire tmp18403;
  wire tmp18404;
  wire tmp18405;
  wire tmp18406;
  wire tmp18407;
  wire tmp18408;
  wire tmp18409;
  wire tmp18410;
  wire tmp18411;
  wire tmp18412;
  wire tmp18413;
  wire tmp18414;
  wire tmp18415;
  wire tmp18416;
  wire tmp18417;
  wire tmp18418;
  wire tmp18419;
  wire tmp18420;
  wire tmp18421;
  wire tmp18422;
  wire tmp18423;
  wire tmp18424;
  wire tmp18425;
  wire tmp18426;
  wire tmp18427;
  wire tmp18428;
  wire tmp18429;
  wire tmp18430;
  wire tmp18431;
  wire tmp18432;
  wire tmp18433;
  wire tmp18434;
  wire tmp18435;
  wire tmp18436;
  wire tmp18437;
  wire tmp18438;
  wire tmp18439;
  wire tmp18440;
  wire tmp18441;
  wire tmp18442;
  wire tmp18443;
  wire tmp18444;
  wire tmp18445;
  wire tmp18446;
  wire tmp18447;
  wire tmp18448;
  wire tmp18449;
  wire tmp18450;
  wire tmp18451;
  wire tmp18452;
  wire tmp18453;
  wire tmp18454;
  wire tmp18455;
  wire tmp18456;
  wire tmp18457;
  wire tmp18458;
  wire tmp18459;
  wire tmp18460;
  wire tmp18461;
  wire tmp18462;
  wire tmp18463;
  wire tmp18464;
  wire tmp18465;
  wire tmp18466;
  wire tmp18467;
  wire tmp18468;
  wire tmp18469;
  wire tmp18470;
  wire tmp18471;
  wire tmp18472;
  wire tmp18473;
  wire tmp18474;
  wire tmp18475;
  wire tmp18476;
  wire tmp18477;
  wire tmp18478;
  wire tmp18479;
  wire tmp18480;
  wire tmp18481;
  wire tmp18482;
  wire tmp18483;
  wire tmp18484;
  wire tmp18485;
  wire tmp18486;
  wire tmp18487;
  wire tmp18488;
  wire tmp18489;
  wire tmp18490;
  wire tmp18491;
  wire tmp18492;
  wire tmp18493;
  wire tmp18494;
  wire tmp18495;
  wire tmp18496;
  wire tmp18497;
  wire tmp18498;
  wire tmp18499;
  wire tmp18500;
  wire tmp18501;
  wire tmp18502;
  wire tmp18503;
  wire tmp18504;
  wire tmp18505;
  wire tmp18506;
  wire tmp18507;
  wire tmp18508;
  wire tmp18509;
  wire tmp18510;
  wire tmp18511;
  wire tmp18512;
  wire tmp18513;
  wire tmp18514;
  wire tmp18515;
  wire tmp18516;
  wire tmp18517;
  wire tmp18518;
  wire tmp18519;
  wire tmp18520;
  wire tmp18521;
  wire tmp18522;
  wire tmp18523;
  wire tmp18524;
  wire tmp18525;
  wire tmp18526;
  wire tmp18527;
  wire tmp18528;
  wire tmp18529;
  wire tmp18530;
  wire tmp18531;
  wire tmp18532;
  wire tmp18533;
  wire tmp18534;
  wire tmp18535;
  wire tmp18536;
  wire tmp18537;
  wire tmp18538;
  wire tmp18539;
  wire tmp18540;
  wire tmp18541;
  wire tmp18542;
  wire tmp18543;
  wire tmp18544;
  wire tmp18545;
  wire tmp18546;
  wire tmp18547;
  wire tmp18548;
  wire tmp18549;
  wire tmp18550;
  wire tmp18551;
  wire tmp18552;
  wire tmp18553;
  wire tmp18554;
  wire tmp18555;
  wire tmp18556;
  wire tmp18557;
  wire tmp18558;
  wire tmp18559;
  wire tmp18560;
  wire tmp18561;
  wire tmp18562;
  wire tmp18563;
  wire tmp18564;
  wire tmp18565;
  wire tmp18566;
  wire tmp18567;
  wire tmp18568;
  wire tmp18569;
  wire tmp18570;
  wire tmp18571;
  wire tmp18572;
  wire tmp18573;
  wire tmp18574;
  wire tmp18575;
  wire tmp18576;
  wire tmp18577;
  wire tmp18578;
  wire tmp18579;
  wire tmp18580;
  wire tmp18581;
  wire tmp18582;
  wire tmp18583;
  wire tmp18584;
  wire tmp18585;
  wire tmp18586;
  wire tmp18587;
  wire tmp18588;
  wire tmp18589;
  wire tmp18590;
  wire tmp18591;
  wire tmp18592;
  wire tmp18593;
  wire tmp18594;
  wire tmp18595;
  wire tmp18596;
  wire tmp18597;
  wire tmp18598;
  wire tmp18599;
  wire tmp18600;
  wire tmp18601;
  wire tmp18602;
  wire tmp18603;
  wire tmp18604;
  wire tmp18605;
  wire tmp18606;
  wire tmp18607;
  wire tmp18608;
  wire tmp18609;
  wire tmp18610;
  wire tmp18611;
  wire tmp18612;
  wire tmp18613;
  wire tmp18614;
  wire tmp18615;
  wire tmp18616;
  wire tmp18617;
  wire tmp18618;
  wire tmp18619;
  wire tmp18620;
  wire tmp18621;
  wire tmp18622;
  wire tmp18623;
  wire tmp18624;
  wire tmp18625;
  wire tmp18626;
  wire tmp18627;
  wire tmp18628;
  wire tmp18629;
  wire tmp18630;
  wire tmp18631;
  wire tmp18632;
  wire tmp18633;
  wire tmp18634;
  wire tmp18635;
  wire tmp18636;
  wire tmp18637;
  wire tmp18638;
  wire tmp18639;
  wire tmp18640;
  wire tmp18641;
  wire tmp18642;
  wire tmp18643;
  wire tmp18644;
  wire tmp18645;
  wire tmp18646;
  wire tmp18647;
  wire tmp18648;
  wire tmp18649;
  wire tmp18650;
  wire tmp18651;
  wire tmp18652;
  wire tmp18653;
  wire tmp18654;
  wire tmp18655;
  wire tmp18656;
  wire tmp18657;
  wire tmp18658;
  wire tmp18659;
  wire tmp18660;
  wire tmp18661;
  wire tmp18662;
  wire tmp18663;
  wire tmp18664;
  wire tmp18665;
  wire tmp18666;
  wire tmp18667;
  wire tmp18668;
  wire tmp18669;
  wire tmp18670;
  wire tmp18671;
  wire tmp18672;
  wire tmp18673;
  wire tmp18674;
  wire tmp18675;
  wire tmp18676;
  wire tmp18677;
  wire tmp18678;
  wire tmp18679;
  wire tmp18680;
  wire tmp18681;
  wire tmp18682;
  wire tmp18683;
  wire tmp18684;
  wire tmp18685;
  wire tmp18686;
  wire tmp18687;
  wire tmp18688;
  wire tmp18689;
  wire tmp18690;
  wire tmp18691;
  wire tmp18692;
  wire tmp18693;
  wire tmp18694;
  wire tmp18695;
  wire tmp18696;
  wire tmp18697;
  wire tmp18698;
  wire tmp18699;
  wire tmp18700;
  wire tmp18701;
  wire tmp18702;
  wire tmp18703;
  wire tmp18704;
  wire tmp18705;
  wire tmp18706;
  wire tmp18707;
  wire tmp18708;
  wire tmp18709;
  wire tmp18710;
  wire tmp18711;
  wire tmp18712;
  wire tmp18713;
  wire tmp18714;
  wire tmp18715;
  wire tmp18716;
  wire tmp18717;
  wire tmp18718;
  wire tmp18719;
  wire tmp18720;
  wire tmp18721;
  wire tmp18722;
  wire tmp18723;
  wire tmp18724;
  wire tmp18725;
  wire tmp18726;
  wire tmp18727;
  wire tmp18728;
  wire tmp18729;
  wire tmp18730;
  wire tmp18731;
  wire tmp18732;
  wire tmp18733;
  wire tmp18734;
  wire tmp18735;
  wire tmp18736;
  wire tmp18737;
  wire tmp18738;
  wire tmp18739;
  wire tmp18740;
  wire tmp18741;
  wire tmp18742;
  wire tmp18743;
  wire tmp18744;
  wire tmp18745;
  wire tmp18746;
  wire tmp18747;
  wire tmp18748;
  wire tmp18749;
  wire tmp18750;
  wire tmp18751;
  wire tmp18752;
  wire tmp18753;
  wire tmp18754;
  wire tmp18755;
  wire tmp18756;
  wire tmp18757;
  wire tmp18758;
  wire tmp18759;
  wire tmp18760;
  wire tmp18761;
  wire tmp18762;
  wire tmp18763;
  wire tmp18764;
  wire tmp18765;
  wire tmp18766;
  wire tmp18767;
  wire tmp18768;
  wire tmp18769;
  wire tmp18770;
  wire tmp18771;
  wire tmp18772;
  wire tmp18773;
  wire tmp18774;
  wire tmp18775;
  wire tmp18776;
  wire tmp18777;
  wire tmp18778;
  wire tmp18779;
  wire tmp18780;
  wire tmp18781;
  wire tmp18782;
  wire tmp18783;
  wire tmp18784;
  wire tmp18785;
  wire tmp18786;
  wire tmp18787;
  wire tmp18788;
  wire tmp18789;
  wire tmp18790;
  wire tmp18791;
  wire tmp18792;
  wire tmp18793;
  wire tmp18794;
  wire tmp18795;
  wire tmp18796;
  wire tmp18797;
  wire tmp18798;
  wire tmp18799;
  wire tmp18800;
  wire tmp18801;
  wire tmp18802;
  wire tmp18803;
  wire tmp18804;
  wire tmp18805;
  wire tmp18806;
  wire tmp18807;
  wire tmp18808;
  wire tmp18809;
  wire tmp18810;
  wire tmp18811;
  wire tmp18812;
  wire tmp18813;
  wire tmp18814;
  wire tmp18815;
  wire tmp18816;
  wire tmp18817;
  wire tmp18818;
  wire tmp18819;
  wire tmp18820;
  wire tmp18821;
  wire tmp18822;
  wire tmp18823;
  wire tmp18824;
  wire tmp18825;
  wire tmp18826;
  wire tmp18827;
  wire tmp18828;
  wire tmp18829;
  wire tmp18830;
  wire tmp18831;
  wire tmp18832;
  wire tmp18833;
  wire tmp18834;
  wire tmp18835;
  wire tmp18836;
  wire tmp18837;
  wire tmp18838;
  wire tmp18839;
  wire tmp18840;
  wire tmp18841;
  wire tmp18842;
  wire tmp18843;
  wire tmp18844;
  wire tmp18845;
  wire tmp18846;
  wire tmp18847;
  wire tmp18848;
  wire tmp18849;
  wire tmp18850;
  wire tmp18851;
  wire tmp18852;
  wire tmp18853;
  wire tmp18854;
  wire tmp18855;
  wire tmp18856;
  wire tmp18857;
  wire tmp18858;
  wire tmp18859;
  wire tmp18860;
  wire tmp18861;
  wire tmp18862;
  wire tmp18863;
  wire tmp18864;
  wire tmp18865;
  wire tmp18866;
  wire tmp18867;
  wire tmp18868;
  wire tmp18869;
  wire tmp18870;
  wire tmp18871;
  wire tmp18872;
  wire tmp18873;
  wire tmp18874;
  wire tmp18875;
  wire tmp18876;
  wire tmp18877;
  wire tmp18878;
  wire tmp18879;
  wire tmp18880;
  wire tmp18881;
  wire tmp18882;
  wire tmp18883;
  wire tmp18884;
  wire tmp18885;
  wire tmp18886;
  wire tmp18887;
  wire tmp18888;
  wire tmp18889;
  wire tmp18890;
  wire tmp18891;
  wire tmp18892;
  wire tmp18893;
  wire tmp18894;
  wire tmp18895;
  wire tmp18896;
  wire tmp18897;
  wire tmp18898;
  wire tmp18899;
  wire tmp18900;
  wire tmp18901;
  wire tmp18902;
  wire tmp18903;
  wire tmp18904;
  wire tmp18905;
  wire tmp18906;
  wire tmp18907;
  wire tmp18908;
  wire tmp18909;
  wire tmp18910;
  wire tmp18911;
  wire tmp18912;
  wire tmp18913;
  wire tmp18914;
  wire tmp18915;
  wire tmp18916;
  wire tmp18917;
  wire tmp18918;
  wire tmp18919;
  wire tmp18920;
  wire tmp18921;
  wire tmp18922;
  wire tmp18923;
  wire tmp18924;
  wire tmp18925;
  wire tmp18926;
  wire tmp18927;
  wire tmp18928;
  wire tmp18929;
  wire tmp18930;
  wire tmp18931;
  wire tmp18932;
  wire tmp18933;
  wire tmp18934;
  wire tmp18935;
  wire tmp18936;
  wire tmp18937;
  wire tmp18938;
  wire tmp18939;
  wire tmp18940;
  wire tmp18941;
  wire tmp18942;
  wire tmp18943;
  wire tmp18944;
  wire tmp18945;
  wire tmp18946;
  wire tmp18947;
  wire tmp18948;
  wire tmp18949;
  wire tmp18950;
  wire tmp18951;
  wire tmp18952;
  wire tmp18953;
  wire tmp18954;
  wire tmp18955;
  wire tmp18956;
  wire tmp18957;
  wire tmp18958;
  wire tmp18959;
  wire tmp18960;
  wire tmp18961;
  wire tmp18962;
  wire tmp18963;
  wire tmp18964;
  wire tmp18965;
  wire tmp18966;
  wire tmp18967;
  wire tmp18968;
  wire tmp18969;
  wire tmp18970;
  wire tmp18971;
  wire tmp18972;
  wire tmp18973;
  wire tmp18974;
  wire tmp18975;
  wire tmp18976;
  wire tmp18977;
  wire tmp18978;
  wire tmp18979;
  wire tmp18980;
  wire tmp18981;
  wire tmp18982;
  wire tmp18983;
  wire tmp18984;
  wire tmp18985;
  wire tmp18986;
  wire tmp18987;
  wire tmp18988;
  wire tmp18989;
  wire tmp18990;
  wire tmp18991;
  wire tmp18992;
  wire tmp18993;
  wire tmp18994;
  wire tmp18995;
  wire tmp18996;
  wire tmp18997;
  wire tmp18998;
  wire tmp18999;
  wire tmp19000;
  wire tmp19001;
  wire tmp19002;
  wire tmp19003;
  wire tmp19004;
  wire tmp19005;
  wire tmp19006;
  wire tmp19007;
  wire tmp19008;
  wire tmp19009;
  wire tmp19010;
  wire tmp19011;
  wire tmp19012;
  wire tmp19013;
  wire tmp19014;
  wire tmp19015;
  wire tmp19016;
  wire tmp19017;
  wire tmp19018;
  wire tmp19019;
  wire tmp19020;
  wire tmp19021;
  wire tmp19022;
  wire tmp19023;
  wire tmp19024;
  wire tmp19025;
  wire tmp19026;
  wire tmp19027;
  wire tmp19028;
  wire tmp19029;
  wire tmp19030;
  wire tmp19031;
  wire tmp19032;
  wire tmp19033;
  wire tmp19034;
  wire tmp19035;
  wire tmp19036;
  wire tmp19037;
  wire tmp19038;
  wire tmp19039;
  wire tmp19040;
  wire tmp19041;
  wire tmp19042;
  wire tmp19043;
  wire tmp19044;
  wire tmp19045;
  wire tmp19046;
  wire tmp19047;
  wire tmp19048;
  wire tmp19049;
  wire tmp19050;
  wire tmp19051;
  wire tmp19052;
  wire tmp19053;
  wire tmp19054;
  wire tmp19055;
  wire tmp19056;
  wire tmp19057;
  wire tmp19058;
  wire tmp19059;
  wire tmp19060;
  wire tmp19061;
  wire tmp19062;
  wire tmp19063;
  wire tmp19064;
  wire tmp19065;
  wire tmp19066;
  wire tmp19067;
  wire tmp19068;
  wire tmp19069;
  wire tmp19070;
  wire tmp19071;
  wire tmp19072;
  wire tmp19073;
  wire tmp19074;
  wire tmp19075;
  wire tmp19076;
  wire tmp19077;
  wire tmp19078;
  wire tmp19079;
  wire tmp19080;
  wire tmp19081;
  wire tmp19082;
  wire tmp19083;
  wire tmp19084;
  wire tmp19085;
  wire tmp19086;
  wire tmp19087;
  wire tmp19088;
  wire tmp19089;
  wire tmp19090;
  wire tmp19091;
  wire tmp19092;
  wire tmp19093;
  wire tmp19094;
  wire tmp19095;
  wire tmp19096;
  wire tmp19097;
  wire tmp19098;
  wire tmp19099;
  wire tmp19100;
  wire tmp19101;
  wire tmp19102;
  wire tmp19103;
  wire tmp19104;
  wire tmp19105;
  wire tmp19106;
  wire tmp19107;
  wire tmp19108;
  wire tmp19109;
  wire tmp19110;
  wire tmp19111;
  wire tmp19112;
  wire tmp19113;
  wire tmp19114;
  wire tmp19115;
  wire tmp19116;
  wire tmp19117;
  wire tmp19118;
  wire tmp19119;
  wire tmp19120;
  wire tmp19121;
  wire tmp19122;
  wire tmp19123;
  wire tmp19124;
  wire tmp19125;
  wire tmp19126;
  wire tmp19127;
  wire tmp19128;
  wire tmp19129;
  wire tmp19130;
  wire tmp19131;
  wire tmp19132;
  wire tmp19133;
  wire tmp19134;
  wire tmp19135;
  wire tmp19136;
  wire tmp19137;
  wire tmp19138;
  wire tmp19139;
  wire tmp19140;
  wire tmp19141;
  wire tmp19142;
  wire tmp19143;
  wire tmp19144;
  wire tmp19145;
  wire tmp19146;
  wire tmp19147;
  wire tmp19148;
  wire tmp19149;
  wire tmp19150;
  wire tmp19151;
  wire tmp19152;
  wire tmp19153;
  wire tmp19154;
  wire tmp19155;
  wire tmp19156;
  wire tmp19157;
  wire tmp19158;
  wire tmp19159;
  wire tmp19160;
  wire tmp19161;
  wire tmp19162;
  wire tmp19163;
  wire tmp19164;
  wire tmp19165;
  wire tmp19166;
  wire tmp19167;
  wire tmp19168;
  wire tmp19169;
  wire tmp19170;
  wire tmp19171;
  wire tmp19172;
  wire tmp19173;
  wire tmp19174;
  wire tmp19175;
  wire tmp19176;
  wire tmp19177;
  wire tmp19178;
  wire tmp19179;
  wire tmp19180;
  wire tmp19181;
  wire tmp19182;
  wire tmp19183;
  wire tmp19184;
  wire tmp19185;
  wire tmp19186;
  wire tmp19187;
  wire tmp19188;
  wire tmp19189;
  wire tmp19190;
  wire tmp19191;
  wire tmp19192;
  wire tmp19193;
  wire tmp19194;
  wire tmp19195;
  wire tmp19196;
  wire tmp19197;
  wire tmp19198;
  wire tmp19199;
  wire tmp19200;
  wire tmp19201;
  wire tmp19202;
  wire tmp19203;
  wire tmp19204;
  wire tmp19205;
  wire tmp19206;
  wire tmp19207;
  wire tmp19208;
  wire tmp19209;
  wire tmp19210;
  wire tmp19211;
  wire tmp19212;
  wire tmp19213;
  wire tmp19214;
  wire tmp19215;
  wire tmp19216;
  wire tmp19217;
  wire tmp19218;
  wire tmp19219;
  wire tmp19220;
  wire tmp19221;
  wire tmp19222;
  wire tmp19223;
  wire tmp19224;
  wire tmp19225;
  wire tmp19226;
  wire tmp19227;
  wire tmp19228;
  wire tmp19229;
  wire tmp19230;
  wire tmp19231;
  wire tmp19232;
  wire tmp19233;
  wire tmp19234;
  wire tmp19235;
  wire tmp19236;
  wire tmp19237;
  wire tmp19238;
  wire tmp19239;
  wire tmp19240;
  wire tmp19241;
  wire tmp19242;
  wire tmp19243;
  wire tmp19244;
  wire tmp19245;
  wire tmp19246;
  wire tmp19247;
  wire tmp19248;
  wire tmp19249;
  wire tmp19250;
  wire tmp19251;
  wire tmp19252;
  wire tmp19253;
  wire tmp19254;
  wire tmp19255;
  wire tmp19256;
  wire tmp19257;
  wire tmp19258;
  wire tmp19259;
  wire tmp19260;
  wire tmp19261;
  wire tmp19262;
  wire tmp19263;
  wire tmp19264;
  wire tmp19265;
  wire tmp19266;
  wire tmp19267;
  wire tmp19268;
  wire tmp19269;
  wire tmp19270;
  wire tmp19271;
  wire tmp19272;
  wire tmp19273;
  wire tmp19274;
  wire tmp19275;
  wire tmp19276;
  wire tmp19277;
  wire tmp19278;
  wire tmp19279;
  wire tmp19280;
  wire tmp19281;
  wire tmp19282;
  wire tmp19283;
  wire tmp19284;
  wire tmp19285;
  wire tmp19286;
  wire tmp19287;
  wire tmp19288;
  wire tmp19289;
  wire tmp19290;
  wire tmp19291;
  wire tmp19292;
  wire tmp19293;
  wire tmp19294;
  wire tmp19295;
  wire tmp19296;
  wire tmp19297;
  wire tmp19298;
  wire tmp19299;
  wire tmp19300;
  wire tmp19301;
  wire tmp19302;
  wire tmp19303;
  wire tmp19304;
  wire tmp19305;
  wire tmp19306;
  wire tmp19307;
  wire tmp19308;
  wire tmp19309;
  wire tmp19310;
  wire tmp19311;
  wire tmp19312;
  wire tmp19313;
  wire tmp19314;
  wire tmp19315;
  wire tmp19316;
  wire tmp19317;
  wire tmp19318;
  wire tmp19319;
  wire tmp19320;
  wire tmp19321;
  wire tmp19322;
  wire tmp19323;
  wire tmp19324;
  wire tmp19325;
  wire tmp19326;
  wire tmp19327;
  wire tmp19328;
  wire tmp19329;
  wire tmp19330;
  wire tmp19331;
  wire tmp19332;
  wire tmp19333;
  wire tmp19334;
  wire tmp19335;
  wire tmp19336;
  wire tmp19337;
  wire tmp19338;
  wire tmp19339;
  wire tmp19340;
  wire tmp19341;
  wire tmp19342;
  wire tmp19343;
  wire tmp19344;
  wire tmp19345;
  wire tmp19346;
  wire tmp19347;
  wire tmp19348;
  wire tmp19349;
  wire tmp19350;
  wire tmp19351;
  wire tmp19352;
  wire tmp19353;
  wire tmp19354;
  wire tmp19355;
  wire tmp19356;
  wire tmp19357;
  wire tmp19358;
  wire tmp19359;
  wire tmp19360;
  wire tmp19361;
  wire tmp19362;
  wire tmp19363;
  wire tmp19364;
  wire tmp19365;
  wire tmp19366;
  wire tmp19367;
  wire tmp19368;
  wire tmp19369;
  wire tmp19370;
  wire tmp19371;
  wire tmp19372;
  wire tmp19373;
  wire tmp19374;
  wire tmp19375;
  wire tmp19376;
  wire tmp19377;
  wire tmp19378;
  wire tmp19379;
  wire tmp19380;
  wire tmp19381;
  wire tmp19382;
  wire tmp19383;
  wire tmp19384;
  wire tmp19385;
  wire tmp19386;
  wire tmp19387;
  wire tmp19388;
  wire tmp19389;
  wire tmp19390;
  wire tmp19391;
  wire tmp19392;
  wire tmp19393;
  wire tmp19394;
  wire tmp19395;
  wire tmp19396;
  wire tmp19397;
  wire tmp19398;
  wire tmp19399;
  wire tmp19400;
  wire tmp19401;
  wire tmp19402;
  wire tmp19403;
  wire tmp19404;
  wire tmp19405;
  wire tmp19406;
  wire tmp19407;
  wire tmp19408;
  wire tmp19409;
  wire tmp19410;
  wire tmp19411;
  wire tmp19412;
  wire tmp19413;
  wire tmp19414;
  wire tmp19415;
  wire tmp19416;
  wire tmp19417;
  wire tmp19418;
  wire tmp19419;
  wire tmp19420;
  wire tmp19421;
  wire tmp19422;
  wire tmp19423;
  wire tmp19424;
  wire tmp19425;
  wire tmp19426;
  wire tmp19427;
  wire tmp19428;
  wire tmp19429;
  wire tmp19430;
  wire tmp19431;
  wire tmp19432;
  wire tmp19433;
  wire tmp19434;
  wire tmp19435;
  wire tmp19436;
  wire tmp19437;
  wire tmp19438;
  wire tmp19439;
  wire tmp19440;
  wire tmp19441;
  wire tmp19442;
  wire tmp19443;
  wire tmp19444;
  wire tmp19445;
  wire tmp19446;
  wire tmp19447;
  wire tmp19448;
  wire tmp19449;
  wire tmp19450;
  wire tmp19451;
  wire tmp19452;
  wire tmp19453;
  wire tmp19454;
  wire tmp19455;
  wire tmp19456;
  wire tmp19457;
  wire tmp19458;
  wire tmp19459;
  wire tmp19460;
  wire tmp19461;
  wire tmp19462;
  wire tmp19463;
  wire tmp19464;
  wire tmp19465;
  wire tmp19466;
  wire tmp19467;
  wire tmp19468;
  wire tmp19469;
  wire tmp19470;
  wire tmp19471;
  wire tmp19472;
  wire tmp19473;
  wire tmp19474;
  wire tmp19475;
  wire tmp19476;
  wire tmp19477;
  wire tmp19478;
  wire tmp19479;
  wire tmp19480;
  wire tmp19481;
  wire tmp19482;
  wire tmp19483;
  wire tmp19484;
  wire tmp19485;
  wire tmp19486;
  wire tmp19487;
  wire tmp19488;
  wire tmp19489;
  wire tmp19490;
  wire tmp19491;
  wire tmp19492;
  wire tmp19493;
  wire tmp19494;
  wire tmp19495;
  wire tmp19496;
  wire tmp19497;
  wire tmp19498;
  wire tmp19499;
  wire tmp19500;
  wire tmp19501;
  wire tmp19502;
  wire tmp19503;
  wire tmp19504;
  wire tmp19505;
  wire tmp19506;
  wire tmp19507;
  wire tmp19508;
  wire tmp19509;
  wire tmp19510;
  wire tmp19511;
  wire tmp19512;
  wire tmp19513;
  wire tmp19514;
  wire tmp19515;
  wire tmp19516;
  wire tmp19517;
  wire tmp19518;
  wire tmp19519;
  wire tmp19520;
  wire tmp19521;
  wire tmp19522;
  wire tmp19523;
  wire tmp19524;
  wire tmp19525;
  wire tmp19526;
  wire tmp19527;
  wire tmp19528;
  wire tmp19529;
  wire tmp19530;
  wire tmp19531;
  wire tmp19532;
  wire tmp19533;
  wire tmp19534;
  wire tmp19535;
  wire tmp19536;
  wire tmp19537;
  wire tmp19538;
  wire tmp19539;
  wire tmp19540;
  wire tmp19541;
  wire tmp19542;
  wire tmp19543;
  wire tmp19544;
  wire tmp19545;
  wire tmp19546;
  wire tmp19547;
  wire tmp19548;
  wire tmp19549;
  wire tmp19550;
  wire tmp19551;
  wire tmp19552;
  wire tmp19553;
  wire tmp19554;
  wire tmp19555;
  wire tmp19556;
  wire tmp19557;
  wire tmp19558;
  wire tmp19559;
  wire tmp19560;
  wire tmp19561;
  wire tmp19562;
  wire tmp19563;
  wire tmp19564;
  wire tmp19565;
  wire tmp19566;
  wire tmp19567;
  wire tmp19568;
  wire tmp19569;
  wire tmp19570;
  wire tmp19571;
  wire tmp19572;
  wire tmp19573;
  wire tmp19574;
  wire tmp19575;
  wire tmp19576;
  wire tmp19577;
  wire tmp19578;
  wire tmp19579;
  wire tmp19580;
  wire tmp19581;
  wire tmp19582;
  wire tmp19583;
  wire tmp19584;
  wire tmp19585;
  wire tmp19586;
  wire tmp19587;
  wire tmp19588;
  wire tmp19589;
  wire tmp19590;
  wire tmp19591;
  wire tmp19592;
  wire tmp19593;
  wire tmp19594;
  wire tmp19595;
  wire tmp19596;
  wire tmp19597;
  wire tmp19598;
  wire tmp19599;
  wire tmp19600;
  wire tmp19601;
  wire tmp19602;
  wire tmp19603;
  wire tmp19604;
  wire tmp19605;
  wire tmp19606;
  wire tmp19607;
  wire tmp19608;
  wire tmp19609;
  wire tmp19610;
  wire tmp19611;
  wire tmp19612;
  wire tmp19613;
  wire tmp19614;
  wire tmp19615;
  wire tmp19616;
  wire tmp19617;
  wire tmp19618;
  wire tmp19619;
  wire tmp19620;
  wire tmp19621;
  wire tmp19622;
  wire tmp19623;
  wire tmp19624;
  wire tmp19625;
  wire tmp19626;
  wire tmp19627;
  wire tmp19628;
  wire tmp19629;
  wire tmp19630;
  wire tmp19631;
  wire tmp19632;
  wire tmp19633;
  wire tmp19634;
  wire tmp19635;
  wire tmp19636;
  wire tmp19637;
  wire tmp19638;
  wire tmp19639;
  wire tmp19640;
  wire tmp19641;
  wire tmp19642;
  wire tmp19643;
  wire tmp19644;
  wire tmp19645;
  wire tmp19646;
  wire tmp19647;
  wire tmp19648;
  wire tmp19649;
  wire tmp19650;
  wire tmp19651;
  wire tmp19652;
  wire tmp19653;
  wire tmp19654;
  wire tmp19655;
  wire tmp19656;
  wire tmp19657;
  wire tmp19658;
  wire tmp19659;
  wire tmp19660;
  wire tmp19661;
  wire tmp19662;
  wire tmp19663;
  wire tmp19664;
  wire tmp19665;
  wire tmp19666;
  wire tmp19667;
  wire tmp19668;
  wire tmp19669;
  wire tmp19670;
  wire tmp19671;
  wire tmp19672;
  wire tmp19673;
  wire tmp19674;
  wire tmp19675;
  wire tmp19676;
  wire tmp19677;
  wire tmp19678;
  wire tmp19679;
  wire tmp19680;
  wire tmp19681;
  wire tmp19682;
  wire tmp19683;
  wire tmp19684;
  wire tmp19685;
  wire tmp19686;
  wire tmp19687;
  wire tmp19688;
  wire tmp19689;
  wire tmp19690;
  wire tmp19691;
  wire tmp19692;
  wire tmp19693;
  wire tmp19694;
  wire tmp19695;
  wire tmp19696;
  wire tmp19697;
  wire tmp19698;
  wire tmp19699;
  wire tmp19700;
  wire tmp19701;
  wire tmp19702;
  wire tmp19703;
  wire tmp19704;
  wire tmp19705;
  wire tmp19706;
  wire tmp19707;
  wire tmp19708;
  wire tmp19709;
  wire tmp19710;
  wire tmp19711;
  wire tmp19712;
  wire tmp19713;
  wire tmp19714;
  wire tmp19715;
  wire tmp19716;
  wire tmp19717;
  wire tmp19718;
  wire tmp19719;
  wire tmp19720;
  wire tmp19721;
  wire tmp19722;
  wire tmp19723;
  wire tmp19724;
  wire tmp19725;
  wire tmp19726;
  wire tmp19727;
  wire tmp19728;
  wire tmp19729;
  wire tmp19730;
  wire tmp19731;
  wire tmp19732;
  wire tmp19733;
  wire tmp19734;
  wire tmp19735;
  wire tmp19736;
  wire tmp19737;
  wire tmp19738;
  wire tmp19739;
  wire tmp19740;
  wire tmp19741;
  wire tmp19742;
  wire tmp19743;
  wire tmp19744;
  wire tmp19745;
  wire tmp19746;
  wire tmp19747;
  wire tmp19748;
  wire tmp19749;
  wire tmp19750;
  wire tmp19751;
  wire tmp19752;
  wire tmp19753;
  wire tmp19754;
  wire tmp19755;
  wire tmp19756;
  wire tmp19757;
  wire tmp19758;
  wire tmp19759;
  wire tmp19760;
  wire tmp19761;
  wire tmp19762;
  wire tmp19763;
  wire tmp19764;
  wire tmp19765;
  wire tmp19766;
  wire tmp19767;
  wire tmp19768;
  wire tmp19769;
  wire tmp19770;
  wire tmp19771;
  wire tmp19772;
  wire tmp19773;
  wire tmp19774;
  wire tmp19775;
  wire tmp19776;
  wire tmp19777;
  wire tmp19778;
  wire tmp19779;
  wire tmp19780;
  wire tmp19781;
  wire tmp19782;
  wire tmp19783;
  wire tmp19784;
  wire tmp19785;
  wire tmp19786;
  wire tmp19787;
  wire tmp19788;
  wire tmp19789;
  wire tmp19790;
  wire tmp19791;
  wire tmp19792;
  wire tmp19793;
  wire tmp19794;
  wire tmp19795;
  wire tmp19796;
  wire tmp19797;
  wire tmp19798;
  wire tmp19799;
  wire tmp19800;
  wire tmp19801;
  wire tmp19802;
  wire tmp19803;
  wire tmp19804;
  wire tmp19805;
  wire tmp19806;
  wire tmp19807;
  wire tmp19808;
  wire tmp19809;
  wire tmp19810;
  wire tmp19811;
  wire tmp19812;
  wire tmp19813;
  wire tmp19814;
  wire tmp19815;
  wire tmp19816;
  wire tmp19817;
  wire tmp19818;
  wire tmp19819;
  wire tmp19820;
  wire tmp19821;
  wire tmp19822;
  wire tmp19823;
  wire tmp19824;
  wire tmp19825;
  wire tmp19826;
  wire tmp19827;
  wire tmp19828;
  wire tmp19829;
  wire tmp19830;
  wire tmp19831;
  wire tmp19832;
  wire tmp19833;
  wire tmp19834;
  wire tmp19835;
  wire tmp19836;
  wire tmp19837;
  wire tmp19838;
  wire tmp19839;
  wire tmp19840;
  wire tmp19841;
  wire tmp19842;
  wire tmp19843;
  wire tmp19844;
  wire tmp19845;
  wire tmp19846;
  wire tmp19847;
  wire tmp19848;
  wire tmp19849;
  wire tmp19850;
  wire tmp19851;
  wire tmp19852;
  wire tmp19853;
  wire tmp19854;
  wire tmp19855;
  wire tmp19856;
  wire tmp19857;
  wire tmp19858;
  wire tmp19859;
  wire tmp19860;
  wire tmp19861;
  wire tmp19862;
  wire tmp19863;
  wire tmp19864;
  wire tmp19865;
  wire tmp19866;
  wire tmp19867;
  wire tmp19868;
  wire tmp19869;
  wire tmp19870;
  wire tmp19871;
  wire tmp19872;
  wire tmp19873;
  wire tmp19874;
  wire tmp19875;
  wire tmp19876;
  wire tmp19877;
  wire tmp19878;
  wire tmp19879;
  wire tmp19880;
  wire tmp19881;
  wire tmp19882;
  wire tmp19883;
  wire tmp19884;
  wire tmp19885;
  wire tmp19886;
  wire tmp19887;
  wire tmp19888;
  wire tmp19889;
  wire tmp19890;
  wire tmp19891;
  wire tmp19892;
  wire tmp19893;
  wire tmp19894;
  wire tmp19895;
  wire tmp19896;
  wire tmp19897;
  wire tmp19898;
  wire tmp19899;
  wire tmp19900;
  wire tmp19901;
  wire tmp19902;
  wire tmp19903;
  wire tmp19904;
  wire tmp19905;
  wire tmp19906;
  wire tmp19907;
  wire tmp19908;
  wire tmp19909;
  wire tmp19910;
  wire tmp19911;
  wire tmp19912;
  wire tmp19913;
  wire tmp19914;
  wire tmp19915;
  wire tmp19916;
  wire tmp19917;
  wire tmp19918;
  wire tmp19919;
  wire tmp19920;
  wire tmp19921;
  wire tmp19922;
  wire tmp19923;
  wire tmp19924;
  wire tmp19925;
  wire tmp19926;
  wire tmp19927;
  wire tmp19928;
  wire tmp19929;
  wire tmp19930;
  wire tmp19931;
  wire tmp19932;
  wire tmp19933;
  wire tmp19934;
  wire tmp19935;
  wire tmp19936;
  wire tmp19937;
  wire tmp19938;
  wire tmp19939;
  wire tmp19940;
  wire tmp19941;
  wire tmp19942;
  wire tmp19943;
  wire tmp19944;
  wire tmp19945;
  wire tmp19946;
  wire tmp19947;
  wire tmp19948;
  wire tmp19949;
  wire tmp19950;
  wire tmp19951;
  wire tmp19952;
  wire tmp19953;
  wire tmp19954;
  wire tmp19955;
  wire tmp19956;
  wire tmp19957;
  wire tmp19958;
  wire tmp19959;
  wire tmp19960;
  wire tmp19961;
  wire tmp19962;
  wire tmp19963;
  wire tmp19964;
  wire tmp19965;
  wire tmp19966;
  wire tmp19967;
  wire tmp19968;
  wire tmp19969;
  wire tmp19970;
  wire tmp19971;
  wire tmp19972;
  wire tmp19973;
  wire tmp19974;
  wire tmp19975;
  wire tmp19976;
  wire tmp19977;
  wire tmp19978;
  wire tmp19979;
  wire tmp19980;
  wire tmp19981;
  wire tmp19982;
  wire tmp19983;
  wire tmp19984;
  wire tmp19985;
  wire tmp19986;
  wire tmp19987;
  wire tmp19988;
  wire tmp19989;
  wire tmp19990;
  wire tmp19991;
  wire tmp19992;
  wire tmp19993;
  wire tmp19994;
  wire tmp19995;
  wire tmp19996;
  wire tmp19997;
  wire tmp19998;
  wire tmp19999;
  wire tmp20000;
  wire tmp20001;
  wire tmp20002;
  wire tmp20003;
  wire tmp20004;
  wire tmp20005;
  wire tmp20006;
  wire tmp20007;
  wire tmp20008;
  wire tmp20009;
  wire tmp20010;
  wire tmp20011;
  wire tmp20012;
  wire tmp20013;
  wire tmp20014;
  wire tmp20015;
  wire tmp20016;
  wire tmp20017;
  wire tmp20018;
  wire tmp20019;
  wire tmp20020;
  wire tmp20021;
  wire tmp20022;
  wire tmp20023;
  wire tmp20024;
  wire tmp20025;
  wire tmp20026;
  wire tmp20027;
  wire tmp20028;
  wire tmp20029;
  wire tmp20030;
  wire tmp20031;
  wire tmp20032;
  wire tmp20033;
  wire tmp20034;
  wire tmp20035;
  wire tmp20036;
  wire tmp20037;
  wire tmp20038;
  wire tmp20039;
  wire tmp20040;
  wire tmp20041;
  wire tmp20042;
  wire tmp20043;
  wire tmp20044;
  wire tmp20045;
  wire tmp20046;
  wire tmp20047;
  wire tmp20048;
  wire tmp20049;
  wire tmp20050;
  wire tmp20051;
  wire tmp20052;
  wire tmp20053;
  wire tmp20054;
  wire tmp20055;
  wire tmp20056;
  wire tmp20057;
  wire tmp20058;
  wire tmp20059;
  wire tmp20060;
  wire tmp20061;
  wire tmp20062;
  wire tmp20063;
  wire tmp20064;
  wire tmp20065;
  wire tmp20066;
  wire tmp20067;
  wire tmp20068;
  wire tmp20069;
  wire tmp20070;
  wire tmp20071;
  wire tmp20072;
  wire tmp20073;
  wire tmp20074;
  wire tmp20075;
  wire tmp20076;
  wire tmp20077;
  wire tmp20078;
  wire tmp20079;
  wire tmp20080;
  wire tmp20081;
  wire tmp20082;
  wire tmp20083;
  wire tmp20084;
  wire tmp20085;
  wire tmp20086;
  wire tmp20087;
  wire tmp20088;
  wire tmp20089;
  wire tmp20090;
  wire tmp20091;
  wire tmp20092;
  wire tmp20093;
  wire tmp20094;
  wire tmp20095;
  wire tmp20096;
  wire tmp20097;
  wire tmp20098;
  wire tmp20099;
  wire tmp20100;
  wire tmp20101;
  wire tmp20102;
  wire tmp20103;
  wire tmp20104;
  wire tmp20105;
  wire tmp20106;
  wire tmp20107;
  wire tmp20108;
  wire tmp20109;
  wire tmp20110;
  wire tmp20111;
  wire tmp20112;
  wire tmp20113;
  wire tmp20114;
  wire tmp20115;
  wire tmp20116;
  wire tmp20117;
  wire tmp20118;
  wire tmp20119;
  wire tmp20120;
  wire tmp20121;
  wire tmp20122;
  wire tmp20123;
  wire tmp20124;
  wire tmp20125;
  wire tmp20126;
  wire tmp20127;
  wire tmp20128;
  wire tmp20129;
  wire tmp20130;
  wire tmp20131;
  wire tmp20132;
  wire tmp20133;
  wire tmp20134;
  wire tmp20135;
  wire tmp20136;
  wire tmp20137;
  wire tmp20138;
  wire tmp20139;
  wire tmp20140;
  wire tmp20141;
  wire tmp20142;
  wire tmp20143;
  wire tmp20144;
  wire tmp20145;
  wire tmp20146;
  wire tmp20147;
  wire tmp20148;
  wire tmp20149;
  wire tmp20150;
  wire tmp20151;
  wire tmp20152;
  wire tmp20153;
  wire tmp20154;
  wire tmp20155;
  wire tmp20156;
  wire tmp20157;
  wire tmp20158;
  wire tmp20159;
  wire tmp20160;
  wire tmp20161;
  wire tmp20162;
  wire tmp20163;
  wire tmp20164;
  wire tmp20165;
  wire tmp20166;
  wire tmp20167;
  wire tmp20168;
  wire tmp20169;
  wire tmp20170;
  wire tmp20171;
  wire tmp20172;
  wire tmp20173;
  wire tmp20174;
  wire tmp20175;
  wire tmp20176;
  wire tmp20177;
  wire tmp20178;
  wire tmp20179;
  wire tmp20180;
  wire tmp20181;
  wire tmp20182;
  wire tmp20183;
  wire tmp20184;
  wire tmp20185;
  wire tmp20186;
  wire tmp20187;
  wire tmp20188;
  wire tmp20189;
  wire tmp20190;
  wire tmp20191;
  wire tmp20192;
  wire tmp20193;
  wire tmp20194;
  wire tmp20195;
  wire tmp20196;
  wire tmp20197;
  wire tmp20198;
  wire tmp20199;
  wire tmp20200;
  wire tmp20201;
  wire tmp20202;
  wire tmp20203;
  wire tmp20204;
  wire tmp20205;
  wire tmp20206;
  wire tmp20207;
  wire tmp20208;
  wire tmp20209;
  wire tmp20210;
  wire tmp20211;
  wire tmp20212;
  wire tmp20213;
  wire tmp20214;
  wire tmp20215;
  wire tmp20216;
  wire tmp20217;
  wire tmp20218;
  wire tmp20219;
  wire tmp20220;
  wire tmp20221;
  wire tmp20222;
  wire tmp20223;
  wire tmp20224;
  wire tmp20225;
  wire tmp20226;
  wire tmp20227;
  wire tmp20228;
  wire tmp20229;
  wire tmp20230;
  wire tmp20231;
  wire tmp20232;
  wire tmp20233;
  wire tmp20234;
  wire tmp20235;
  wire tmp20236;
  wire tmp20237;
  wire tmp20238;
  wire tmp20239;
  wire tmp20240;
  wire tmp20241;
  wire tmp20242;
  wire tmp20243;
  wire tmp20244;
  wire tmp20245;
  wire tmp20246;
  wire tmp20247;
  wire tmp20248;
  wire tmp20249;
  wire tmp20250;
  wire tmp20251;
  wire tmp20252;
  wire tmp20253;
  wire tmp20254;
  wire tmp20255;
  wire tmp20256;
  wire tmp20257;
  wire tmp20258;
  wire tmp20259;
  wire tmp20260;
  wire tmp20261;
  wire tmp20262;
  wire tmp20263;
  wire tmp20264;
  wire tmp20265;
  wire tmp20266;
  wire tmp20267;
  wire tmp20268;
  wire tmp20269;
  wire tmp20270;
  wire tmp20271;
  wire tmp20272;
  wire tmp20273;
  wire tmp20274;
  wire tmp20275;
  wire tmp20276;
  wire tmp20277;
  wire tmp20278;
  wire tmp20279;
  wire tmp20280;
  wire tmp20281;
  wire tmp20282;
  wire tmp20283;
  wire tmp20284;
  wire tmp20285;
  wire tmp20286;
  wire tmp20287;
  wire tmp20288;
  wire tmp20289;
  wire tmp20290;
  wire tmp20291;
  wire tmp20292;
  wire tmp20293;
  wire tmp20294;
  wire tmp20295;
  wire tmp20296;
  wire tmp20297;
  wire tmp20298;
  wire tmp20299;
  wire tmp20300;
  wire tmp20301;
  wire tmp20302;
  wire tmp20303;
  wire tmp20304;
  wire tmp20305;
  wire tmp20306;
  wire tmp20307;
  wire tmp20308;
  wire tmp20309;
  wire tmp20310;
  wire tmp20311;
  wire tmp20312;
  wire tmp20313;
  wire tmp20314;
  wire tmp20315;
  wire tmp20316;
  wire tmp20317;
  wire tmp20318;
  wire tmp20319;
  wire tmp20320;
  wire tmp20321;
  wire tmp20322;
  wire tmp20323;
  wire tmp20324;
  wire tmp20325;
  wire tmp20326;
  wire tmp20327;
  wire tmp20328;
  wire tmp20329;
  wire tmp20330;
  wire tmp20331;
  wire tmp20332;
  wire tmp20333;
  wire tmp20334;
  wire tmp20335;
  wire tmp20336;
  wire tmp20337;
  wire tmp20338;
  wire tmp20339;
  wire tmp20340;
  wire tmp20341;
  wire tmp20342;
  wire tmp20343;
  wire tmp20344;
  wire tmp20345;
  wire tmp20346;
  wire tmp20347;
  wire tmp20348;
  wire tmp20349;
  wire tmp20350;
  wire tmp20351;
  wire tmp20352;
  wire tmp20353;
  wire tmp20354;
  wire tmp20355;
  wire tmp20356;
  wire tmp20357;
  wire tmp20358;
  wire tmp20359;
  wire tmp20360;
  wire tmp20361;
  wire tmp20362;
  wire tmp20363;
  wire tmp20364;
  wire tmp20365;
  wire tmp20366;
  wire tmp20367;
  wire tmp20368;
  wire tmp20369;
  wire tmp20370;
  wire tmp20371;
  wire tmp20372;
  wire tmp20373;
  wire tmp20374;
  wire tmp20375;
  wire tmp20376;
  wire tmp20377;
  wire tmp20378;
  wire tmp20379;
  wire tmp20380;
  wire tmp20381;
  wire tmp20382;
  wire tmp20383;
  wire tmp20384;
  wire tmp20385;
  wire tmp20386;
  wire tmp20387;
  wire tmp20388;
  wire tmp20389;
  wire tmp20390;
  wire tmp20391;
  wire tmp20392;
  wire tmp20393;
  wire tmp20394;
  wire tmp20395;
  wire tmp20396;
  wire tmp20397;
  wire tmp20398;
  wire tmp20399;
  wire tmp20400;
  wire tmp20401;
  wire tmp20402;
  wire tmp20403;
  wire tmp20404;
  wire tmp20405;
  wire tmp20406;
  wire tmp20407;
  wire tmp20408;
  wire tmp20409;
  wire tmp20410;
  wire tmp20411;
  wire tmp20412;
  wire tmp20413;
  wire tmp20414;
  wire tmp20415;
  wire tmp20416;
  wire tmp20417;
  wire tmp20418;
  wire tmp20419;
  wire tmp20420;
  wire tmp20421;
  wire tmp20422;
  wire tmp20423;
  wire tmp20424;
  wire tmp20425;
  wire tmp20426;
  wire tmp20427;
  wire tmp20428;
  wire tmp20429;
  wire tmp20430;
  wire tmp20431;
  wire tmp20432;
  wire tmp20433;
  wire tmp20434;
  wire tmp20435;
  wire tmp20436;
  wire tmp20437;
  wire tmp20438;
  wire tmp20439;
  wire tmp20440;
  wire tmp20441;
  wire tmp20442;
  wire tmp20443;
  wire tmp20444;
  wire tmp20445;
  wire tmp20446;
  wire tmp20447;
  wire tmp20448;
  wire tmp20449;
  wire tmp20450;
  wire tmp20451;
  wire tmp20452;
  wire tmp20453;
  wire tmp20454;
  wire tmp20455;
  wire tmp20456;
  wire tmp20457;
  wire tmp20458;
  wire tmp20459;
  wire tmp20460;
  wire tmp20461;
  wire tmp20462;
  wire tmp20463;
  wire tmp20464;
  wire tmp20465;
  wire tmp20466;
  wire tmp20467;
  wire tmp20468;
  wire tmp20469;
  wire tmp20470;
  wire tmp20471;
  wire tmp20472;
  wire tmp20473;
  wire tmp20474;
  wire tmp20475;
  wire tmp20476;
  wire tmp20477;
  wire tmp20478;
  wire tmp20479;
  wire tmp20480;
  wire tmp20481;
  wire tmp20482;
  wire tmp20483;
  wire tmp20484;
  wire tmp20485;
  wire tmp20486;
  wire tmp20487;
  wire tmp20488;
  wire tmp20489;
  wire tmp20490;
  wire tmp20491;
  wire tmp20492;
  wire tmp20493;
  wire tmp20494;
  wire tmp20495;
  wire tmp20496;
  wire tmp20497;
  wire tmp20498;
  wire tmp20499;
  wire tmp20500;
  wire tmp20501;
  wire tmp20502;
  wire tmp20503;
  wire tmp20504;
  wire tmp20505;
  wire tmp20506;
  wire tmp20507;
  wire tmp20508;
  wire tmp20509;
  wire tmp20510;
  wire tmp20511;
  wire tmp20512;
  wire tmp20513;
  wire tmp20514;
  wire tmp20515;
  wire tmp20516;
  wire tmp20517;
  wire tmp20518;
  wire tmp20519;
  wire tmp20520;
  wire tmp20521;
  wire tmp20522;
  wire tmp20523;
  wire tmp20524;
  wire tmp20525;
  wire tmp20526;
  wire tmp20527;
  wire tmp20528;
  wire tmp20529;
  wire tmp20530;
  wire tmp20531;
  wire tmp20532;
  wire tmp20533;
  wire tmp20534;
  wire tmp20535;
  wire tmp20536;
  wire tmp20537;
  wire tmp20538;
  wire tmp20539;
  wire tmp20540;
  wire tmp20541;
  wire tmp20542;
  wire tmp20543;
  wire tmp20544;
  wire tmp20545;
  wire tmp20546;
  wire tmp20547;
  wire tmp20548;
  wire tmp20549;
  wire tmp20550;
  wire tmp20551;
  wire tmp20552;
  wire tmp20553;
  wire tmp20554;
  wire tmp20555;
  wire tmp20556;
  wire tmp20557;
  wire tmp20558;
  wire tmp20559;
  wire tmp20560;
  wire tmp20561;
  wire tmp20562;
  wire tmp20563;
  wire tmp20564;
  wire tmp20565;
  wire tmp20566;
  wire tmp20567;
  wire tmp20568;
  wire tmp20569;
  wire tmp20570;
  wire tmp20571;
  wire tmp20572;
  wire tmp20573;
  wire tmp20574;
  wire tmp20575;
  wire tmp20576;
  wire tmp20577;
  wire tmp20578;
  wire tmp20579;
  wire tmp20580;
  wire tmp20581;
  wire tmp20582;
  wire tmp20583;
  wire tmp20584;
  wire tmp20585;
  wire tmp20586;
  wire tmp20587;
  wire tmp20588;
  wire tmp20589;
  wire tmp20590;
  wire tmp20591;
  wire tmp20592;
  wire tmp20593;
  wire tmp20594;
  wire tmp20595;
  wire tmp20596;
  wire tmp20597;
  wire tmp20598;
  wire tmp20599;
  wire tmp20600;
  wire tmp20601;
  wire tmp20602;
  wire tmp20603;
  wire tmp20604;
  wire tmp20605;
  wire tmp20606;
  wire tmp20607;
  wire tmp20608;
  wire tmp20609;
  wire tmp20610;
  wire tmp20611;
  wire tmp20612;
  wire tmp20613;
  wire tmp20614;
  wire tmp20615;
  wire tmp20616;
  wire tmp20617;
  wire tmp20618;
  wire tmp20619;
  wire tmp20620;
  wire tmp20621;
  wire tmp20622;
  wire tmp20623;
  wire tmp20624;
  wire tmp20625;
  wire tmp20626;
  wire tmp20627;
  wire tmp20628;
  wire tmp20629;
  wire tmp20630;
  wire tmp20631;
  wire tmp20632;
  wire tmp20633;
  wire tmp20634;
  wire tmp20635;
  wire tmp20636;
  wire tmp20637;
  wire tmp20638;
  wire tmp20639;
  wire tmp20640;
  wire tmp20641;
  wire tmp20642;
  wire tmp20643;
  wire tmp20644;
  wire tmp20645;
  wire tmp20646;
  wire tmp20647;
  wire tmp20648;
  wire tmp20649;
  wire tmp20650;
  wire tmp20651;
  wire tmp20652;
  wire tmp20653;
  wire tmp20654;
  wire tmp20655;
  wire tmp20656;
  wire tmp20657;
  wire tmp20658;
  wire tmp20659;
  wire tmp20660;
  wire tmp20661;
  wire tmp20662;
  wire tmp20663;
  wire tmp20664;
  wire tmp20665;
  wire tmp20666;
  wire tmp20667;
  wire tmp20668;
  wire tmp20669;
  wire tmp20670;
  wire tmp20671;
  wire tmp20672;
  wire tmp20673;
  wire tmp20674;
  wire tmp20675;
  wire tmp20676;
  wire tmp20677;
  wire tmp20678;
  wire tmp20679;
  wire tmp20680;
  wire tmp20681;
  wire tmp20682;
  wire tmp20683;
  wire tmp20684;
  wire tmp20685;
  wire tmp20686;
  wire tmp20687;
  wire tmp20688;
  wire tmp20689;
  wire tmp20690;
  wire tmp20691;
  wire tmp20692;
  wire tmp20693;
  wire tmp20694;
  wire tmp20695;
  wire tmp20696;
  wire tmp20697;
  wire tmp20698;
  wire tmp20699;
  wire tmp20700;
  wire tmp20701;
  wire tmp20702;
  wire tmp20703;
  wire tmp20704;
  wire tmp20705;
  wire tmp20706;
  wire tmp20707;
  wire tmp20708;
  wire tmp20709;
  wire tmp20710;
  wire tmp20711;
  wire tmp20712;
  wire tmp20713;
  wire tmp20714;
  wire tmp20715;
  wire tmp20716;
  wire tmp20717;
  wire tmp20718;
  wire tmp20719;
  wire tmp20720;
  wire tmp20721;
  wire tmp20722;
  wire tmp20723;
  wire tmp20724;
  wire tmp20725;
  wire tmp20726;
  wire tmp20727;
  wire tmp20728;
  wire tmp20729;
  wire tmp20730;
  wire tmp20731;
  wire tmp20732;
  wire tmp20733;
  wire tmp20734;
  wire tmp20735;
  wire tmp20736;
  wire tmp20737;
  wire tmp20738;
  wire tmp20739;
  wire tmp20740;
  wire tmp20741;
  wire tmp20742;
  wire tmp20743;
  wire tmp20744;
  wire tmp20745;
  wire tmp20746;
  wire tmp20747;
  wire tmp20748;
  wire tmp20749;
  wire tmp20750;
  wire tmp20751;
  wire tmp20752;
  wire tmp20753;
  wire tmp20754;
  wire tmp20755;
  wire tmp20756;
  wire tmp20757;
  wire tmp20758;
  wire tmp20759;
  wire tmp20760;
  wire tmp20761;
  wire tmp20762;
  wire tmp20763;
  wire tmp20764;
  wire tmp20765;
  wire tmp20766;
  wire tmp20767;
  wire tmp20768;
  wire tmp20769;
  wire tmp20770;
  wire tmp20771;
  wire tmp20772;
  wire tmp20773;
  wire tmp20774;
  wire tmp20775;
  wire tmp20776;
  wire tmp20777;
  wire tmp20778;
  wire tmp20779;
  wire tmp20780;
  wire tmp20781;
  wire tmp20782;
  wire tmp20783;
  wire tmp20784;
  wire tmp20785;
  wire tmp20786;
  wire tmp20787;
  wire tmp20788;
  wire tmp20789;
  wire tmp20790;
  wire tmp20791;
  wire tmp20792;
  wire tmp20793;
  wire tmp20794;
  wire tmp20795;
  wire tmp20796;
  wire tmp20797;
  wire tmp20798;
  wire tmp20799;
  wire tmp20800;
  wire tmp20801;
  wire tmp20802;
  wire tmp20803;
  wire tmp20804;
  wire tmp20805;
  wire tmp20806;
  wire tmp20807;
  wire tmp20808;
  wire tmp20809;
  wire tmp20810;
  wire tmp20811;
  wire tmp20812;
  wire tmp20813;
  wire tmp20814;
  wire tmp20815;
  wire tmp20816;
  wire tmp20817;
  wire tmp20818;
  wire tmp20819;
  wire tmp20820;
  wire tmp20821;
  wire tmp20822;
  wire tmp20823;
  wire tmp20824;
  wire tmp20825;
  wire tmp20826;
  wire tmp20827;
  wire tmp20828;
  wire tmp20829;
  wire tmp20830;
  wire tmp20831;
  wire tmp20832;
  wire tmp20833;
  wire tmp20834;
  wire tmp20835;
  wire tmp20836;
  wire tmp20837;
  wire tmp20838;
  wire tmp20839;
  wire tmp20840;
  wire tmp20841;
  wire tmp20842;
  wire tmp20843;
  wire tmp20844;
  wire tmp20845;
  wire tmp20846;
  wire tmp20847;
  wire tmp20848;
  wire tmp20849;
  wire tmp20850;
  wire tmp20851;
  wire tmp20852;
  wire tmp20853;
  wire tmp20854;
  wire tmp20855;
  wire tmp20856;
  wire tmp20857;
  wire tmp20858;
  wire tmp20859;
  wire tmp20860;
  wire tmp20861;
  wire tmp20862;
  wire tmp20863;
  wire tmp20864;
  wire tmp20865;
  wire tmp20866;
  wire tmp20867;
  wire tmp20868;
  wire tmp20869;
  wire tmp20870;
  wire tmp20871;
  wire tmp20872;
  wire tmp20873;
  wire tmp20874;
  wire tmp20875;
  wire tmp20876;
  wire tmp20877;
  wire tmp20878;
  wire tmp20879;
  wire tmp20880;
  wire tmp20881;
  wire tmp20882;
  wire tmp20883;
  wire tmp20884;
  wire tmp20885;
  wire tmp20886;
  wire tmp20887;
  wire tmp20888;
  wire tmp20889;
  wire tmp20890;
  wire tmp20891;
  wire tmp20892;
  wire tmp20893;
  wire tmp20894;
  wire tmp20895;
  wire tmp20896;
  wire tmp20897;
  wire tmp20898;
  wire tmp20899;
  wire tmp20900;
  wire tmp20901;
  wire tmp20902;
  wire tmp20903;
  wire tmp20904;
  wire tmp20905;
  wire tmp20906;
  wire tmp20907;
  wire tmp20908;
  wire tmp20909;
  wire tmp20910;
  wire tmp20911;
  wire tmp20912;
  wire tmp20913;
  wire tmp20914;
  wire tmp20915;
  wire tmp20916;
  wire tmp20917;
  wire tmp20918;
  wire tmp20919;
  wire tmp20920;
  wire tmp20921;
  wire tmp20922;
  wire tmp20923;
  wire tmp20924;
  wire tmp20925;
  wire tmp20926;
  wire tmp20927;
  wire tmp20928;
  wire tmp20929;
  wire tmp20930;
  wire tmp20931;
  wire tmp20932;
  wire tmp20933;
  wire tmp20934;
  wire tmp20935;
  wire tmp20936;
  wire tmp20937;
  wire tmp20938;
  wire tmp20939;
  wire tmp20940;
  wire tmp20941;
  wire tmp20942;
  wire tmp20943;
  wire tmp20944;
  wire tmp20945;
  wire tmp20946;
  wire tmp20947;
  wire tmp20948;
  wire tmp20949;
  wire tmp20950;
  wire tmp20951;
  wire tmp20952;
  wire tmp20953;
  wire tmp20954;
  wire tmp20955;
  wire tmp20956;
  wire tmp20957;
  wire tmp20958;
  wire tmp20959;
  wire tmp20960;
  wire tmp20961;
  wire tmp20962;
  wire tmp20963;
  wire tmp20964;
  wire tmp20965;
  wire tmp20966;
  wire tmp20967;
  wire tmp20968;
  wire tmp20969;
  wire tmp20970;
  wire tmp20971;
  wire tmp20972;
  wire tmp20973;
  wire tmp20974;
  wire tmp20975;
  wire tmp20976;
  wire tmp20977;
  wire tmp20978;
  wire tmp20979;
  wire tmp20980;
  wire tmp20981;
  wire tmp20982;
  wire tmp20983;
  wire tmp20984;
  wire tmp20985;
  wire tmp20986;
  wire tmp20987;
  wire tmp20988;
  wire tmp20989;
  wire tmp20990;
  wire tmp20991;
  wire tmp20992;
  wire tmp20993;
  wire tmp20994;
  wire tmp20995;
  wire tmp20996;
  wire tmp20997;
  wire tmp20998;
  wire tmp20999;
  wire tmp21000;
  wire tmp21001;
  wire tmp21002;
  wire tmp21003;
  wire tmp21004;
  wire tmp21005;
  wire tmp21006;
  wire tmp21007;
  wire tmp21008;
  wire tmp21009;
  wire tmp21010;
  wire tmp21011;
  wire tmp21012;
  wire tmp21013;
  wire tmp21014;
  wire tmp21015;
  wire tmp21016;
  wire tmp21017;
  wire tmp21018;
  wire tmp21019;
  wire tmp21020;
  wire tmp21021;
  wire tmp21022;
  wire tmp21023;
  wire tmp21024;
  wire tmp21025;
  wire tmp21026;
  wire tmp21027;
  wire tmp21028;
  wire tmp21029;
  wire tmp21030;
  wire tmp21031;
  wire tmp21032;
  wire tmp21033;
  wire tmp21034;
  wire tmp21035;
  wire tmp21036;
  wire tmp21037;
  wire tmp21038;
  wire tmp21039;
  wire tmp21040;
  wire tmp21041;
  wire tmp21042;
  wire tmp21043;
  wire tmp21044;
  wire tmp21045;
  wire tmp21046;
  wire tmp21047;
  wire tmp21048;
  wire tmp21049;
  wire tmp21050;
  wire tmp21051;
  wire tmp21052;
  wire tmp21053;
  wire tmp21054;
  wire tmp21055;
  wire tmp21056;
  wire tmp21057;
  wire tmp21058;
  wire tmp21059;
  wire tmp21060;
  wire tmp21061;
  wire tmp21062;
  wire tmp21063;
  wire tmp21064;
  wire tmp21065;
  wire tmp21066;
  wire tmp21067;
  wire tmp21068;
  wire tmp21069;
  wire tmp21070;
  wire tmp21071;
  wire tmp21072;
  wire tmp21073;
  wire tmp21074;
  wire tmp21075;
  wire tmp21076;
  wire tmp21077;
  wire tmp21078;
  wire tmp21079;
  wire tmp21080;
  wire tmp21081;
  wire tmp21082;
  wire tmp21083;
  wire tmp21084;
  wire tmp21085;
  wire tmp21086;
  wire tmp21087;
  wire tmp21088;
  wire tmp21089;
  wire tmp21090;
  wire tmp21091;
  wire tmp21092;
  wire tmp21093;
  wire tmp21094;
  wire tmp21095;
  wire tmp21096;
  wire tmp21097;
  wire tmp21098;
  wire tmp21099;
  wire tmp21100;
  wire tmp21101;
  wire tmp21102;
  wire tmp21103;
  wire tmp21104;
  wire tmp21105;
  wire tmp21106;
  wire tmp21107;
  wire tmp21108;
  wire tmp21109;
  wire tmp21110;
  wire tmp21111;
  wire tmp21112;
  wire tmp21113;
  wire tmp21114;
  wire tmp21115;
  wire tmp21116;
  wire tmp21117;
  wire tmp21118;
  wire tmp21119;
  wire tmp21120;
  wire tmp21121;
  wire tmp21122;
  wire tmp21123;
  wire tmp21124;
  wire tmp21125;
  wire tmp21126;
  wire tmp21127;
  wire tmp21128;
  wire tmp21129;
  wire tmp21130;
  wire tmp21131;
  wire tmp21132;
  wire tmp21133;
  wire tmp21134;
  wire tmp21135;
  wire tmp21136;
  wire tmp21137;
  wire tmp21138;
  wire tmp21139;
  wire tmp21140;
  wire tmp21141;
  wire tmp21142;
  wire tmp21143;
  wire tmp21144;
  wire tmp21145;
  wire tmp21146;
  wire tmp21147;
  wire tmp21148;
  wire tmp21149;
  wire tmp21150;
  wire tmp21151;
  wire tmp21152;
  wire tmp21153;
  wire tmp21154;
  wire tmp21155;
  wire tmp21156;
  wire tmp21157;
  wire tmp21158;
  wire tmp21159;
  wire tmp21160;
  wire tmp21161;
  wire tmp21162;
  wire tmp21163;
  wire tmp21164;
  wire tmp21165;
  wire tmp21166;
  wire tmp21167;
  wire tmp21168;
  wire tmp21169;
  wire tmp21170;
  wire tmp21171;
  wire tmp21172;
  wire tmp21173;
  wire tmp21174;
  wire tmp21175;
  wire tmp21176;
  wire tmp21177;
  wire tmp21178;
  wire tmp21179;
  wire tmp21180;
  wire tmp21181;
  wire tmp21182;
  wire tmp21183;
  wire tmp21184;
  wire tmp21185;
  wire tmp21186;
  wire tmp21187;
  wire tmp21188;
  wire tmp21189;
  wire tmp21190;
  wire tmp21191;
  wire tmp21192;
  wire tmp21193;
  wire tmp21194;
  wire tmp21195;
  wire tmp21196;
  wire tmp21197;
  wire tmp21198;
  wire tmp21199;
  wire tmp21200;
  wire tmp21201;
  wire tmp21202;
  wire tmp21203;
  wire tmp21204;
  wire tmp21205;
  wire tmp21206;
  wire tmp21207;
  wire tmp21208;
  wire tmp21209;
  wire tmp21210;
  wire tmp21211;
  wire tmp21212;
  wire tmp21213;
  wire tmp21214;
  wire tmp21215;
  wire tmp21216;
  wire tmp21217;
  wire tmp21218;
  wire tmp21219;
  wire tmp21220;
  wire tmp21221;
  wire tmp21222;
  wire tmp21223;
  wire tmp21224;
  wire tmp21225;
  wire tmp21226;
  wire tmp21227;
  wire tmp21228;
  wire tmp21229;
  wire tmp21230;
  wire tmp21231;
  wire tmp21232;
  wire tmp21233;
  wire tmp21234;
  wire tmp21235;
  wire tmp21236;
  wire tmp21237;
  wire tmp21238;
  wire tmp21239;
  wire tmp21240;
  wire tmp21241;
  wire tmp21242;
  wire tmp21243;
  wire tmp21244;
  wire tmp21245;
  wire tmp21246;
  wire tmp21247;
  wire tmp21248;
  wire tmp21249;
  wire tmp21250;
  wire tmp21251;
  wire tmp21252;
  wire tmp21253;
  wire tmp21254;
  wire tmp21255;
  wire tmp21256;
  wire tmp21257;
  wire tmp21258;
  wire tmp21259;
  wire tmp21260;
  wire tmp21261;
  wire tmp21262;
  wire tmp21263;
  wire tmp21264;
  wire tmp21265;
  wire tmp21266;
  wire tmp21267;
  wire tmp21268;
  wire tmp21269;
  wire tmp21270;
  wire tmp21271;
  wire tmp21272;
  wire tmp21273;
  wire tmp21274;
  wire tmp21275;
  wire tmp21276;
  wire tmp21277;
  wire tmp21278;
  wire tmp21279;
  wire tmp21280;
  wire tmp21281;
  wire tmp21282;
  wire tmp21283;
  wire tmp21284;
  wire tmp21285;
  wire tmp21286;
  wire tmp21287;
  wire tmp21288;
  wire tmp21289;
  wire tmp21290;
  wire tmp21291;
  wire tmp21292;
  wire tmp21293;
  wire tmp21294;
  wire tmp21295;
  wire tmp21296;
  wire tmp21297;
  wire tmp21298;
  wire tmp21299;
  wire tmp21300;
  wire tmp21301;
  wire tmp21302;
  wire tmp21303;
  wire tmp21304;
  wire tmp21305;
  wire tmp21306;
  wire tmp21307;
  wire tmp21308;
  wire tmp21309;
  wire tmp21310;
  wire tmp21311;
  wire tmp21312;
  wire tmp21313;
  wire tmp21314;
  wire tmp21315;
  wire tmp21316;
  wire tmp21317;
  wire tmp21318;
  wire tmp21319;
  wire tmp21320;
  wire tmp21321;
  wire tmp21322;
  wire tmp21323;
  wire tmp21324;
  wire tmp21325;
  wire tmp21326;
  wire tmp21327;
  wire tmp21328;
  wire tmp21329;
  wire tmp21330;
  wire tmp21331;
  wire tmp21332;
  wire tmp21333;
  wire tmp21334;
  wire tmp21335;
  wire tmp21336;
  wire tmp21337;
  wire tmp21338;
  wire tmp21339;
  wire tmp21340;
  wire tmp21341;
  wire tmp21342;
  wire tmp21343;
  wire tmp21344;
  wire tmp21345;
  wire tmp21346;
  wire tmp21347;
  wire tmp21348;
  wire tmp21349;
  wire tmp21350;
  wire tmp21351;
  wire tmp21352;
  wire tmp21353;
  wire tmp21354;
  wire tmp21355;
  wire tmp21356;
  wire tmp21357;
  wire tmp21358;
  wire tmp21359;
  wire tmp21360;
  wire tmp21361;
  wire tmp21362;
  wire tmp21363;
  wire tmp21364;
  wire tmp21365;
  wire tmp21366;
  wire tmp21367;
  wire tmp21368;
  wire tmp21369;
  wire tmp21370;
  wire tmp21371;
  wire tmp21372;
  wire tmp21373;
  wire tmp21374;
  wire tmp21375;
  wire tmp21376;
  wire tmp21377;
  wire tmp21378;
  wire tmp21379;
  wire tmp21380;
  wire tmp21381;
  wire tmp21382;
  wire tmp21383;
  wire tmp21384;
  wire tmp21385;
  wire tmp21386;
  wire tmp21387;
  wire tmp21388;
  wire tmp21389;
  wire tmp21390;
  wire tmp21391;
  wire tmp21392;
  wire tmp21393;
  wire tmp21394;
  wire tmp21395;
  wire tmp21396;
  wire tmp21397;
  wire tmp21398;
  wire tmp21399;
  wire tmp21400;
  wire tmp21401;
  wire tmp21402;
  wire tmp21403;
  wire tmp21404;
  wire tmp21405;
  wire tmp21406;
  wire tmp21407;
  wire tmp21408;
  wire tmp21409;
  wire tmp21410;
  wire tmp21411;
  wire tmp21412;
  wire tmp21413;
  wire tmp21414;
  wire tmp21415;
  wire tmp21416;
  wire tmp21417;
  wire tmp21418;
  wire tmp21419;
  wire tmp21420;
  wire tmp21421;
  wire tmp21422;
  wire tmp21423;
  wire tmp21424;
  wire tmp21425;
  wire tmp21426;
  wire tmp21427;
  wire tmp21428;
  wire tmp21429;
  wire tmp21430;
  wire tmp21431;
  wire tmp21432;
  wire tmp21433;
  wire tmp21434;
  wire tmp21435;
  wire tmp21436;
  wire tmp21437;
  wire tmp21438;
  wire tmp21439;
  wire tmp21440;
  wire tmp21441;
  wire tmp21442;
  wire tmp21443;
  wire tmp21444;
  wire tmp21445;
  wire tmp21446;
  wire tmp21447;
  wire tmp21448;
  wire tmp21449;
  wire tmp21450;
  wire tmp21451;
  wire tmp21452;
  wire tmp21453;
  wire tmp21454;
  wire tmp21455;
  wire tmp21456;
  wire tmp21457;
  wire tmp21458;
  wire tmp21459;
  wire tmp21460;
  wire tmp21461;
  wire tmp21462;
  wire tmp21463;
  wire tmp21464;
  wire tmp21465;
  wire tmp21466;
  wire tmp21467;
  wire tmp21468;
  wire tmp21469;
  wire tmp21470;
  wire tmp21471;
  wire tmp21472;
  wire tmp21473;
  wire tmp21474;
  wire tmp21475;
  wire tmp21476;
  wire tmp21477;
  wire tmp21478;
  wire tmp21479;
  wire tmp21480;
  wire tmp21481;
  wire tmp21482;
  wire tmp21483;
  wire tmp21484;
  wire tmp21485;
  wire tmp21486;
  wire tmp21487;
  wire tmp21488;
  wire tmp21489;
  wire tmp21490;
  wire tmp21491;
  wire tmp21492;
  wire tmp21493;
  wire tmp21494;
  wire tmp21495;
  wire tmp21496;
  wire tmp21497;
  wire tmp21498;
  wire tmp21499;
  wire tmp21500;
  wire tmp21501;
  wire tmp21502;
  wire tmp21503;
  wire tmp21504;
  wire tmp21505;
  wire tmp21506;
  wire tmp21507;
  wire tmp21508;
  wire tmp21509;
  wire tmp21510;
  wire tmp21511;
  wire tmp21512;
  wire tmp21513;
  wire tmp21514;
  wire tmp21515;
  wire tmp21516;
  wire tmp21517;
  wire tmp21518;
  wire tmp21519;
  wire tmp21520;
  wire tmp21521;
  wire tmp21522;
  wire tmp21523;
  wire tmp21524;
  wire tmp21525;
  wire tmp21526;
  wire tmp21527;
  wire tmp21528;
  wire tmp21529;
  wire tmp21530;
  wire tmp21531;
  wire tmp21532;
  wire tmp21533;
  wire tmp21534;
  wire tmp21535;
  wire tmp21536;
  wire tmp21537;
  wire tmp21538;
  wire tmp21539;
  wire tmp21540;
  wire tmp21541;
  wire tmp21542;
  wire tmp21543;
  wire tmp21544;
  wire tmp21545;
  wire tmp21546;
  wire tmp21547;
  wire tmp21548;
  wire tmp21549;
  wire tmp21550;
  wire tmp21551;
  wire tmp21552;
  wire tmp21553;
  wire tmp21554;
  wire tmp21555;
  wire tmp21556;
  wire tmp21557;
  wire tmp21558;
  wire tmp21559;
  wire tmp21560;
  wire tmp21561;
  wire tmp21562;
  wire tmp21563;
  wire tmp21564;
  wire tmp21565;
  wire tmp21566;
  wire tmp21567;
  wire tmp21568;
  wire tmp21569;
  wire tmp21570;
  wire tmp21571;
  wire tmp21572;
  wire tmp21573;
  wire tmp21574;
  wire tmp21575;
  wire tmp21576;
  wire tmp21577;
  wire tmp21578;
  wire tmp21579;
  wire tmp21580;
  wire tmp21581;
  wire tmp21582;
  wire tmp21583;
  wire tmp21584;
  wire tmp21585;
  wire tmp21586;
  wire tmp21587;
  wire tmp21588;
  wire tmp21589;
  wire tmp21590;
  wire tmp21591;
  wire tmp21592;
  wire tmp21593;
  wire tmp21594;
  wire tmp21595;
  wire tmp21596;
  wire tmp21597;
  wire tmp21598;
  wire tmp21599;
  wire tmp21600;
  wire tmp21601;
  wire tmp21602;
  wire tmp21603;
  wire tmp21604;
  wire tmp21605;
  wire tmp21606;
  wire tmp21607;
  wire tmp21608;
  wire tmp21609;
  wire tmp21610;
  wire tmp21611;
  wire tmp21612;
  wire tmp21613;
  wire tmp21614;
  wire tmp21615;
  wire tmp21616;
  wire tmp21617;
  wire tmp21618;
  wire tmp21619;
  wire tmp21620;
  wire tmp21621;
  wire tmp21622;
  wire tmp21623;
  wire tmp21624;
  wire tmp21625;
  wire tmp21626;
  wire tmp21627;
  wire tmp21628;
  wire tmp21629;
  wire tmp21630;
  wire tmp21631;
  wire tmp21632;
  wire tmp21633;
  wire tmp21634;
  wire tmp21635;
  wire tmp21636;
  wire tmp21637;
  wire tmp21638;
  wire tmp21639;
  wire tmp21640;
  wire tmp21641;
  wire tmp21642;
  wire tmp21643;
  wire tmp21644;
  wire tmp21645;
  wire tmp21646;
  wire tmp21647;
  wire tmp21648;
  wire tmp21649;
  wire tmp21650;
  wire tmp21651;
  wire tmp21652;
  wire tmp21653;
  wire tmp21654;
  wire tmp21655;
  wire tmp21656;
  wire tmp21657;
  wire tmp21658;
  wire tmp21659;
  wire tmp21660;
  wire tmp21661;
  wire tmp21662;
  wire tmp21663;
  wire tmp21664;
  wire tmp21665;
  wire tmp21666;
  wire tmp21667;
  wire tmp21668;
  wire tmp21669;
  wire tmp21670;
  wire tmp21671;
  wire tmp21672;
  wire tmp21673;
  wire tmp21674;
  wire tmp21675;
  wire tmp21676;
  wire tmp21677;
  wire tmp21678;
  wire tmp21679;
  wire tmp21680;
  wire tmp21681;
  wire tmp21682;
  wire tmp21683;
  wire tmp21684;
  wire tmp21685;
  wire tmp21686;
  wire tmp21687;
  wire tmp21688;
  wire tmp21689;
  wire tmp21690;
  wire tmp21691;
  wire tmp21692;
  wire tmp21693;
  wire tmp21694;
  wire tmp21695;
  wire tmp21696;
  wire tmp21697;
  wire tmp21698;
  wire tmp21699;
  wire tmp21700;
  wire tmp21701;
  wire tmp21702;
  wire tmp21703;
  wire tmp21704;
  wire tmp21705;
  wire tmp21706;
  wire tmp21707;
  wire tmp21708;
  wire tmp21709;
  wire tmp21710;
  wire tmp21711;
  wire tmp21712;
  wire tmp21713;
  wire tmp21714;
  wire tmp21715;
  wire tmp21716;
  wire tmp21717;
  wire tmp21718;
  wire tmp21719;
  wire tmp21720;
  wire tmp21721;
  wire tmp21722;
  wire tmp21723;
  wire tmp21724;
  wire tmp21725;
  wire tmp21726;
  wire tmp21727;
  wire tmp21728;
  wire tmp21729;
  wire tmp21730;
  wire tmp21731;
  wire tmp21732;
  wire tmp21733;
  wire tmp21734;
  wire tmp21735;
  wire tmp21736;
  wire tmp21737;
  wire tmp21738;
  wire tmp21739;
  wire tmp21740;
  wire tmp21741;
  wire tmp21742;
  wire tmp21743;
  wire tmp21744;
  wire tmp21745;
  wire tmp21746;
  wire tmp21747;
  wire tmp21748;
  wire tmp21749;
  wire tmp21750;
  wire tmp21751;
  wire tmp21752;
  wire tmp21753;
  wire tmp21754;
  wire tmp21755;
  wire tmp21756;
  wire tmp21757;
  wire tmp21758;
  wire tmp21759;
  wire tmp21760;
  wire tmp21761;
  wire tmp21762;
  wire tmp21763;
  wire tmp21764;
  wire tmp21765;
  wire tmp21766;
  wire tmp21767;
  wire tmp21768;
  wire tmp21769;
  wire tmp21770;
  wire tmp21771;
  wire tmp21772;
  wire tmp21773;
  wire tmp21774;
  wire tmp21775;
  wire tmp21776;
  wire tmp21777;
  wire tmp21778;
  wire tmp21779;
  wire tmp21780;
  wire tmp21781;
  wire tmp21782;
  wire tmp21783;
  wire tmp21784;
  wire tmp21785;
  wire tmp21786;
  wire tmp21787;
  wire tmp21788;
  wire tmp21789;
  wire tmp21790;
  wire tmp21791;
  wire tmp21792;
  wire tmp21793;
  wire tmp21794;
  wire tmp21795;
  wire tmp21796;
  wire tmp21797;
  wire tmp21798;
  wire tmp21799;
  wire tmp21800;
  wire tmp21801;
  wire tmp21802;
  wire tmp21803;
  wire tmp21804;
  wire tmp21805;
  wire tmp21806;
  wire tmp21807;
  wire tmp21808;
  wire tmp21809;
  wire tmp21810;
  wire tmp21811;
  wire tmp21812;
  wire tmp21813;
  wire tmp21814;
  wire tmp21815;
  wire tmp21816;
  wire tmp21817;
  wire tmp21818;
  wire tmp21819;
  wire tmp21820;
  wire tmp21821;
  wire tmp21822;
  wire tmp21823;
  wire tmp21824;
  wire tmp21825;
  wire tmp21826;
  wire tmp21827;
  wire tmp21828;
  wire tmp21829;
  wire tmp21830;
  wire tmp21831;
  wire tmp21832;
  wire tmp21833;
  wire tmp21834;
  wire tmp21835;
  wire tmp21836;
  wire tmp21837;
  wire tmp21838;
  wire tmp21839;
  wire tmp21840;
  wire tmp21841;
  wire tmp21842;
  wire tmp21843;
  wire tmp21844;
  wire tmp21845;
  wire tmp21846;
  wire tmp21847;
  wire tmp21848;
  wire tmp21849;
  wire tmp21850;
  wire tmp21851;
  wire tmp21852;
  wire tmp21853;
  wire tmp21854;
  wire tmp21855;
  wire tmp21856;
  wire tmp21857;
  wire tmp21858;
  wire tmp21859;
  wire tmp21860;
  wire tmp21861;
  wire tmp21862;
  wire tmp21863;
  wire tmp21864;
  wire tmp21865;
  wire tmp21866;
  wire tmp21867;
  wire tmp21868;
  wire tmp21869;
  wire tmp21870;
  wire tmp21871;
  wire tmp21872;
  wire tmp21873;
  wire tmp21874;
  wire tmp21875;
  wire tmp21876;
  wire tmp21877;
  wire tmp21878;
  wire tmp21879;
  wire tmp21880;
  wire tmp21881;
  wire tmp21882;
  wire tmp21883;
  wire tmp21884;
  wire tmp21885;
  wire tmp21886;
  wire tmp21887;
  wire tmp21888;
  wire tmp21889;
  wire tmp21890;
  wire tmp21891;
  wire tmp21892;
  wire tmp21893;
  wire tmp21894;
  wire tmp21895;
  wire tmp21896;
  wire tmp21897;
  wire tmp21898;
  wire tmp21899;
  wire tmp21900;
  wire tmp21901;
  wire tmp21902;
  wire tmp21903;
  wire tmp21904;
  wire tmp21905;
  wire tmp21906;
  wire tmp21907;
  wire tmp21908;
  wire tmp21909;
  wire tmp21910;
  wire tmp21911;
  wire tmp21912;
  wire tmp21913;
  wire tmp21914;
  wire tmp21915;
  wire tmp21916;
  wire tmp21917;
  wire tmp21918;
  wire tmp21919;
  wire tmp21920;
  wire tmp21921;
  wire tmp21922;
  wire tmp21923;
  wire tmp21924;
  wire tmp21925;
  wire tmp21926;
  wire tmp21927;
  wire tmp21928;
  wire tmp21929;
  wire tmp21930;
  wire tmp21931;
  wire tmp21932;
  wire tmp21933;
  wire tmp21934;
  wire tmp21935;
  wire tmp21936;
  wire tmp21937;
  wire tmp21938;
  wire tmp21939;
  wire tmp21940;
  wire tmp21941;
  wire tmp21942;
  wire tmp21943;
  wire tmp21944;
  wire tmp21945;
  wire tmp21946;
  wire tmp21947;
  wire tmp21948;
  wire tmp21949;
  wire tmp21950;
  wire tmp21951;
  wire tmp21952;
  wire tmp21953;
  wire tmp21954;
  wire tmp21955;
  wire tmp21956;
  wire tmp21957;
  wire tmp21958;
  wire tmp21959;
  wire tmp21960;
  wire tmp21961;
  wire tmp21962;
  wire tmp21963;
  wire tmp21964;
  wire tmp21965;
  wire tmp21966;
  wire tmp21967;
  wire tmp21968;
  wire tmp21969;
  wire tmp21970;
  wire tmp21971;
  wire tmp21972;
  wire tmp21973;
  wire tmp21974;
  wire tmp21975;
  wire tmp21976;
  wire tmp21977;
  wire tmp21978;
  wire tmp21979;
  wire tmp21980;
  wire tmp21981;
  wire tmp21982;
  wire tmp21983;
  wire tmp21984;
  wire tmp21985;
  wire tmp21986;
  wire tmp21987;
  wire tmp21988;
  wire tmp21989;
  wire tmp21990;
  wire tmp21991;
  wire tmp21992;
  wire tmp21993;
  wire tmp21994;
  wire tmp21995;
  wire tmp21996;
  wire tmp21997;
  wire tmp21998;
  wire tmp21999;
  wire tmp22000;
  wire tmp22001;
  wire tmp22002;
  wire tmp22003;
  wire tmp22004;
  wire tmp22005;
  wire tmp22006;
  wire tmp22007;
  wire tmp22008;
  wire tmp22009;
  wire tmp22010;
  wire tmp22011;
  wire tmp22012;
  wire tmp22013;
  wire tmp22014;
  wire tmp22015;
  wire tmp22016;
  wire tmp22017;
  wire tmp22018;
  wire tmp22019;
  wire tmp22020;
  wire tmp22021;
  wire tmp22022;
  wire tmp22023;
  wire tmp22024;
  wire tmp22025;
  wire tmp22026;
  wire tmp22027;
  wire tmp22028;
  wire tmp22029;
  wire tmp22030;
  wire tmp22031;
  wire tmp22032;
  wire tmp22033;
  wire tmp22034;
  wire tmp22035;
  wire tmp22036;
  wire tmp22037;
  wire tmp22038;
  wire tmp22039;
  wire tmp22040;
  wire tmp22041;
  wire tmp22042;
  wire tmp22043;
  wire tmp22044;
  wire tmp22045;
  wire tmp22046;
  wire tmp22047;
  wire tmp22048;
  wire tmp22049;
  wire tmp22050;
  wire tmp22051;
  wire tmp22052;
  wire tmp22053;
  wire tmp22054;
  wire tmp22055;
  wire tmp22056;
  wire tmp22057;
  wire tmp22058;
  wire tmp22059;
  wire tmp22060;
  wire tmp22061;
  wire tmp22062;
  wire tmp22063;
  wire tmp22064;
  wire tmp22065;
  wire tmp22066;
  wire tmp22067;
  wire tmp22068;
  wire tmp22069;
  wire tmp22070;
  wire tmp22071;
  wire tmp22072;
  wire tmp22073;
  wire tmp22074;
  wire tmp22075;
  wire tmp22076;
  wire tmp22077;
  wire tmp22078;
  wire tmp22079;
  wire tmp22080;
  wire tmp22081;
  wire tmp22082;
  wire tmp22083;
  wire tmp22084;
  wire tmp22085;
  wire tmp22086;
  wire tmp22087;
  wire tmp22088;
  wire tmp22089;
  wire tmp22090;
  wire tmp22091;
  wire tmp22092;
  wire tmp22093;
  wire tmp22094;
  wire tmp22095;
  wire tmp22096;
  wire tmp22097;
  wire tmp22098;
  wire tmp22099;
  wire tmp22100;
  wire tmp22101;
  wire tmp22102;
  wire tmp22103;
  wire tmp22104;
  wire tmp22105;
  wire tmp22106;
  wire tmp22107;
  wire tmp22108;
  wire tmp22109;
  wire tmp22110;
  wire tmp22111;
  wire tmp22112;
  wire tmp22113;
  wire tmp22114;
  wire tmp22115;
  wire tmp22116;
  wire tmp22117;
  wire tmp22118;
  wire tmp22119;
  wire tmp22120;
  wire tmp22121;
  wire tmp22122;
  wire tmp22123;
  wire tmp22124;
  wire tmp22125;
  wire tmp22126;
  wire tmp22127;
  wire tmp22128;
  wire tmp22129;
  wire tmp22130;
  wire tmp22131;
  wire tmp22132;
  wire tmp22133;
  wire tmp22134;
  wire tmp22135;
  wire tmp22136;
  wire tmp22137;
  wire tmp22138;
  wire tmp22139;
  wire tmp22140;
  wire tmp22141;
  wire tmp22142;
  wire tmp22143;
  wire tmp22144;
  wire tmp22145;
  wire tmp22146;
  wire tmp22147;
  wire tmp22148;
  wire tmp22149;
  wire tmp22150;
  wire tmp22151;
  wire tmp22152;
  wire tmp22153;
  wire tmp22154;
  wire tmp22155;
  wire tmp22156;
  wire tmp22157;
  wire tmp22158;
  wire tmp22159;
  wire tmp22160;
  wire tmp22161;
  wire tmp22162;
  wire tmp22163;
  wire tmp22164;
  wire tmp22165;
  wire tmp22166;
  wire tmp22167;
  wire tmp22168;
  wire tmp22169;
  wire tmp22170;
  wire tmp22171;
  wire tmp22172;
  wire tmp22173;
  wire tmp22174;
  wire tmp22175;
  wire tmp22176;
  wire tmp22177;
  wire tmp22178;
  wire tmp22179;
  wire tmp22180;
  wire tmp22181;
  wire tmp22182;
  wire tmp22183;
  wire tmp22184;
  wire tmp22185;
  wire tmp22186;
  wire tmp22187;
  wire tmp22188;
  wire tmp22189;
  wire tmp22190;
  wire tmp22191;
  wire tmp22192;
  wire tmp22193;
  wire tmp22194;
  wire tmp22195;
  wire tmp22196;
  wire tmp22197;
  wire tmp22198;
  wire tmp22199;
  wire tmp22200;
  wire tmp22201;
  wire tmp22202;
  wire tmp22203;
  wire tmp22204;
  wire tmp22205;
  wire tmp22206;
  wire tmp22207;
  wire tmp22208;
  wire tmp22209;
  wire tmp22210;
  wire tmp22211;
  wire tmp22212;
  wire tmp22213;
  wire tmp22214;
  wire tmp22215;
  wire tmp22216;
  wire tmp22217;
  wire tmp22218;
  wire tmp22219;
  wire tmp22220;
  wire tmp22221;
  wire tmp22222;
  wire tmp22223;
  wire tmp22224;
  wire tmp22225;
  wire tmp22226;
  wire tmp22227;
  wire tmp22228;
  wire tmp22229;
  wire tmp22230;
  wire tmp22231;
  wire tmp22232;
  wire tmp22233;
  wire tmp22234;
  wire tmp22235;
  wire tmp22236;
  wire tmp22237;
  wire tmp22238;
  wire tmp22239;
  wire tmp22240;
  wire tmp22241;
  wire tmp22242;
  wire tmp22243;
  wire tmp22244;
  wire tmp22245;
  wire tmp22246;
  wire tmp22247;
  wire tmp22248;
  wire tmp22249;
  wire tmp22250;
  wire tmp22251;
  wire tmp22252;
  wire tmp22253;
  wire tmp22254;
  wire tmp22255;
  wire tmp22256;
  wire tmp22257;
  wire tmp22258;
  wire tmp22259;
  wire tmp22260;
  wire tmp22261;
  wire tmp22262;
  wire tmp22263;
  wire tmp22264;
  wire tmp22265;
  wire tmp22266;
  wire tmp22267;
  wire tmp22268;
  wire tmp22269;
  wire tmp22270;
  wire tmp22271;
  wire tmp22272;
  wire tmp22273;
  wire tmp22274;
  wire tmp22275;
  wire tmp22276;
  wire tmp22277;
  wire tmp22278;
  wire tmp22279;
  wire tmp22280;
  wire tmp22281;
  wire tmp22282;
  wire tmp22283;
  wire tmp22284;
  wire tmp22285;
  wire tmp22286;
  wire tmp22287;
  wire tmp22288;
  wire tmp22289;
  wire tmp22290;
  wire tmp22291;
  wire tmp22292;
  wire tmp22293;
  wire tmp22294;
  wire tmp22295;
  wire tmp22296;
  wire tmp22297;
  wire tmp22298;
  wire tmp22299;
  wire tmp22300;
  wire tmp22301;
  wire tmp22302;
  wire tmp22303;
  wire tmp22304;
  wire tmp22305;
  wire tmp22306;
  wire tmp22307;
  wire tmp22308;
  wire tmp22309;
  wire tmp22310;
  wire tmp22311;
  wire tmp22312;
  wire tmp22313;
  wire tmp22314;
  wire tmp22315;
  wire tmp22316;
  wire tmp22317;
  wire tmp22318;
  wire tmp22319;
  wire tmp22320;
  wire tmp22321;
  wire tmp22322;
  wire tmp22323;
  wire tmp22324;
  wire tmp22325;
  wire tmp22326;
  wire tmp22327;
  wire tmp22328;
  wire tmp22329;
  wire tmp22330;
  wire tmp22331;
  wire tmp22332;
  wire tmp22333;
  wire tmp22334;
  wire tmp22335;
  wire tmp22336;
  wire tmp22337;
  wire tmp22338;
  wire tmp22339;
  wire tmp22340;
  wire tmp22341;
  wire tmp22342;
  wire tmp22343;
  wire tmp22344;
  wire tmp22345;
  wire tmp22346;
  wire tmp22347;
  wire tmp22348;
  wire tmp22349;
  wire tmp22350;
  wire tmp22351;
  wire tmp22352;
  wire tmp22353;
  wire tmp22354;
  wire tmp22355;
  wire tmp22356;
  wire tmp22357;
  wire tmp22358;
  wire tmp22359;
  wire tmp22360;
  wire tmp22361;
  wire tmp22362;
  wire tmp22363;
  wire tmp22364;
  wire tmp22365;
  wire tmp22366;
  wire tmp22367;
  wire tmp22368;
  wire tmp22369;
  wire tmp22370;
  wire tmp22371;
  wire tmp22372;
  wire tmp22373;
  wire tmp22374;
  wire tmp22375;
  wire tmp22376;
  wire tmp22377;
  wire tmp22378;
  wire tmp22379;
  wire tmp22380;
  wire tmp22381;
  wire tmp22382;
  wire tmp22383;
  wire tmp22384;
  wire tmp22385;
  wire tmp22386;
  wire tmp22387;
  wire tmp22388;
  wire tmp22389;
  wire tmp22390;
  wire tmp22391;
  wire tmp22392;
  wire tmp22393;
  wire tmp22394;
  wire tmp22395;
  wire tmp22396;
  wire tmp22397;
  wire tmp22398;
  wire tmp22399;
  wire tmp22400;
  wire tmp22401;
  wire tmp22402;
  wire tmp22403;
  wire tmp22404;
  wire tmp22405;
  wire tmp22406;
  wire tmp22407;
  wire tmp22408;
  wire tmp22409;
  wire tmp22410;
  wire tmp22411;
  wire tmp22412;
  wire tmp22413;
  wire tmp22414;
  wire tmp22415;
  wire tmp22416;
  wire tmp22417;
  wire tmp22418;
  wire tmp22419;
  wire tmp22420;
  wire tmp22421;
  wire tmp22422;
  wire tmp22423;
  wire tmp22424;
  wire tmp22425;
  wire tmp22426;
  wire tmp22427;
  wire tmp22428;
  wire tmp22429;
  wire tmp22430;
  wire tmp22431;
  wire tmp22432;
  wire tmp22433;
  wire tmp22434;
  wire tmp22435;
  wire tmp22436;
  wire tmp22437;
  wire tmp22438;
  wire tmp22439;
  wire tmp22440;
  wire tmp22441;
  wire tmp22442;
  wire tmp22443;
  wire tmp22444;
  wire tmp22445;
  wire tmp22446;
  wire tmp22447;
  wire tmp22448;
  wire tmp22449;
  wire tmp22450;
  wire tmp22451;
  wire tmp22452;
  wire tmp22453;
  wire tmp22454;
  wire tmp22455;
  wire tmp22456;
  wire tmp22457;
  wire tmp22458;
  wire tmp22459;
  wire tmp22460;
  wire tmp22461;
  wire tmp22462;
  wire tmp22463;
  wire tmp22464;
  wire tmp22465;
  wire tmp22466;
  wire tmp22467;
  wire tmp22468;
  wire tmp22469;
  wire tmp22470;
  wire tmp22471;
  wire tmp22472;
  wire tmp22473;
  wire tmp22474;
  wire tmp22475;
  wire tmp22476;
  wire tmp22477;
  wire tmp22478;
  wire tmp22479;
  wire tmp22480;
  wire tmp22481;
  wire tmp22482;
  wire tmp22483;
  wire tmp22484;
  wire tmp22485;
  wire tmp22486;
  wire tmp22487;
  wire tmp22488;
  wire tmp22489;
  wire tmp22490;
  wire tmp22491;
  wire tmp22492;
  wire tmp22493;
  wire tmp22494;
  wire tmp22495;
  wire tmp22496;
  wire tmp22497;
  wire tmp22498;
  wire tmp22499;
  wire tmp22500;
  wire tmp22501;
  wire tmp22502;
  wire tmp22503;
  wire tmp22504;
  wire tmp22505;
  wire tmp22506;
  wire tmp22507;
  wire tmp22508;
  wire tmp22509;
  wire tmp22510;
  wire tmp22511;
  wire tmp22512;
  wire tmp22513;
  wire tmp22514;
  wire tmp22515;
  wire tmp22516;
  wire tmp22517;
  wire tmp22518;
  wire tmp22519;
  wire tmp22520;
  wire tmp22521;
  wire tmp22522;
  wire tmp22523;
  wire tmp22524;
  wire tmp22525;
  wire tmp22526;
  wire tmp22527;
  wire tmp22528;
  wire tmp22529;
  wire tmp22530;
  wire tmp22531;
  wire tmp22532;
  wire tmp22533;
  wire tmp22534;
  wire tmp22535;
  wire tmp22536;
  wire tmp22537;
  wire tmp22538;
  wire tmp22539;
  wire tmp22540;
  wire tmp22541;
  wire tmp22542;
  wire tmp22543;
  wire tmp22544;
  wire tmp22545;
  wire tmp22546;
  wire tmp22547;
  wire tmp22548;
  wire tmp22549;
  wire tmp22550;
  wire tmp22551;
  wire tmp22552;
  wire tmp22553;
  wire tmp22554;
  wire tmp22555;
  wire tmp22556;
  wire tmp22557;
  wire tmp22558;
  wire tmp22559;
  wire tmp22560;
  wire tmp22561;
  wire tmp22562;
  wire tmp22563;
  wire tmp22564;
  wire tmp22565;
  wire tmp22566;
  wire tmp22567;
  wire tmp22568;
  wire tmp22569;
  wire tmp22570;
  wire tmp22571;
  wire tmp22572;
  wire tmp22573;
  wire tmp22574;
  wire tmp22575;
  wire tmp22576;
  wire tmp22577;
  wire tmp22578;
  wire tmp22579;
  wire tmp22580;
  wire tmp22581;
  wire tmp22582;
  wire tmp22583;
  wire tmp22584;
  wire tmp22585;
  wire tmp22586;
  wire tmp22587;
  wire tmp22588;
  wire tmp22589;
  wire tmp22590;
  wire tmp22591;
  wire tmp22592;
  wire tmp22593;
  wire tmp22594;
  wire tmp22595;
  wire tmp22596;
  wire tmp22597;
  wire tmp22598;
  wire tmp22599;
  wire tmp22600;
  wire tmp22601;
  wire tmp22602;
  wire tmp22603;
  wire tmp22604;
  wire tmp22605;
  wire tmp22606;
  wire tmp22607;
  wire tmp22608;
  wire tmp22609;
  wire tmp22610;
  wire tmp22611;
  wire tmp22612;
  wire tmp22613;
  wire tmp22614;
  wire tmp22615;
  wire tmp22616;
  wire tmp22617;
  wire tmp22618;
  wire tmp22619;
  wire tmp22620;
  wire tmp22621;
  wire tmp22622;
  wire tmp22623;
  wire tmp22624;
  wire tmp22625;
  wire tmp22626;
  wire tmp22627;
  wire tmp22628;
  wire tmp22629;
  wire tmp22630;
  wire tmp22631;
  wire tmp22632;
  wire tmp22633;
  wire tmp22634;
  wire tmp22635;
  wire tmp22636;
  wire tmp22637;
  wire tmp22638;
  wire tmp22639;
  wire tmp22640;
  wire tmp22641;
  wire tmp22642;
  wire tmp22643;
  wire tmp22644;
  wire tmp22645;
  wire tmp22646;
  wire tmp22647;
  wire tmp22648;
  wire tmp22649;
  wire tmp22650;
  wire tmp22651;
  wire tmp22652;
  wire tmp22653;
  wire tmp22654;
  wire tmp22655;
  wire tmp22656;
  wire tmp22657;
  wire tmp22658;
  wire tmp22659;
  wire tmp22660;
  wire tmp22661;
  wire tmp22662;
  wire tmp22663;
  wire tmp22664;
  wire tmp22665;
  wire tmp22666;
  wire tmp22667;
  wire tmp22668;
  wire tmp22669;
  wire tmp22670;
  wire tmp22671;
  wire tmp22672;
  wire tmp22673;
  wire tmp22674;
  wire tmp22675;
  wire tmp22676;
  wire tmp22677;
  wire tmp22678;
  wire tmp22679;
  wire tmp22680;
  wire tmp22681;
  wire tmp22682;
  wire tmp22683;
  wire tmp22684;
  wire tmp22685;
  wire tmp22686;
  wire tmp22687;
  wire tmp22688;
  wire tmp22689;
  wire tmp22690;
  wire tmp22691;
  wire tmp22692;
  wire tmp22693;
  wire tmp22694;
  wire tmp22695;
  wire tmp22696;
  wire tmp22697;
  wire tmp22698;
  wire tmp22699;
  wire tmp22700;
  wire tmp22701;
  wire tmp22702;
  wire tmp22703;
  wire tmp22704;
  wire tmp22705;
  wire tmp22706;
  wire tmp22707;
  wire tmp22708;
  wire tmp22709;
  wire tmp22710;
  wire tmp22711;
  wire tmp22712;
  wire tmp22713;
  wire tmp22714;
  wire tmp22715;
  wire tmp22716;
  wire tmp22717;
  wire tmp22718;
  wire tmp22719;
  wire tmp22720;
  wire tmp22721;
  wire tmp22722;
  wire tmp22723;
  wire tmp22724;
  wire tmp22725;
  wire tmp22726;
  wire tmp22727;
  wire tmp22728;
  wire tmp22729;
  wire tmp22730;
  wire tmp22731;
  wire tmp22732;
  wire tmp22733;
  wire tmp22734;
  wire tmp22735;
  wire tmp22736;
  wire tmp22737;
  wire tmp22738;
  wire tmp22739;
  wire tmp22740;
  wire tmp22741;
  wire tmp22742;
  wire tmp22743;
  wire tmp22744;
  wire tmp22745;
  wire tmp22746;
  wire tmp22747;
  wire tmp22748;
  wire tmp22749;
  wire tmp22750;
  wire tmp22751;
  wire tmp22752;
  wire tmp22753;
  wire tmp22754;
  wire tmp22755;
  wire tmp22756;
  wire tmp22757;
  wire tmp22758;
  wire tmp22759;
  wire tmp22760;
  wire tmp22761;
  wire tmp22762;
  wire tmp22763;
  wire tmp22764;
  wire tmp22765;
  wire tmp22766;
  wire tmp22767;
  wire tmp22768;
  wire tmp22769;
  wire tmp22770;
  wire tmp22771;
  wire tmp22772;
  wire tmp22773;
  wire tmp22774;
  wire tmp22775;
  wire tmp22776;
  wire tmp22777;
  wire tmp22778;
  wire tmp22779;
  wire tmp22780;
  wire tmp22781;
  wire tmp22782;
  wire tmp22783;
  wire tmp22784;
  wire tmp22785;
  wire tmp22786;
  wire tmp22787;
  wire tmp22788;
  wire tmp22789;
  wire tmp22790;
  wire tmp22791;
  wire tmp22792;
  wire tmp22793;
  wire tmp22794;
  wire tmp22795;
  wire tmp22796;
  wire tmp22797;
  wire tmp22798;
  wire tmp22799;
  wire tmp22800;
  wire tmp22801;
  wire tmp22802;
  wire tmp22803;
  wire tmp22804;
  wire tmp22805;
  wire tmp22806;
  wire tmp22807;
  wire tmp22808;
  wire tmp22809;
  wire tmp22810;
  wire tmp22811;
  wire tmp22812;
  wire tmp22813;
  wire tmp22814;
  wire tmp22815;
  wire tmp22816;
  wire tmp22817;
  wire tmp22818;
  wire tmp22819;
  wire tmp22820;
  wire tmp22821;
  wire tmp22822;
  wire tmp22823;
  wire tmp22824;
  wire tmp22825;
  wire tmp22826;
  wire tmp22827;
  wire tmp22828;
  wire tmp22829;
  wire tmp22830;
  wire tmp22831;
  wire tmp22832;
  wire tmp22833;
  wire tmp22834;
  wire tmp22835;
  wire tmp22836;
  wire tmp22837;
  wire tmp22838;
  wire tmp22839;
  wire tmp22840;
  wire tmp22841;
  wire tmp22842;
  wire tmp22843;
  wire tmp22844;
  wire tmp22845;
  wire tmp22846;
  wire tmp22847;
  wire tmp22848;
  wire tmp22849;
  wire tmp22850;
  wire tmp22851;
  wire tmp22852;
  wire tmp22853;
  wire tmp22854;
  wire tmp22855;
  wire tmp22856;
  wire tmp22857;
  wire tmp22858;
  wire tmp22859;
  wire tmp22860;
  wire tmp22861;
  wire tmp22862;
  wire tmp22863;
  wire tmp22864;
  wire tmp22865;
  wire tmp22866;
  wire tmp22867;
  wire tmp22868;
  wire tmp22869;
  wire tmp22870;
  wire tmp22871;
  wire tmp22872;
  wire tmp22873;
  wire tmp22874;
  wire tmp22875;
  wire tmp22876;
  wire tmp22877;
  wire tmp22878;
  wire tmp22879;
  wire tmp22880;
  wire tmp22881;
  wire tmp22882;
  wire tmp22883;
  wire tmp22884;
  wire tmp22885;
  wire tmp22886;
  wire tmp22887;
  wire tmp22888;
  wire tmp22889;
  wire tmp22890;
  wire tmp22891;
  wire tmp22892;
  wire tmp22893;
  wire tmp22894;
  wire tmp22895;
  wire tmp22896;
  wire tmp22897;
  wire tmp22898;
  wire tmp22899;
  wire tmp22900;
  wire tmp22901;
  wire tmp22902;
  wire tmp22903;
  wire tmp22904;
  wire tmp22905;
  wire tmp22906;
  wire tmp22907;
  wire tmp22908;
  wire tmp22909;
  wire tmp22910;
  wire tmp22911;
  wire tmp22912;
  wire tmp22913;
  wire tmp22914;
  wire tmp22915;
  wire tmp22916;
  wire tmp22917;
  wire tmp22918;
  wire tmp22919;
  wire tmp22920;
  wire tmp22921;
  wire tmp22922;
  wire tmp22923;
  wire tmp22924;
  wire tmp22925;
  wire tmp22926;
  wire tmp22927;
  wire tmp22928;
  wire tmp22929;
  wire tmp22930;
  wire tmp22931;
  wire tmp22932;
  wire tmp22933;
  wire tmp22934;
  wire tmp22935;
  wire tmp22936;
  wire tmp22937;
  wire tmp22938;
  wire tmp22939;
  wire tmp22940;
  wire tmp22941;
  wire tmp22942;
  wire tmp22943;
  wire tmp22944;
  wire tmp22945;
  wire tmp22946;
  wire tmp22947;
  wire tmp22948;
  wire tmp22949;
  wire tmp22950;
  wire tmp22951;
  wire tmp22952;
  wire tmp22953;
  wire tmp22954;
  wire tmp22955;
  wire tmp22956;
  wire tmp22957;
  wire tmp22958;
  wire tmp22959;
  wire tmp22960;
  wire tmp22961;
  wire tmp22962;
  wire tmp22963;
  wire tmp22964;
  wire tmp22965;
  wire tmp22966;
  wire tmp22967;
  wire tmp22968;
  wire tmp22969;
  wire tmp22970;
  wire tmp22971;
  wire tmp22972;
  wire tmp22973;
  wire tmp22974;
  wire tmp22975;
  wire tmp22976;
  wire tmp22977;
  wire tmp22978;
  wire tmp22979;
  wire tmp22980;
  wire tmp22981;
  wire tmp22982;
  wire tmp22983;
  wire tmp22984;
  wire tmp22985;
  wire tmp22986;
  wire tmp22987;
  wire tmp22988;
  wire tmp22989;
  wire tmp22990;
  wire tmp22991;
  wire tmp22992;
  wire tmp22993;
  wire tmp22994;
  wire tmp22995;
  wire tmp22996;
  wire tmp22997;
  wire tmp22998;
  wire tmp22999;
  wire tmp23000;
  wire tmp23001;
  wire tmp23002;
  wire tmp23003;
  wire tmp23004;
  wire tmp23005;
  wire tmp23006;
  wire tmp23007;
  wire tmp23008;
  wire tmp23009;
  wire tmp23010;
  wire tmp23011;
  wire tmp23012;
  wire tmp23013;
  wire tmp23014;
  wire tmp23015;
  wire tmp23016;
  wire tmp23017;
  wire tmp23018;
  wire tmp23019;
  wire tmp23020;
  wire tmp23021;
  wire tmp23022;
  wire tmp23023;
  wire tmp23024;
  wire tmp23025;
  wire tmp23026;
  wire tmp23027;
  wire tmp23028;
  wire tmp23029;
  wire tmp23030;
  wire tmp23031;
  wire tmp23032;
  wire tmp23033;
  wire tmp23034;
  wire tmp23035;
  wire tmp23036;
  wire tmp23037;
  wire tmp23038;
  wire tmp23039;
  wire tmp23040;
  wire tmp23041;
  wire tmp23042;
  wire tmp23043;
  wire tmp23044;
  wire tmp23045;
  wire tmp23046;
  wire tmp23047;
  wire tmp23048;
  wire tmp23049;
  wire tmp23050;
  wire tmp23051;
  wire tmp23052;
  wire tmp23053;
  wire tmp23054;
  wire tmp23055;
  wire tmp23056;
  wire tmp23057;
  wire tmp23058;
  wire tmp23059;
  wire tmp23060;
  wire tmp23061;
  wire tmp23062;
  wire tmp23063;
  wire tmp23064;
  wire tmp23065;
  wire tmp23066;
  wire tmp23067;
  wire tmp23068;
  wire tmp23069;
  wire tmp23070;
  wire tmp23071;
  wire tmp23072;
  wire tmp23073;
  wire tmp23074;
  wire tmp23075;
  wire tmp23076;
  wire tmp23077;
  wire tmp23078;
  wire tmp23079;
  wire tmp23080;
  wire tmp23081;
  wire tmp23082;
  wire tmp23083;
  wire tmp23084;
  wire tmp23085;
  wire tmp23086;
  wire tmp23087;
  wire tmp23088;
  wire tmp23089;
  wire tmp23090;
  wire tmp23091;
  wire tmp23092;
  wire tmp23093;
  wire tmp23094;
  wire tmp23095;
  wire tmp23096;
  wire tmp23097;
  wire tmp23098;
  wire tmp23099;
  wire tmp23100;
  wire tmp23101;
  wire tmp23102;
  wire tmp23103;
  wire tmp23104;
  wire tmp23105;
  wire tmp23106;
  wire tmp23107;
  wire tmp23108;
  wire tmp23109;
  wire tmp23110;
  wire tmp23111;
  wire tmp23112;
  wire tmp23113;
  wire tmp23114;
  wire tmp23115;
  wire tmp23116;
  wire tmp23117;
  wire tmp23118;
  wire tmp23119;
  wire tmp23120;
  wire tmp23121;
  wire tmp23122;
  wire tmp23123;
  wire tmp23124;
  wire tmp23125;
  wire tmp23126;
  wire tmp23127;
  wire tmp23128;
  wire tmp23129;
  wire tmp23130;
  wire tmp23131;
  wire tmp23132;
  wire tmp23133;
  wire tmp23134;
  wire tmp23135;
  wire tmp23136;
  wire tmp23137;
  wire tmp23138;
  wire tmp23139;
  wire tmp23140;
  wire tmp23141;
  wire tmp23142;
  wire tmp23143;
  wire tmp23144;
  wire tmp23145;
  wire tmp23146;
  wire tmp23147;
  wire tmp23148;
  wire tmp23149;
  wire tmp23150;
  wire tmp23151;
  wire tmp23152;
  wire tmp23153;
  wire tmp23154;
  wire tmp23155;
  wire tmp23156;
  wire tmp23157;
  wire tmp23158;
  wire tmp23159;
  wire tmp23160;
  wire tmp23161;
  wire tmp23162;
  wire tmp23163;
  wire tmp23164;
  wire tmp23165;
  wire tmp23166;
  wire tmp23167;
  wire tmp23168;
  wire tmp23169;
  wire tmp23170;
  wire tmp23171;
  wire tmp23172;
  wire tmp23173;
  wire tmp23174;
  wire tmp23175;
  wire tmp23176;
  wire tmp23177;
  wire tmp23178;
  wire tmp23179;
  wire tmp23180;
  wire tmp23181;
  wire tmp23182;
  wire tmp23183;
  wire tmp23184;
  wire tmp23185;
  wire tmp23186;
  wire tmp23187;
  wire tmp23188;
  wire tmp23189;
  wire tmp23190;
  wire tmp23191;
  wire tmp23192;
  wire tmp23193;
  wire tmp23194;
  wire tmp23195;
  wire tmp23196;
  wire tmp23197;
  wire tmp23198;
  wire tmp23199;
  wire tmp23200;
  wire tmp23201;
  wire tmp23202;
  wire tmp23203;
  wire tmp23204;
  wire tmp23205;
  wire tmp23206;
  wire tmp23207;
  wire tmp23208;
  wire tmp23209;
  wire tmp23210;
  wire tmp23211;
  wire tmp23212;
  wire tmp23213;
  wire tmp23214;
  wire tmp23215;
  wire tmp23216;
  wire tmp23217;
  wire tmp23218;
  wire tmp23219;
  wire tmp23220;
  wire tmp23221;
  wire tmp23222;
  wire tmp23223;
  wire tmp23224;
  wire tmp23225;
  wire tmp23226;
  wire tmp23227;
  wire tmp23228;
  wire tmp23229;
  wire tmp23230;
  wire tmp23231;
  wire tmp23232;
  wire tmp23233;
  wire tmp23234;
  wire tmp23235;
  wire tmp23236;
  wire tmp23237;
  wire tmp23238;
  wire tmp23239;
  wire tmp23240;
  wire tmp23241;
  wire tmp23242;
  wire tmp23243;
  wire tmp23244;
  wire tmp23245;
  wire tmp23246;
  wire tmp23247;
  wire tmp23248;
  wire tmp23249;
  wire tmp23250;
  wire tmp23251;
  wire tmp23252;
  wire tmp23253;
  wire tmp23254;
  wire tmp23255;
  wire tmp23256;
  wire tmp23257;
  wire tmp23258;
  wire tmp23259;
  wire tmp23260;
  wire tmp23261;
  wire tmp23262;
  wire tmp23263;
  wire tmp23264;
  wire tmp23265;
  wire tmp23266;
  wire tmp23267;
  wire tmp23268;
  wire tmp23269;
  wire tmp23270;
  wire tmp23271;
  wire tmp23272;
  wire tmp23273;
  wire tmp23274;
  wire tmp23275;
  wire tmp23276;
  wire tmp23277;
  wire tmp23278;
  wire tmp23279;
  wire tmp23280;
  wire tmp23281;
  wire tmp23282;
  wire tmp23283;
  wire tmp23284;
  wire tmp23285;
  wire tmp23286;
  wire tmp23287;
  wire tmp23288;
  wire tmp23289;
  wire tmp23290;
  wire tmp23291;
  wire tmp23292;
  wire tmp23293;
  wire tmp23294;
  wire tmp23295;
  wire tmp23296;
  wire tmp23297;
  wire tmp23298;
  wire tmp23299;
  wire tmp23300;
  wire tmp23301;
  wire tmp23302;
  wire tmp23303;
  wire tmp23304;
  wire tmp23305;
  wire tmp23306;
  wire tmp23307;
  wire tmp23308;
  wire tmp23309;
  wire tmp23310;
  wire tmp23311;
  wire tmp23312;
  wire tmp23313;
  wire tmp23314;
  wire tmp23315;
  wire tmp23316;
  wire tmp23317;
  wire tmp23318;
  wire tmp23319;
  wire tmp23320;
  wire tmp23321;
  wire tmp23322;
  wire tmp23323;
  wire tmp23324;
  wire tmp23325;
  wire tmp23326;
  wire tmp23327;
  wire tmp23328;
  wire tmp23329;
  wire tmp23330;
  wire tmp23331;
  wire tmp23332;
  wire tmp23333;
  wire tmp23334;
  wire tmp23335;
  wire tmp23336;
  wire tmp23337;
  wire tmp23338;
  wire tmp23339;
  wire tmp23340;
  wire tmp23341;
  wire tmp23342;
  wire tmp23343;
  wire tmp23344;
  wire tmp23345;
  wire tmp23346;
  wire tmp23347;
  wire tmp23348;
  wire tmp23349;
  wire tmp23350;
  wire tmp23351;
  wire tmp23352;
  wire tmp23353;
  wire tmp23354;
  wire tmp23355;
  wire tmp23356;
  wire tmp23357;
  wire tmp23358;
  wire tmp23359;
  wire tmp23360;
  wire tmp23361;
  wire tmp23362;
  wire tmp23363;
  wire tmp23364;
  wire tmp23365;
  wire tmp23366;
  wire tmp23367;
  wire tmp23368;
  wire tmp23369;
  wire tmp23370;
  wire tmp23371;
  wire tmp23372;
  wire tmp23373;
  wire tmp23374;
  wire tmp23375;
  wire tmp23376;
  wire tmp23377;
  wire tmp23378;
  wire tmp23379;
  wire tmp23380;
  wire tmp23381;
  wire tmp23382;
  wire tmp23383;
  wire tmp23384;
  wire tmp23385;
  wire tmp23386;
  wire tmp23387;
  wire tmp23388;
  wire tmp23389;
  wire tmp23390;
  wire tmp23391;
  wire tmp23392;
  wire tmp23393;
  wire tmp23394;
  wire tmp23395;
  wire tmp23396;
  wire tmp23397;
  wire tmp23398;
  wire tmp23399;
  wire tmp23400;
  wire tmp23401;
  wire tmp23402;
  wire tmp23403;
  wire tmp23404;
  wire tmp23405;
  wire tmp23406;
  wire tmp23407;
  wire tmp23408;
  wire tmp23409;
  wire tmp23410;
  wire tmp23411;
  wire tmp23412;
  wire tmp23413;
  wire tmp23414;
  wire tmp23415;
  wire tmp23416;
  wire tmp23417;
  wire tmp23418;
  wire tmp23419;
  wire tmp23420;
  wire tmp23421;
  wire tmp23422;
  wire tmp23423;
  wire tmp23424;
  wire tmp23425;
  wire tmp23426;
  wire tmp23427;
  wire tmp23428;
  wire tmp23429;
  wire tmp23430;
  wire tmp23431;
  wire tmp23432;
  wire tmp23433;
  wire tmp23434;
  wire tmp23435;
  wire tmp23436;
  wire tmp23437;
  wire tmp23438;
  wire tmp23439;
  wire tmp23440;
  wire tmp23441;
  wire tmp23442;
  wire tmp23443;
  wire tmp23444;
  wire tmp23445;
  wire tmp23446;
  wire tmp23447;
  wire tmp23448;
  wire tmp23449;
  wire tmp23450;
  wire tmp23451;
  wire tmp23452;
  wire tmp23453;
  wire tmp23454;
  wire tmp23455;
  wire tmp23456;
  wire tmp23457;
  wire tmp23458;
  wire tmp23459;
  wire tmp23460;
  wire tmp23461;
  wire tmp23462;
  wire tmp23463;
  wire tmp23464;
  wire tmp23465;
  wire tmp23466;
  wire tmp23467;
  wire tmp23468;
  wire tmp23469;
  wire tmp23470;
  wire tmp23471;
  wire tmp23472;
  wire tmp23473;
  wire tmp23474;
  wire tmp23475;
  wire tmp23476;
  wire tmp23477;
  wire tmp23478;
  wire tmp23479;
  wire tmp23480;
  wire tmp23481;
  wire tmp23482;
  wire tmp23483;
  wire tmp23484;
  wire tmp23485;
  wire tmp23486;
  wire tmp23487;
  wire tmp23488;
  wire tmp23489;
  wire tmp23490;
  wire tmp23491;
  wire tmp23492;
  wire tmp23493;
  wire tmp23494;
  wire tmp23495;
  wire tmp23496;
  wire tmp23497;
  wire tmp23498;
  wire tmp23499;
  wire tmp23500;
  wire tmp23501;
  wire tmp23502;
  wire tmp23503;
  wire tmp23504;
  wire tmp23505;
  wire tmp23506;
  wire tmp23507;
  wire tmp23508;
  wire tmp23509;
  wire tmp23510;
  wire tmp23511;
  wire tmp23512;
  wire tmp23513;
  wire tmp23514;
  wire tmp23515;
  wire tmp23516;
  wire tmp23517;
  wire tmp23518;
  wire tmp23519;
  wire tmp23520;
  wire tmp23521;
  wire tmp23522;
  wire tmp23523;
  wire tmp23524;
  wire tmp23525;
  wire tmp23526;
  wire tmp23527;
  wire tmp23528;
  wire tmp23529;
  wire tmp23530;
  wire tmp23531;
  wire tmp23532;
  wire tmp23533;
  wire tmp23534;
  wire tmp23535;
  wire tmp23536;
  wire tmp23537;
  wire tmp23538;
  wire tmp23539;
  wire tmp23540;
  wire tmp23541;
  wire tmp23542;
  wire tmp23543;
  wire tmp23544;
  wire tmp23545;
  wire tmp23546;
  wire tmp23547;
  wire tmp23548;
  wire tmp23549;
  wire tmp23550;
  wire tmp23551;
  wire tmp23552;
  wire tmp23553;
  wire tmp23554;
  wire tmp23555;
  wire tmp23556;
  wire tmp23557;
  wire tmp23558;
  wire tmp23559;
  wire tmp23560;
  wire tmp23561;
  wire tmp23562;
  wire tmp23563;
  wire tmp23564;
  wire tmp23565;
  wire tmp23566;
  wire tmp23567;
  wire tmp23568;
  wire tmp23569;
  wire tmp23570;
  wire tmp23571;
  wire tmp23572;
  wire tmp23573;
  wire tmp23574;
  wire tmp23575;
  wire tmp23576;
  wire tmp23577;
  wire tmp23578;
  wire tmp23579;
  wire tmp23580;
  wire tmp23581;
  wire tmp23582;
  wire tmp23583;
  wire tmp23584;
  wire tmp23585;
  wire tmp23586;
  wire tmp23587;
  wire tmp23588;
  wire tmp23589;
  wire tmp23590;
  wire tmp23591;
  wire tmp23592;
  wire tmp23593;
  wire tmp23594;
  wire tmp23595;
  wire tmp23596;
  wire tmp23597;
  wire tmp23598;
  wire tmp23599;
  wire tmp23600;
  wire tmp23601;
  wire tmp23602;
  wire tmp23603;
  wire tmp23604;
  wire tmp23605;
  wire tmp23606;
  wire tmp23607;
  wire tmp23608;
  wire tmp23609;
  wire tmp23610;
  wire tmp23611;
  wire tmp23612;
  wire tmp23613;
  wire tmp23614;
  wire tmp23615;
  wire tmp23616;
  wire tmp23617;
  wire tmp23618;
  wire tmp23619;
  wire tmp23620;
  wire tmp23621;
  wire tmp23622;
  wire tmp23623;
  wire tmp23624;
  wire tmp23625;
  wire tmp23626;
  wire tmp23627;
  wire tmp23628;
  wire tmp23629;
  wire tmp23630;
  wire tmp23631;
  wire tmp23632;
  wire tmp23633;
  wire tmp23634;
  wire tmp23635;
  wire tmp23636;
  wire tmp23637;
  wire tmp23638;
  wire tmp23639;
  wire tmp23640;
  wire tmp23641;
  wire tmp23642;
  wire tmp23643;
  wire tmp23644;
  wire tmp23645;
  wire tmp23646;
  wire tmp23647;
  wire tmp23648;
  wire tmp23649;
  wire tmp23650;
  wire tmp23651;
  wire tmp23652;
  wire tmp23653;
  wire tmp23654;
  wire tmp23655;
  wire tmp23656;
  wire tmp23657;
  wire tmp23658;
  wire tmp23659;
  wire tmp23660;
  wire tmp23661;
  wire tmp23662;
  wire tmp23663;
  wire tmp23664;
  wire tmp23665;
  wire tmp23666;
  wire tmp23667;
  wire tmp23668;
  wire tmp23669;
  wire tmp23670;
  wire tmp23671;
  wire tmp23672;
  wire tmp23673;
  wire tmp23674;
  wire tmp23675;
  wire tmp23676;
  wire tmp23677;
  wire tmp23678;
  wire tmp23679;
  wire tmp23680;
  wire tmp23681;
  wire tmp23682;
  wire tmp23683;
  wire tmp23684;
  wire tmp23685;
  wire tmp23686;
  wire tmp23687;
  wire tmp23688;
  wire tmp23689;
  wire tmp23690;
  wire tmp23691;
  wire tmp23692;
  wire tmp23693;
  wire tmp23694;
  wire tmp23695;
  wire tmp23696;
  wire tmp23697;
  wire tmp23698;
  wire tmp23699;
  wire tmp23700;
  wire tmp23701;
  wire tmp23702;
  wire tmp23703;
  wire tmp23704;
  wire tmp23705;
  wire tmp23706;
  wire tmp23707;
  wire tmp23708;
  wire tmp23709;
  wire tmp23710;
  wire tmp23711;
  wire tmp23712;
  wire tmp23713;
  wire tmp23714;
  wire tmp23715;
  wire tmp23716;
  wire tmp23717;
  wire tmp23718;
  wire tmp23719;
  wire tmp23720;
  wire tmp23721;
  wire tmp23722;
  wire tmp23723;
  wire tmp23724;
  wire tmp23725;
  wire tmp23726;
  wire tmp23727;
  wire tmp23728;
  wire tmp23729;
  wire tmp23730;
  wire tmp23731;
  wire tmp23732;
  wire tmp23733;
  wire tmp23734;
  wire tmp23735;
  wire tmp23736;
  wire tmp23737;
  wire tmp23738;
  wire tmp23739;
  wire tmp23740;
  wire tmp23741;
  wire tmp23742;
  wire tmp23743;
  wire tmp23744;
  wire tmp23745;
  wire tmp23746;
  wire tmp23747;
  wire tmp23748;
  wire tmp23749;
  wire tmp23750;
  wire tmp23751;
  wire tmp23752;
  wire tmp23753;
  wire tmp23754;
  wire tmp23755;
  wire tmp23756;
  wire tmp23757;
  wire tmp23758;
  wire tmp23759;
  wire tmp23760;
  wire tmp23761;
  wire tmp23762;
  wire tmp23763;
  wire tmp23764;
  wire tmp23765;
  wire tmp23766;
  wire tmp23767;
  wire tmp23768;
  wire tmp23769;
  wire tmp23770;
  wire tmp23771;
  wire tmp23772;
  wire tmp23773;
  wire tmp23774;
  wire tmp23775;
  wire tmp23776;
  wire tmp23777;
  wire tmp23778;
  wire tmp23779;
  wire tmp23780;
  wire tmp23781;
  wire tmp23782;
  wire tmp23783;
  wire tmp23784;
  wire tmp23785;
  wire tmp23786;
  wire tmp23787;
  wire tmp23788;
  wire tmp23789;
  wire tmp23790;
  wire tmp23791;
  wire tmp23792;
  wire tmp23793;
  wire tmp23794;
  wire tmp23795;
  wire tmp23796;
  wire tmp23797;
  wire tmp23798;
  wire tmp23799;
  wire tmp23800;
  wire tmp23801;
  wire tmp23802;
  wire tmp23803;
  wire tmp23804;
  wire tmp23805;
  wire tmp23806;
  wire tmp23807;
  wire tmp23808;
  wire tmp23809;
  wire tmp23810;
  wire tmp23811;
  wire tmp23812;
  wire tmp23813;
  wire tmp23814;
  wire tmp23815;
  wire tmp23816;
  wire tmp23817;
  wire tmp23818;
  wire tmp23819;
  wire tmp23820;
  wire tmp23821;
  wire tmp23822;
  wire tmp23823;
  wire tmp23824;
  wire tmp23825;
  wire tmp23826;
  wire tmp23827;
  wire tmp23828;
  wire tmp23829;
  wire tmp23830;
  wire tmp23831;
  wire tmp23832;
  wire tmp23833;
  wire tmp23834;
  wire tmp23835;
  wire tmp23836;
  wire tmp23837;
  wire tmp23838;
  wire tmp23839;
  wire tmp23840;
  wire tmp23841;
  wire tmp23842;
  wire tmp23843;
  wire tmp23844;
  wire tmp23845;
  wire tmp23846;
  wire tmp23847;
  wire tmp23848;
  wire tmp23849;
  wire tmp23850;
  wire tmp23851;
  wire tmp23852;
  wire tmp23853;
  wire tmp23854;
  wire tmp23855;
  wire tmp23856;
  wire tmp23857;
  wire tmp23858;
  wire tmp23859;
  wire tmp23860;
  wire tmp23861;
  wire tmp23862;
  wire tmp23863;
  wire tmp23864;
  wire tmp23865;
  wire tmp23866;
  wire tmp23867;
  wire tmp23868;
  wire tmp23869;
  wire tmp23870;
  wire tmp23871;
  wire tmp23872;
  wire tmp23873;
  wire tmp23874;
  wire tmp23875;
  wire tmp23876;
  wire tmp23877;
  wire tmp23878;
  wire tmp23879;
  wire tmp23880;
  wire tmp23881;
  wire tmp23882;
  wire tmp23883;
  wire tmp23884;
  wire tmp23885;
  wire tmp23886;
  wire tmp23887;
  wire tmp23888;
  wire tmp23889;
  wire tmp23890;
  wire tmp23891;
  wire tmp23892;
  wire tmp23893;
  wire tmp23894;
  wire tmp23895;
  wire tmp23896;
  wire tmp23897;
  wire tmp23898;
  wire tmp23899;
  wire tmp23900;
  wire tmp23901;
  wire tmp23902;
  wire tmp23903;
  wire tmp23904;
  wire tmp23905;
  wire tmp23906;
  wire tmp23907;
  wire tmp23908;
  wire tmp23909;
  wire tmp23910;
  wire tmp23911;
  wire tmp23912;
  wire tmp23913;
  wire tmp23914;
  wire tmp23915;
  wire tmp23916;
  wire tmp23917;
  wire tmp23918;
  wire tmp23919;
  wire tmp23920;
  wire tmp23921;
  wire tmp23922;
  wire tmp23923;
  wire tmp23924;
  wire tmp23925;
  wire tmp23926;
  wire tmp23927;
  wire tmp23928;
  wire tmp23929;
  wire tmp23930;
  wire tmp23931;
  wire tmp23932;
  wire tmp23933;
  wire tmp23934;
  wire tmp23935;
  wire tmp23936;
  wire tmp23937;
  wire tmp23938;
  wire tmp23939;
  wire tmp23940;
  wire tmp23941;
  wire tmp23942;
  wire tmp23943;
  wire tmp23944;
  wire tmp23945;
  wire tmp23946;
  wire tmp23947;
  wire tmp23948;
  wire tmp23949;
  wire tmp23950;
  wire tmp23951;
  wire tmp23952;
  wire tmp23953;
  wire tmp23954;
  wire tmp23955;
  wire tmp23956;
  wire tmp23957;
  wire tmp23958;
  wire tmp23959;
  wire tmp23960;
  wire tmp23961;
  wire tmp23962;
  wire tmp23963;
  wire tmp23964;
  wire tmp23965;
  wire tmp23966;
  wire tmp23967;
  wire tmp23968;
  wire tmp23969;
  wire tmp23970;
  wire tmp23971;
  wire tmp23972;
  wire tmp23973;
  wire tmp23974;
  wire tmp23975;
  wire tmp23976;
  wire tmp23977;
  wire tmp23978;
  wire tmp23979;
  wire tmp23980;
  wire tmp23981;
  wire tmp23982;
  wire tmp23983;
  wire tmp23984;
  wire tmp23985;
  wire tmp23986;
  wire tmp23987;
  wire tmp23988;
  wire tmp23989;
  wire tmp23990;
  wire tmp23991;
  wire tmp23992;
  wire tmp23993;
  wire tmp23994;
  wire tmp23995;
  wire tmp23996;
  wire tmp23997;
  wire tmp23998;
  wire tmp23999;
  wire tmp24000;
  wire tmp24001;
  wire tmp24002;
  wire tmp24003;
  wire tmp24004;
  wire tmp24005;
  wire tmp24006;
  wire tmp24007;
  wire tmp24008;
  wire tmp24009;
  wire tmp24010;
  wire tmp24011;
  wire tmp24012;
  wire tmp24013;
  wire tmp24014;
  wire tmp24015;
  wire tmp24016;
  wire tmp24017;
  wire tmp24018;
  wire tmp24019;
  wire tmp24020;
  wire tmp24021;
  wire tmp24022;
  wire tmp24023;
  wire tmp24024;
  wire tmp24025;
  wire tmp24026;
  wire tmp24027;
  wire tmp24028;
  wire tmp24029;
  wire tmp24030;
  wire tmp24031;
  wire tmp24032;
  wire tmp24033;
  wire tmp24034;
  wire tmp24035;
  wire tmp24036;
  wire tmp24037;
  wire tmp24038;
  wire tmp24039;
  wire tmp24040;
  wire tmp24041;
  wire tmp24042;
  wire tmp24043;
  wire tmp24044;
  wire tmp24045;
  wire tmp24046;
  wire tmp24047;
  wire tmp24048;
  wire tmp24049;
  wire tmp24050;
  wire tmp24051;
  wire tmp24052;
  wire tmp24053;
  wire tmp24054;
  wire tmp24055;
  wire tmp24056;
  wire tmp24057;
  wire tmp24058;
  wire tmp24059;
  wire tmp24060;
  wire tmp24061;
  wire tmp24062;
  wire tmp24063;
  wire tmp24064;
  wire tmp24065;
  wire tmp24066;
  wire tmp24067;
  wire tmp24068;
  wire tmp24069;
  wire tmp24070;
  wire tmp24071;
  wire tmp24072;
  wire tmp24073;
  wire tmp24074;
  wire tmp24075;
  wire tmp24076;
  wire tmp24077;
  wire tmp24078;
  wire tmp24079;
  wire tmp24080;
  wire tmp24081;
  wire tmp24082;
  wire tmp24083;
  wire tmp24084;
  wire tmp24085;
  wire tmp24086;
  wire tmp24087;
  wire tmp24088;
  wire tmp24089;
  wire tmp24090;
  wire tmp24091;
  wire tmp24092;
  wire tmp24093;
  wire tmp24094;
  wire tmp24095;
  wire tmp24096;
  wire tmp24097;
  wire tmp24098;
  wire tmp24099;
  wire tmp24100;
  wire tmp24101;
  wire tmp24102;
  wire tmp24103;
  wire tmp24104;
  wire tmp24105;
  wire tmp24106;
  wire tmp24107;
  wire tmp24108;
  wire tmp24109;
  wire tmp24110;
  wire tmp24111;
  wire tmp24112;
  wire tmp24113;
  wire tmp24114;
  wire tmp24115;
  wire tmp24116;
  wire tmp24117;
  wire tmp24118;
  wire tmp24119;
  wire tmp24120;
  wire tmp24121;
  wire tmp24122;
  wire tmp24123;
  wire tmp24124;
  wire tmp24125;
  wire tmp24126;
  wire tmp24127;
  wire tmp24128;
  wire tmp24129;
  wire tmp24130;
  wire tmp24131;
  wire tmp24132;
  wire tmp24133;
  wire tmp24134;
  wire tmp24135;
  wire tmp24136;
  wire tmp24137;
  wire tmp24138;
  wire tmp24139;
  wire tmp24140;
  wire tmp24141;
  wire tmp24142;
  wire tmp24143;
  wire tmp24144;
  wire tmp24145;
  wire tmp24146;
  wire tmp24147;
  wire tmp24148;
  wire tmp24149;
  wire tmp24150;
  wire tmp24151;
  wire tmp24152;
  wire tmp24153;
  wire tmp24154;
  wire tmp24155;
  wire tmp24156;
  wire tmp24157;
  wire tmp24158;
  wire tmp24159;
  wire tmp24160;
  wire tmp24161;
  wire tmp24162;
  wire tmp24163;
  wire tmp24164;
  wire tmp24165;
  wire tmp24166;
  wire tmp24167;
  wire tmp24168;
  wire tmp24169;
  wire tmp24170;
  wire tmp24171;
  wire tmp24172;
  wire tmp24173;
  wire tmp24174;
  wire tmp24175;
  wire tmp24176;
  wire tmp24177;
  wire tmp24178;
  wire tmp24179;
  wire tmp24180;
  wire tmp24181;
  wire tmp24182;
  wire tmp24183;
  wire tmp24184;
  wire tmp24185;
  wire tmp24186;
  wire tmp24187;
  wire tmp24188;
  wire tmp24189;
  wire tmp24190;
  wire tmp24191;
  wire tmp24192;
  wire tmp24193;
  wire tmp24194;
  wire tmp24195;
  wire tmp24196;
  wire tmp24197;
  wire tmp24198;
  wire tmp24199;
  wire tmp24200;
  wire tmp24201;
  wire tmp24202;
  wire tmp24203;
  wire tmp24204;
  wire tmp24205;
  wire tmp24206;
  wire tmp24207;
  wire tmp24208;
  wire tmp24209;
  wire tmp24210;
  wire tmp24211;
  wire tmp24212;
  wire tmp24213;
  wire tmp24214;
  wire tmp24215;
  wire tmp24216;
  wire tmp24217;
  wire tmp24218;
  wire tmp24219;
  wire tmp24220;
  wire tmp24221;
  wire tmp24222;
  wire tmp24223;
  wire tmp24224;
  wire tmp24225;
  wire tmp24226;
  wire tmp24227;
  wire tmp24228;
  wire tmp24229;
  wire tmp24230;
  wire tmp24231;
  wire tmp24232;
  wire tmp24233;
  wire tmp24234;
  wire tmp24235;
  wire tmp24236;
  wire tmp24237;
  wire tmp24238;
  wire tmp24239;
  wire tmp24240;
  wire tmp24241;
  wire tmp24242;
  wire tmp24243;
  wire tmp24244;
  wire tmp24245;
  wire tmp24246;
  wire tmp24247;
  wire tmp24248;
  wire tmp24249;
  wire tmp24250;
  wire tmp24251;
  wire tmp24252;
  wire tmp24253;
  wire tmp24254;
  wire tmp24255;
  wire tmp24256;
  wire tmp24257;
  wire tmp24258;
  wire tmp24259;
  wire tmp24260;
  wire tmp24261;
  wire tmp24262;
  wire tmp24263;
  wire tmp24264;
  wire tmp24265;
  wire tmp24266;
  wire tmp24267;
  wire tmp24268;
  wire tmp24269;
  wire tmp24270;
  wire tmp24271;
  wire tmp24272;
  wire tmp24273;
  wire tmp24274;
  wire tmp24275;
  wire tmp24276;
  wire tmp24277;
  wire tmp24278;
  wire tmp24279;
  wire tmp24280;
  wire tmp24281;
  wire tmp24282;
  wire tmp24283;
  wire tmp24284;
  wire tmp24285;
  wire tmp24286;
  wire tmp24287;
  wire tmp24288;
  wire tmp24289;
  wire tmp24290;
  wire tmp24291;
  wire tmp24292;
  wire tmp24293;
  wire tmp24294;
  wire tmp24295;
  wire tmp24296;
  wire tmp24297;
  wire tmp24298;
  wire tmp24299;
  wire tmp24300;
  wire tmp24301;
  wire tmp24302;
  wire tmp24303;
  wire tmp24304;
  wire tmp24305;
  wire tmp24306;
  wire tmp24307;
  wire tmp24308;
  wire tmp24309;
  wire tmp24310;
  wire tmp24311;
  wire tmp24312;
  wire tmp24313;
  wire tmp24314;
  wire tmp24315;
  wire tmp24316;
  wire tmp24317;
  wire tmp24318;
  wire tmp24319;
  wire tmp24320;
  wire tmp24321;
  wire tmp24322;
  wire tmp24323;
  wire tmp24324;
  wire tmp24325;
  wire tmp24326;
  wire tmp24327;
  wire tmp24328;
  wire tmp24329;
  wire tmp24330;
  wire tmp24331;
  wire tmp24332;
  wire tmp24333;
  wire tmp24334;
  wire tmp24335;
  wire tmp24336;
  wire tmp24337;
  wire tmp24338;
  wire tmp24339;
  wire tmp24340;
  wire tmp24341;
  wire tmp24342;
  wire tmp24343;
  wire tmp24344;
  wire tmp24345;
  wire tmp24346;
  wire tmp24347;
  wire tmp24348;
  wire tmp24349;
  wire tmp24350;
  wire tmp24351;
  wire tmp24352;
  wire tmp24353;
  wire tmp24354;
  wire tmp24355;
  wire tmp24356;
  wire tmp24357;
  wire tmp24358;
  wire tmp24359;
  wire tmp24360;
  wire tmp24361;
  wire tmp24362;
  wire tmp24363;
  wire tmp24364;
  wire tmp24365;
  wire tmp24366;
  wire tmp24367;
  wire tmp24368;
  wire tmp24369;
  wire tmp24370;
  wire tmp24371;
  wire tmp24372;
  wire tmp24373;
  wire tmp24374;
  wire tmp24375;
  wire tmp24376;
  wire tmp24377;
  wire tmp24378;
  wire tmp24379;
  wire tmp24380;
  wire tmp24381;
  wire tmp24382;
  wire tmp24383;
  wire tmp24384;
  wire tmp24385;
  wire tmp24386;
  wire tmp24387;
  wire tmp24388;
  wire tmp24389;
  wire tmp24390;
  wire tmp24391;
  wire tmp24392;
  wire tmp24393;
  wire tmp24394;
  wire tmp24395;
  wire tmp24396;
  wire tmp24397;
  wire tmp24398;
  wire tmp24399;
  wire tmp24400;
  wire tmp24401;
  wire tmp24402;
  wire tmp24403;
  wire tmp24404;
  wire tmp24405;
  wire tmp24406;
  wire tmp24407;
  wire tmp24408;
  wire tmp24409;
  wire tmp24410;
  wire tmp24411;
  wire tmp24412;
  wire tmp24413;
  wire tmp24414;
  wire tmp24415;
  wire tmp24416;
  wire tmp24417;
  wire tmp24418;
  wire tmp24419;
  wire tmp24420;
  wire tmp24421;
  wire tmp24422;
  wire tmp24423;
  wire tmp24424;
  wire tmp24425;
  wire tmp24426;
  wire tmp24427;
  wire tmp24428;
  wire tmp24429;
  wire tmp24430;
  wire tmp24431;
  wire tmp24432;
  wire tmp24433;
  wire tmp24434;
  wire tmp24435;
  wire tmp24436;
  wire tmp24437;
  wire tmp24438;
  wire tmp24439;
  wire tmp24440;
  wire tmp24441;
  wire tmp24442;
  wire tmp24443;
  wire tmp24444;
  wire tmp24445;
  wire tmp24446;
  wire tmp24447;
  wire tmp24448;
  wire tmp24449;
  wire tmp24450;
  wire tmp24451;
  wire tmp24452;
  wire tmp24453;
  wire tmp24454;
  wire tmp24455;
  wire tmp24456;
  wire tmp24457;
  wire tmp24458;
  wire tmp24459;
  wire tmp24460;
  wire tmp24461;
  wire tmp24462;
  wire tmp24463;
  wire tmp24464;
  wire tmp24465;
  wire tmp24466;
  wire tmp24467;
  wire tmp24468;
  wire tmp24469;
  wire tmp24470;
  wire tmp24471;
  wire tmp24472;
  wire tmp24473;
  wire tmp24474;
  wire tmp24475;
  wire tmp24476;
  wire tmp24477;
  wire tmp24478;
  wire tmp24479;
  wire tmp24480;
  wire tmp24481;
  wire tmp24482;
  wire tmp24483;
  wire tmp24484;
  wire tmp24485;
  wire tmp24486;
  wire tmp24487;
  wire tmp24488;
  wire tmp24489;
  wire tmp24490;
  wire tmp24491;
  wire tmp24492;
  wire tmp24493;
  wire tmp24494;
  wire tmp24495;
  wire tmp24496;
  wire tmp24497;
  wire tmp24498;
  wire tmp24499;
  wire tmp24500;
  wire tmp24501;
  wire tmp24502;
  wire tmp24503;
  wire tmp24504;
  wire tmp24505;
  wire tmp24506;
  wire tmp24507;
  wire tmp24508;
  wire tmp24509;
  wire tmp24510;
  wire tmp24511;
  wire tmp24512;
  wire tmp24513;
  wire tmp24514;
  wire tmp24515;
  wire tmp24516;
  wire tmp24517;
  wire tmp24518;
  wire tmp24519;
  wire tmp24520;
  wire tmp24521;
  wire tmp24522;
  wire tmp24523;
  wire tmp24524;
  wire tmp24525;
  wire tmp24526;
  wire tmp24527;
  wire tmp24528;
  wire tmp24529;
  wire tmp24530;
  wire tmp24531;
  wire tmp24532;
  wire tmp24533;
  wire tmp24534;
  wire tmp24535;
  wire tmp24536;
  wire tmp24537;
  wire tmp24538;
  wire tmp24539;
  wire tmp24540;
  wire tmp24541;
  wire tmp24542;
  wire tmp24543;
  wire tmp24544;
  wire tmp24545;
  wire tmp24546;
  wire tmp24547;
  wire tmp24548;
  wire tmp24549;
  wire tmp24550;
  wire tmp24551;
  wire tmp24552;
  wire tmp24553;
  wire tmp24554;
  wire tmp24555;
  wire tmp24556;
  wire tmp24557;
  wire tmp24558;
  wire tmp24559;
  wire tmp24560;
  wire tmp24561;
  wire tmp24562;
  wire tmp24563;
  wire tmp24564;
  wire tmp24565;
  wire tmp24566;
  wire tmp24567;
  wire tmp24568;
  wire tmp24569;
  wire tmp24570;
  wire tmp24571;
  wire tmp24572;
  wire tmp24573;
  wire tmp24574;
  wire tmp24575;
  wire tmp24576;
  wire tmp24577;
  wire tmp24578;
  wire tmp24579;
  wire tmp24580;
  wire tmp24581;
  wire tmp24582;
  wire tmp24583;
  wire tmp24584;
  wire tmp24585;
  wire tmp24586;
  wire tmp24587;
  wire tmp24588;
  wire tmp24589;
  wire tmp24590;
  wire tmp24591;
  wire tmp24592;
  wire tmp24593;
  wire tmp24594;
  wire tmp24595;
  wire tmp24596;
  wire tmp24597;
  wire tmp24598;
  wire tmp24599;
  wire tmp24600;
  wire tmp24601;
  wire tmp24602;
  wire tmp24603;
  wire tmp24604;
  wire tmp24605;
  wire tmp24606;
  wire tmp24607;
  wire tmp24608;
  wire tmp24609;
  wire tmp24610;
  wire tmp24611;
  wire tmp24612;
  wire tmp24613;
  wire tmp24614;
  wire tmp24615;
  wire tmp24616;
  wire tmp24617;
  wire tmp24618;
  wire tmp24619;
  wire tmp24620;
  wire tmp24621;
  wire tmp24622;
  wire tmp24623;
  wire tmp24624;
  wire tmp24625;
  wire tmp24626;
  wire tmp24627;
  wire tmp24628;
  wire tmp24629;
  wire tmp24630;
  wire tmp24631;
  wire tmp24632;
  wire tmp24633;
  wire tmp24634;
  wire tmp24635;
  wire tmp24636;
  wire tmp24637;
  wire tmp24638;
  wire tmp24639;
  wire tmp24640;
  wire tmp24641;
  wire tmp24642;
  wire tmp24643;
  wire tmp24644;
  wire tmp24645;
  wire tmp24646;
  wire tmp24647;
  wire tmp24648;
  wire tmp24649;
  wire tmp24650;
  wire tmp24651;
  wire tmp24652;
  wire tmp24653;
  wire tmp24654;
  wire tmp24655;
  wire tmp24656;
  wire tmp24657;
  wire tmp24658;
  wire tmp24659;
  wire tmp24660;
  wire tmp24661;
  wire tmp24662;
  wire tmp24663;
  wire tmp24664;
  wire tmp24665;
  wire tmp24666;
  wire tmp24667;
  wire tmp24668;
  wire tmp24669;
  wire tmp24670;
  wire tmp24671;
  wire tmp24672;
  wire tmp24673;
  wire tmp24674;
  wire tmp24675;
  wire tmp24676;
  wire tmp24677;
  wire tmp24678;
  wire tmp24679;
  wire tmp24680;
  wire tmp24681;
  wire tmp24682;
  wire tmp24683;
  wire tmp24684;
  wire tmp24685;
  wire tmp24686;
  wire tmp24687;
  wire tmp24688;
  wire tmp24689;
  wire tmp24690;
  wire tmp24691;
  wire tmp24692;
  wire tmp24693;
  wire tmp24694;
  wire tmp24695;
  wire tmp24696;
  wire tmp24697;
  wire tmp24698;
  wire tmp24699;
  wire tmp24700;
  wire tmp24701;
  wire tmp24702;
  wire tmp24703;
  wire tmp24704;
  wire tmp24705;
  wire tmp24706;
  wire tmp24707;
  wire tmp24708;
  wire tmp24709;
  wire tmp24710;
  wire tmp24711;
  wire tmp24712;
  wire tmp24713;
  wire tmp24714;
  wire tmp24715;
  wire tmp24716;
  wire tmp24717;
  wire tmp24718;
  wire tmp24719;
  wire tmp24720;
  wire tmp24721;
  wire tmp24722;
  wire tmp24723;
  wire tmp24724;
  wire tmp24725;
  wire tmp24726;
  wire tmp24727;
  wire tmp24728;
  wire tmp24729;
  wire tmp24730;
  wire tmp24731;
  wire tmp24732;
  wire tmp24733;
  wire tmp24734;
  wire tmp24735;
  wire tmp24736;
  wire tmp24737;
  wire tmp24738;
  wire tmp24739;
  wire tmp24740;
  wire tmp24741;
  wire tmp24742;
  wire tmp24743;
  wire tmp24744;
  wire tmp24745;
  wire tmp24746;
  wire tmp24747;
  wire tmp24748;
  wire tmp24749;
  wire tmp24750;
  wire tmp24751;
  wire tmp24752;
  wire tmp24753;
  wire tmp24754;
  wire tmp24755;
  wire tmp24756;
  wire tmp24757;
  wire tmp24758;
  wire tmp24759;
  wire tmp24760;
  wire tmp24761;
  wire tmp24762;
  wire tmp24763;
  wire tmp24764;
  wire tmp24765;
  wire tmp24766;
  wire tmp24767;
  wire tmp24768;
  wire tmp24769;
  wire tmp24770;
  wire tmp24771;
  wire tmp24772;
  wire tmp24773;
  wire tmp24774;
  wire tmp24775;
  wire tmp24776;
  wire tmp24777;
  wire tmp24778;
  wire tmp24779;
  wire tmp24780;
  wire tmp24781;
  wire tmp24782;
  wire tmp24783;
  wire tmp24784;
  wire tmp24785;
  wire tmp24786;
  wire tmp24787;
  wire tmp24788;
  wire tmp24789;
  wire tmp24790;
  wire tmp24791;
  wire tmp24792;
  wire tmp24793;
  wire tmp24794;
  wire tmp24795;
  wire tmp24796;
  wire tmp24797;
  wire tmp24798;
  wire tmp24799;
  wire tmp24800;
  wire tmp24801;
  wire tmp24802;
  wire tmp24803;
  wire tmp24804;
  wire tmp24805;
  wire tmp24806;
  wire tmp24807;
  wire tmp24808;
  wire tmp24809;
  wire tmp24810;
  wire tmp24811;
  wire tmp24812;
  wire tmp24813;
  wire tmp24814;
  wire tmp24815;
  wire tmp24816;
  wire tmp24817;
  wire tmp24818;
  wire tmp24819;
  wire tmp24820;
  wire tmp24821;
  wire tmp24822;
  wire tmp24823;
  wire tmp24824;
  wire tmp24825;
  wire tmp24826;
  wire tmp24827;
  wire tmp24828;
  wire tmp24829;
  wire tmp24830;
  wire tmp24831;
  wire tmp24832;
  wire tmp24833;
  wire tmp24834;
  wire tmp24835;
  wire tmp24836;
  wire tmp24837;
  wire tmp24838;
  wire tmp24839;
  wire tmp24840;
  wire tmp24841;
  wire tmp24842;
  wire tmp24843;
  wire tmp24844;
  wire tmp24845;
  wire tmp24846;
  wire tmp24847;
  wire tmp24848;
  wire tmp24849;
  wire tmp24850;
  wire tmp24851;
  wire tmp24852;
  wire tmp24853;
  wire tmp24854;
  wire tmp24855;
  wire tmp24856;
  wire tmp24857;
  wire tmp24858;
  wire tmp24859;
  wire tmp24860;
  wire tmp24861;
  wire tmp24862;
  wire tmp24863;
  wire tmp24864;
  wire tmp24865;
  wire tmp24866;
  wire tmp24867;
  wire tmp24868;
  wire tmp24869;
  wire tmp24870;
  wire tmp24871;
  wire tmp24872;
  wire tmp24873;
  wire tmp24874;
  wire tmp24875;
  wire tmp24876;
  wire tmp24877;
  wire tmp24878;
  wire tmp24879;
  wire tmp24880;
  wire tmp24881;
  wire tmp24882;
  wire tmp24883;
  wire tmp24884;
  wire tmp24885;
  wire tmp24886;
  wire tmp24887;
  wire tmp24888;
  wire tmp24889;
  wire tmp24890;
  wire tmp24891;
  wire tmp24892;
  wire tmp24893;
  wire tmp24894;
  wire tmp24895;
  wire tmp24896;
  wire tmp24897;
  wire tmp24898;
  wire tmp24899;
  wire tmp24900;
  wire tmp24901;
  wire tmp24902;
  wire tmp24903;
  wire tmp24904;
  wire tmp24905;
  wire tmp24906;
  wire tmp24907;
  wire tmp24908;
  wire tmp24909;
  wire tmp24910;
  wire tmp24911;
  wire tmp24912;
  wire tmp24913;
  wire tmp24914;
  wire tmp24915;
  wire tmp24916;
  wire tmp24917;
  wire tmp24918;
  wire tmp24919;
  wire tmp24920;
  wire tmp24921;
  wire tmp24922;
  wire tmp24923;
  wire tmp24924;
  wire tmp24925;
  wire tmp24926;
  wire tmp24927;
  wire tmp24928;
  wire tmp24929;
  wire tmp24930;
  wire tmp24931;
  wire tmp24932;
  wire tmp24933;
  wire tmp24934;
  wire tmp24935;
  wire tmp24936;
  wire tmp24937;
  wire tmp24938;
  wire tmp24939;
  wire tmp24940;
  wire tmp24941;
  wire tmp24942;
  wire tmp24943;
  wire tmp24944;
  wire tmp24945;
  wire tmp24946;
  wire tmp24947;
  wire tmp24948;
  wire tmp24949;
  wire tmp24950;
  wire tmp24951;
  wire tmp24952;
  wire tmp24953;
  wire tmp24954;
  wire tmp24955;
  wire tmp24956;
  wire tmp24957;
  wire tmp24958;
  wire tmp24959;
  wire tmp24960;
  wire tmp24961;
  wire tmp24962;
  wire tmp24963;
  wire tmp24964;
  wire tmp24965;
  wire tmp24966;
  wire tmp24967;
  wire tmp24968;
  wire tmp24969;
  wire tmp24970;
  wire tmp24971;
  wire tmp24972;
  wire tmp24973;
  wire tmp24974;
  wire tmp24975;
  wire tmp24976;
  wire tmp24977;
  wire tmp24978;
  wire tmp24979;
  wire tmp24980;
  wire tmp24981;
  wire tmp24982;
  wire tmp24983;
  wire tmp24984;
  wire tmp24985;
  wire tmp24986;
  wire tmp24987;
  wire tmp24988;
  wire tmp24989;
  wire tmp24990;
  wire tmp24991;
  wire tmp24992;
  wire tmp24993;
  wire tmp24994;
  wire tmp24995;
  wire tmp24996;
  wire tmp24997;
  wire tmp24998;
  wire tmp24999;
  wire tmp25000;
  wire tmp25001;
  wire tmp25002;
  wire tmp25003;
  wire tmp25004;
  wire tmp25005;
  wire tmp25006;
  wire tmp25007;
  wire tmp25008;
  wire tmp25009;
  wire tmp25010;
  wire tmp25011;
  wire tmp25012;
  wire tmp25013;
  wire tmp25014;
  wire tmp25015;
  wire tmp25016;
  wire tmp25017;
  wire tmp25018;
  wire tmp25019;
  wire tmp25020;
  wire tmp25021;
  wire tmp25022;
  wire tmp25023;
  wire tmp25024;
  wire tmp25025;
  wire tmp25026;
  wire tmp25027;
  wire tmp25028;
  wire tmp25029;
  wire tmp25030;
  wire tmp25031;
  wire tmp25032;
  wire tmp25033;
  wire tmp25034;
  wire tmp25035;
  wire tmp25036;
  wire tmp25037;
  wire tmp25038;
  wire tmp25039;
  wire tmp25040;
  wire tmp25041;
  wire tmp25042;
  wire tmp25043;
  wire tmp25044;
  wire tmp25045;
  wire tmp25046;
  wire tmp25047;
  wire tmp25048;
  wire tmp25049;
  wire tmp25050;
  wire tmp25051;
  wire tmp25052;
  wire tmp25053;
  wire tmp25054;
  wire tmp25055;
  wire tmp25056;
  wire tmp25057;
  wire tmp25058;
  wire tmp25059;
  wire tmp25060;
  wire tmp25061;
  wire tmp25062;
  wire tmp25063;
  wire tmp25064;
  wire tmp25065;
  wire tmp25066;
  wire tmp25067;
  wire tmp25068;
  wire tmp25069;
  wire tmp25070;
  wire tmp25071;
  wire tmp25072;
  wire tmp25073;
  wire tmp25074;
  wire tmp25075;
  wire tmp25076;
  wire tmp25077;
  wire tmp25078;
  wire tmp25079;
  wire tmp25080;
  wire tmp25081;
  wire tmp25082;
  wire tmp25083;
  wire tmp25084;
  wire tmp25085;
  wire tmp25086;
  wire tmp25087;
  wire tmp25088;
  wire tmp25089;
  wire tmp25090;
  wire tmp25091;
  wire tmp25092;
  wire tmp25093;
  wire tmp25094;
  wire tmp25095;
  wire tmp25096;
  wire tmp25097;
  wire tmp25098;
  wire tmp25099;
  wire tmp25100;
  wire tmp25101;
  wire tmp25102;
  wire tmp25103;
  wire tmp25104;
  wire tmp25105;
  wire tmp25106;
  wire tmp25107;
  wire tmp25108;
  wire tmp25109;
  wire tmp25110;
  wire tmp25111;
  wire tmp25112;
  wire tmp25113;
  wire tmp25114;
  wire tmp25115;
  wire tmp25116;
  wire tmp25117;
  wire tmp25118;
  wire tmp25119;
  wire tmp25120;
  wire tmp25121;
  wire tmp25122;
  wire tmp25123;
  wire tmp25124;
  wire tmp25125;
  wire tmp25126;
  wire tmp25127;
  wire tmp25128;
  wire tmp25129;
  wire tmp25130;
  wire tmp25131;
  wire tmp25132;
  wire tmp25133;
  wire tmp25134;
  wire tmp25135;
  wire tmp25136;
  wire tmp25137;
  wire tmp25138;
  wire tmp25139;
  wire tmp25140;
  wire tmp25141;
  wire tmp25142;
  wire tmp25143;
  wire tmp25144;
  wire tmp25145;
  wire tmp25146;
  wire tmp25147;
  wire tmp25148;
  wire tmp25149;
  wire tmp25150;
  wire tmp25151;
  wire tmp25152;
  wire tmp25153;
  wire tmp25154;
  wire tmp25155;
  wire tmp25156;
  wire tmp25157;
  wire tmp25158;
  wire tmp25159;
  wire tmp25160;
  wire tmp25161;
  wire tmp25162;
  wire tmp25163;
  wire tmp25164;
  wire tmp25165;
  wire tmp25166;
  wire tmp25167;
  wire tmp25168;
  wire tmp25169;
  wire tmp25170;
  wire tmp25171;
  wire tmp25172;
  wire tmp25173;
  wire tmp25174;
  wire tmp25175;
  wire tmp25176;
  wire tmp25177;
  wire tmp25178;
  wire tmp25179;
  wire tmp25180;
  wire tmp25181;
  wire tmp25182;
  wire tmp25183;
  wire tmp25184;
  wire tmp25185;
  wire tmp25186;
  wire tmp25187;
  wire tmp25188;
  wire tmp25189;
  wire tmp25190;
  wire tmp25191;
  wire tmp25192;
  wire tmp25193;
  wire tmp25194;
  wire tmp25195;
  wire tmp25196;
  wire tmp25197;
  wire tmp25198;
  wire tmp25199;
  wire tmp25200;
  wire tmp25201;
  wire tmp25202;
  wire tmp25203;
  wire tmp25204;
  wire tmp25205;
  wire tmp25206;
  wire tmp25207;
  wire tmp25208;
  wire tmp25209;
  wire tmp25210;
  wire tmp25211;
  wire tmp25212;
  wire tmp25213;
  wire tmp25214;
  wire tmp25215;
  wire tmp25216;
  wire tmp25217;
  wire tmp25218;
  wire tmp25219;
  wire tmp25220;
  wire tmp25221;
  wire tmp25222;
  wire tmp25223;
  wire tmp25224;
  wire tmp25225;
  wire tmp25226;
  wire tmp25227;
  wire tmp25228;
  wire tmp25229;
  wire tmp25230;
  wire tmp25231;
  wire tmp25232;
  wire tmp25233;
  wire tmp25234;
  wire tmp25235;
  wire tmp25236;
  wire tmp25237;
  wire tmp25238;
  wire tmp25239;
  wire tmp25240;
  wire tmp25241;
  wire tmp25242;
  wire tmp25243;
  wire tmp25244;
  wire tmp25245;
  wire tmp25246;
  wire tmp25247;
  wire tmp25248;
  wire tmp25249;
  wire tmp25250;
  wire tmp25251;
  wire tmp25252;
  wire tmp25253;
  wire tmp25254;
  wire tmp25255;
  wire tmp25256;
  wire tmp25257;
  wire tmp25258;
  wire tmp25259;
  wire tmp25260;
  wire tmp25261;
  wire tmp25262;
  wire tmp25263;
  wire tmp25264;
  wire tmp25265;
  wire tmp25266;
  wire tmp25267;
  wire tmp25268;
  wire tmp25269;
  wire tmp25270;
  wire tmp25271;
  wire tmp25272;
  wire tmp25273;
  wire tmp25274;
  wire tmp25275;
  wire tmp25276;
  wire tmp25277;
  wire tmp25278;
  wire tmp25279;
  wire tmp25280;
  wire tmp25281;
  wire tmp25282;
  wire tmp25283;
  wire tmp25284;
  wire tmp25285;
  wire tmp25286;
  wire tmp25287;
  wire tmp25288;
  wire tmp25289;
  wire tmp25290;
  wire tmp25291;
  wire tmp25292;
  wire tmp25293;
  wire tmp25294;
  wire tmp25295;
  wire tmp25296;
  wire tmp25297;
  wire tmp25298;
  wire tmp25299;
  wire tmp25300;
  wire tmp25301;
  wire tmp25302;
  wire tmp25303;
  wire tmp25304;
  wire tmp25305;
  wire tmp25306;
  wire tmp25307;
  wire tmp25308;
  wire tmp25309;
  wire tmp25310;
  wire tmp25311;
  wire tmp25312;
  wire tmp25313;
  wire tmp25314;
  wire tmp25315;
  wire tmp25316;
  wire tmp25317;
  wire tmp25318;
  wire tmp25319;
  wire tmp25320;
  wire tmp25321;
  wire tmp25322;
  wire tmp25323;
  wire tmp25324;
  wire tmp25325;
  wire tmp25326;
  wire tmp25327;
  wire tmp25328;
  wire tmp25329;
  wire tmp25330;
  wire tmp25331;
  wire tmp25332;
  wire tmp25333;
  wire tmp25334;
  wire tmp25335;
  wire tmp25336;
  wire tmp25337;
  wire tmp25338;
  wire tmp25339;
  wire tmp25340;
  wire tmp25341;
  wire tmp25342;
  wire tmp25343;
  wire tmp25344;
  wire tmp25345;
  wire tmp25346;
  wire tmp25347;
  wire tmp25348;
  wire tmp25349;
  wire tmp25350;
  wire tmp25351;
  wire tmp25352;
  wire tmp25353;
  wire tmp25354;
  wire tmp25355;
  wire tmp25356;
  wire tmp25357;
  wire tmp25358;
  wire tmp25359;
  wire tmp25360;
  wire tmp25361;
  wire tmp25362;
  wire tmp25363;
  wire tmp25364;
  wire tmp25365;
  wire tmp25366;
  wire tmp25367;
  wire tmp25368;
  wire tmp25369;
  wire tmp25370;
  wire tmp25371;
  wire tmp25372;
  wire tmp25373;
  wire tmp25374;
  wire tmp25375;
  wire tmp25376;
  wire tmp25377;
  wire tmp25378;
  wire tmp25379;
  wire tmp25380;
  wire tmp25381;
  wire tmp25382;
  wire tmp25383;
  wire tmp25384;
  wire tmp25385;
  wire tmp25386;
  wire tmp25387;
  wire tmp25388;
  wire tmp25389;
  wire tmp25390;
  wire tmp25391;
  wire tmp25392;
  wire tmp25393;
  wire tmp25394;
  wire tmp25395;
  wire tmp25396;
  wire tmp25397;
  wire tmp25398;
  wire tmp25399;
  wire tmp25400;
  wire tmp25401;
  wire tmp25402;
  wire tmp25403;
  wire tmp25404;
  wire tmp25405;
  wire tmp25406;
  wire tmp25407;
  wire tmp25408;
  wire tmp25409;
  wire tmp25410;
  wire tmp25411;
  wire tmp25412;
  wire tmp25413;
  wire tmp25414;
  wire tmp25415;
  wire tmp25416;
  wire tmp25417;
  wire tmp25418;
  wire tmp25419;
  wire tmp25420;
  wire tmp25421;
  wire tmp25422;
  wire tmp25423;
  wire tmp25424;
  wire tmp25425;
  wire tmp25426;
  wire tmp25427;
  wire tmp25428;
  wire tmp25429;
  wire tmp25430;
  wire tmp25431;
  wire tmp25432;
  wire tmp25433;
  wire tmp25434;
  wire tmp25435;
  wire tmp25436;
  wire tmp25437;
  wire tmp25438;
  wire tmp25439;
  wire tmp25440;
  wire tmp25441;
  wire tmp25442;
  wire tmp25443;
  wire tmp25444;
  wire tmp25445;
  wire tmp25446;
  wire tmp25447;
  wire tmp25448;
  wire tmp25449;
  wire tmp25450;
  wire tmp25451;
  wire tmp25452;
  wire tmp25453;
  wire tmp25454;
  wire tmp25455;
  wire tmp25456;
  wire tmp25457;
  wire tmp25458;
  wire tmp25459;
  wire tmp25460;
  wire tmp25461;
  wire tmp25462;
  wire tmp25463;
  wire tmp25464;
  wire tmp25465;
  wire tmp25466;
  wire tmp25467;
  wire tmp25468;
  wire tmp25469;
  wire tmp25470;
  wire tmp25471;
  wire tmp25472;
  wire tmp25473;
  wire tmp25474;
  wire tmp25475;
  wire tmp25476;
  wire tmp25477;
  wire tmp25478;
  wire tmp25479;
  wire tmp25480;
  wire tmp25481;
  wire tmp25482;
  wire tmp25483;
  wire tmp25484;
  wire tmp25485;
  wire tmp25486;
  wire tmp25487;
  wire tmp25488;
  wire tmp25489;
  wire tmp25490;
  wire tmp25491;
  wire tmp25492;
  wire tmp25493;
  wire tmp25494;
  wire tmp25495;
  wire tmp25496;
  wire tmp25497;
  wire tmp25498;
  wire tmp25499;
  wire tmp25500;
  wire tmp25501;
  wire tmp25502;
  wire tmp25503;
  wire tmp25504;
  wire tmp25505;
  wire tmp25506;
  wire tmp25507;
  wire tmp25508;
  wire tmp25509;
  wire tmp25510;
  wire tmp25511;
  wire tmp25512;
  wire tmp25513;
  wire tmp25514;
  wire tmp25515;
  wire tmp25516;
  wire tmp25517;
  wire tmp25518;
  wire tmp25519;
  wire tmp25520;
  wire tmp25521;
  wire tmp25522;
  wire tmp25523;
  wire tmp25524;
  wire tmp25525;
  wire tmp25526;
  wire tmp25527;
  wire tmp25528;
  wire tmp25529;
  wire tmp25530;
  wire tmp25531;
  wire tmp25532;
  wire tmp25533;
  wire tmp25534;
  wire tmp25535;
  wire tmp25536;
  wire tmp25537;
  wire tmp25538;
  wire tmp25539;
  wire tmp25540;
  wire tmp25541;
  wire tmp25542;
  wire tmp25543;
  wire tmp25544;
  wire tmp25545;
  wire tmp25546;
  wire tmp25547;
  wire tmp25548;
  wire tmp25549;
  wire tmp25550;
  wire tmp25551;
  wire tmp25552;
  wire tmp25553;
  wire tmp25554;
  wire tmp25555;
  wire tmp25556;
  wire tmp25557;
  wire tmp25558;
  wire tmp25559;
  wire tmp25560;
  wire tmp25561;
  wire tmp25562;
  wire tmp25563;
  wire tmp25564;
  wire tmp25565;
  wire tmp25566;
  wire tmp25567;
  wire tmp25568;
  wire tmp25569;
  wire tmp25570;
  wire tmp25571;
  wire tmp25572;
  wire tmp25573;
  wire tmp25574;
  wire tmp25575;
  wire tmp25576;
  wire tmp25577;
  wire tmp25578;
  wire tmp25579;
  wire tmp25580;
  wire tmp25581;
  wire tmp25582;
  wire tmp25583;
  wire tmp25584;
  wire tmp25585;
  wire tmp25586;
  wire tmp25587;
  wire tmp25588;
  wire tmp25589;
  wire tmp25590;
  wire tmp25591;
  wire tmp25592;
  wire tmp25593;
  wire tmp25594;
  wire tmp25595;
  wire tmp25596;
  wire tmp25597;
  wire tmp25598;
  wire tmp25599;
  wire tmp25600;
  wire tmp25601;
  wire tmp25602;
  wire tmp25603;
  wire tmp25604;
  wire tmp25605;
  wire tmp25606;
  wire tmp25607;
  wire tmp25608;
  wire tmp25609;
  wire tmp25610;
  wire tmp25611;
  wire tmp25612;
  wire tmp25613;
  wire tmp25614;
  wire tmp25615;
  wire tmp25616;
  wire tmp25617;
  wire tmp25618;
  wire tmp25619;
  wire tmp25620;
  wire tmp25621;
  wire tmp25622;
  wire tmp25623;
  wire tmp25624;
  wire tmp25625;
  wire tmp25626;
  wire tmp25627;
  wire tmp25628;
  wire tmp25629;
  wire tmp25630;
  wire tmp25631;
  wire tmp25632;
  wire tmp25633;
  wire tmp25634;
  wire tmp25635;
  wire tmp25636;
  wire tmp25637;
  wire tmp25638;
  wire tmp25639;
  wire tmp25640;
  wire tmp25641;
  wire tmp25642;
  wire tmp25643;
  wire tmp25644;
  wire tmp25645;
  wire tmp25646;
  wire tmp25647;
  wire tmp25648;
  wire tmp25649;
  wire tmp25650;
  wire tmp25651;
  wire tmp25652;
  wire tmp25653;
  wire tmp25654;
  wire tmp25655;
  wire tmp25656;
  wire tmp25657;
  wire tmp25658;
  wire tmp25659;
  wire tmp25660;
  wire tmp25661;
  wire tmp25662;
  wire tmp25663;
  wire tmp25664;
  wire tmp25665;
  wire tmp25666;
  wire tmp25667;
  wire tmp25668;
  wire tmp25669;
  wire tmp25670;
  wire tmp25671;
  wire tmp25672;
  wire tmp25673;
  wire tmp25674;
  wire tmp25675;
  wire tmp25676;
  wire tmp25677;
  wire tmp25678;
  wire tmp25679;
  wire tmp25680;
  wire tmp25681;
  wire tmp25682;
  wire tmp25683;
  wire tmp25684;
  wire tmp25685;
  wire tmp25686;
  wire tmp25687;
  wire tmp25688;
  wire tmp25689;
  wire tmp25690;
  wire tmp25691;
  wire tmp25692;
  wire tmp25693;
  wire tmp25694;
  wire tmp25695;
  wire tmp25696;
  wire tmp25697;
  wire tmp25698;
  wire tmp25699;
  wire tmp25700;
  wire tmp25701;
  wire tmp25702;
  wire tmp25703;
  wire tmp25704;
  wire tmp25705;
  wire tmp25706;
  wire tmp25707;
  wire tmp25708;
  wire tmp25709;
  wire tmp25710;
  wire tmp25711;
  wire tmp25712;
  wire tmp25713;
  wire tmp25714;
  wire tmp25715;
  wire tmp25716;
  wire tmp25717;
  wire tmp25718;
  wire tmp25719;
  wire tmp25720;
  wire tmp25721;
  wire tmp25722;
  wire tmp25723;
  wire tmp25724;
  wire tmp25725;
  wire tmp25726;
  wire tmp25727;
  wire tmp25728;
  wire tmp25729;
  wire tmp25730;
  wire tmp25731;
  wire tmp25732;
  wire tmp25733;
  wire tmp25734;
  wire tmp25735;
  wire tmp25736;
  wire tmp25737;
  wire tmp25738;
  wire tmp25739;
  wire tmp25740;
  wire tmp25741;
  wire tmp25742;
  wire tmp25743;
  wire tmp25744;
  wire tmp25745;
  wire tmp25746;
  wire tmp25747;
  wire tmp25748;
  wire tmp25749;
  wire tmp25750;
  wire tmp25751;
  wire tmp25752;
  wire tmp25753;
  wire tmp25754;
  wire tmp25755;
  wire tmp25756;
  wire tmp25757;
  wire tmp25758;
  wire tmp25759;
  wire tmp25760;
  wire tmp25761;
  wire tmp25762;
  wire tmp25763;
  wire tmp25764;
  wire tmp25765;
  wire tmp25766;
  wire tmp25767;
  wire tmp25768;
  wire tmp25769;
  wire tmp25770;
  wire tmp25771;
  wire tmp25772;
  wire tmp25773;
  wire tmp25774;
  wire tmp25775;
  wire tmp25776;
  wire tmp25777;
  wire tmp25778;
  wire tmp25779;
  wire tmp25780;
  wire tmp25781;
  wire tmp25782;
  wire tmp25783;
  wire tmp25784;
  wire tmp25785;
  wire tmp25786;
  wire tmp25787;
  wire tmp25788;
  wire tmp25789;
  wire tmp25790;
  wire tmp25791;
  wire tmp25792;
  wire tmp25793;
  wire tmp25794;
  wire tmp25795;
  wire tmp25796;
  wire tmp25797;
  wire tmp25798;
  wire tmp25799;
  wire tmp25800;
  wire tmp25801;
  wire tmp25802;
  wire tmp25803;
  wire tmp25804;
  wire tmp25805;
  wire tmp25806;
  wire tmp25807;
  wire tmp25808;
  wire tmp25809;
  wire tmp25810;
  wire tmp25811;
  wire tmp25812;
  wire tmp25813;
  wire tmp25814;
  wire tmp25815;
  wire tmp25816;
  wire tmp25817;
  wire tmp25818;
  wire tmp25819;
  wire tmp25820;
  wire tmp25821;
  wire tmp25822;
  wire tmp25823;
  wire tmp25824;
  wire tmp25825;
  wire tmp25826;
  wire tmp25827;
  wire tmp25828;
  wire tmp25829;
  wire tmp25830;
  wire tmp25831;
  wire tmp25832;
  wire tmp25833;
  wire tmp25834;
  wire tmp25835;
  wire tmp25836;
  wire tmp25837;
  wire tmp25838;
  wire tmp25839;
  wire tmp25840;
  wire tmp25841;
  wire tmp25842;
  wire tmp25843;
  wire tmp25844;
  wire tmp25845;
  wire tmp25846;
  wire tmp25847;
  wire tmp25848;
  wire tmp25849;
  wire tmp25850;
  wire tmp25851;
  wire tmp25852;
  wire tmp25853;
  wire tmp25854;
  wire tmp25855;
  wire tmp25856;
  wire tmp25857;
  wire tmp25858;
  wire tmp25859;
  wire tmp25860;
  wire tmp25861;
  wire tmp25862;
  wire tmp25863;
  wire tmp25864;
  wire tmp25865;
  wire tmp25866;
  wire tmp25867;
  wire tmp25868;
  wire tmp25869;
  wire tmp25870;
  wire tmp25871;
  wire tmp25872;
  wire tmp25873;
  wire tmp25874;
  wire tmp25875;
  wire tmp25876;
  wire tmp25877;
  wire tmp25878;
  wire tmp25879;
  wire tmp25880;
  wire tmp25881;
  wire tmp25882;
  wire tmp25883;
  wire tmp25884;
  wire tmp25885;
  wire tmp25886;
  wire tmp25887;
  wire tmp25888;
  wire tmp25889;
  wire tmp25890;
  wire tmp25891;
  wire tmp25892;
  wire tmp25893;
  wire tmp25894;
  wire tmp25895;
  wire tmp25896;
  wire tmp25897;
  wire tmp25898;
  wire tmp25899;
  wire tmp25900;
  wire tmp25901;
  wire tmp25902;
  wire tmp25903;
  wire tmp25904;
  wire tmp25905;
  wire tmp25906;
  wire tmp25907;
  wire tmp25908;
  wire tmp25909;
  wire tmp25910;
  wire tmp25911;
  wire tmp25912;
  wire tmp25913;
  wire tmp25914;
  wire tmp25915;
  wire tmp25916;
  wire tmp25917;
  wire tmp25918;
  wire tmp25919;
  wire tmp25920;
  wire tmp25921;
  wire tmp25922;
  wire tmp25923;
  wire tmp25924;
  wire tmp25925;
  wire tmp25926;
  wire tmp25927;
  wire tmp25928;
  wire tmp25929;
  wire tmp25930;
  wire tmp25931;
  wire tmp25932;
  wire tmp25933;
  wire tmp25934;
  wire tmp25935;
  wire tmp25936;
  wire tmp25937;
  wire tmp25938;
  wire tmp25939;
  wire tmp25940;
  wire tmp25941;
  wire tmp25942;
  wire tmp25943;
  wire tmp25944;
  wire tmp25945;
  wire tmp25946;
  wire tmp25947;
  wire tmp25948;
  wire tmp25949;
  wire tmp25950;
  wire tmp25951;
  wire tmp25952;
  wire tmp25953;
  wire tmp25954;
  wire tmp25955;
  wire tmp25956;
  wire tmp25957;
  wire tmp25958;
  wire tmp25959;
  wire tmp25960;
  wire tmp25961;
  wire tmp25962;
  wire tmp25963;
  wire tmp25964;
  wire tmp25965;
  wire tmp25966;
  wire tmp25967;
  wire tmp25968;
  wire tmp25969;
  wire tmp25970;
  wire tmp25971;
  wire tmp25972;
  wire tmp25973;
  wire tmp25974;
  wire tmp25975;
  wire tmp25976;
  wire tmp25977;
  wire tmp25978;
  wire tmp25979;
  wire tmp25980;
  wire tmp25981;
  wire tmp25982;
  wire tmp25983;
  wire tmp25984;
  wire tmp25985;
  wire tmp25986;
  wire tmp25987;
  wire tmp25988;
  wire tmp25989;
  wire tmp25990;
  wire tmp25991;
  wire tmp25992;
  wire tmp25993;
  wire tmp25994;
  wire tmp25995;
  wire tmp25996;
  wire tmp25997;
  wire tmp25998;
  wire tmp25999;
  wire tmp26000;
  wire tmp26001;
  wire tmp26002;
  wire tmp26003;
  wire tmp26004;
  wire tmp26005;
  wire tmp26006;
  wire tmp26007;
  wire tmp26008;
  wire tmp26009;
  wire tmp26010;
  wire tmp26011;
  wire tmp26012;
  wire tmp26013;
  wire tmp26014;
  wire tmp26015;
  wire tmp26016;
  wire tmp26017;
  wire tmp26018;
  wire tmp26019;
  wire tmp26020;
  wire tmp26021;
  wire tmp26022;
  wire tmp26023;
  wire tmp26024;
  wire tmp26025;
  wire tmp26026;
  wire tmp26027;
  wire tmp26028;
  wire tmp26029;
  wire tmp26030;
  wire tmp26031;
  wire tmp26032;
  wire tmp26033;
  wire tmp26034;
  wire tmp26035;
  wire tmp26036;
  wire tmp26037;
  wire tmp26038;
  wire tmp26039;
  wire tmp26040;
  wire tmp26041;
  wire tmp26042;
  wire tmp26043;
  wire tmp26044;
  wire tmp26045;
  wire tmp26046;
  wire tmp26047;
  wire tmp26048;
  wire tmp26049;
  wire tmp26050;
  wire tmp26051;
  wire tmp26052;
  wire tmp26053;
  wire tmp26054;
  wire tmp26055;
  wire tmp26056;
  wire tmp26057;
  wire tmp26058;
  wire tmp26059;
  wire tmp26060;
  wire tmp26061;
  wire tmp26062;
  wire tmp26063;
  wire tmp26064;
  wire tmp26065;
  wire tmp26066;
  wire tmp26067;
  wire tmp26068;
  wire tmp26069;
  wire tmp26070;
  wire tmp26071;
  wire tmp26072;
  wire tmp26073;
  wire tmp26074;
  wire tmp26075;
  wire tmp26076;
  wire tmp26077;
  wire tmp26078;
  wire tmp26079;
  wire tmp26080;
  wire tmp26081;
  wire tmp26082;
  wire tmp26083;
  wire tmp26084;
  wire tmp26085;
  wire tmp26086;
  wire tmp26087;
  wire tmp26088;
  wire tmp26089;
  wire tmp26090;
  wire tmp26091;
  wire tmp26092;
  wire tmp26093;
  wire tmp26094;
  wire tmp26095;
  wire tmp26096;
  wire tmp26097;
  wire tmp26098;
  wire tmp26099;
  wire tmp26100;
  wire tmp26101;
  wire tmp26102;
  wire tmp26103;
  wire tmp26104;
  wire tmp26105;
  wire tmp26106;
  wire tmp26107;
  wire tmp26108;
  wire tmp26109;
  wire tmp26110;
  wire tmp26111;
  wire tmp26112;
  wire tmp26113;
  wire tmp26114;
  wire tmp26115;
  wire tmp26116;
  wire tmp26117;
  wire tmp26118;
  wire tmp26119;
  wire tmp26120;
  wire tmp26121;
  wire tmp26122;
  wire tmp26123;
  wire tmp26124;
  wire tmp26125;
  wire tmp26126;
  wire tmp26127;
  wire tmp26128;
  wire tmp26129;
  wire tmp26130;
  wire tmp26131;
  wire tmp26132;
  wire tmp26133;
  wire tmp26134;
  wire tmp26135;
  wire tmp26136;
  wire tmp26137;
  wire tmp26138;
  wire tmp26139;
  wire tmp26140;
  wire tmp26141;
  wire tmp26142;
  wire tmp26143;
  wire tmp26144;
  wire tmp26145;
  wire tmp26146;
  wire tmp26147;
  wire tmp26148;
  wire tmp26149;
  wire tmp26150;
  wire tmp26151;
  wire tmp26152;
  wire tmp26153;
  wire tmp26154;
  wire tmp26155;
  wire tmp26156;
  wire tmp26157;
  wire tmp26158;
  wire tmp26159;
  wire tmp26160;
  wire tmp26161;
  wire tmp26162;
  wire tmp26163;
  wire tmp26164;
  wire tmp26165;
  wire tmp26166;
  wire tmp26167;
  wire tmp26168;
  wire tmp26169;
  wire tmp26170;
  wire tmp26171;
  wire tmp26172;
  wire tmp26173;
  wire tmp26174;
  wire tmp26175;
  wire tmp26176;
  wire tmp26177;
  wire tmp26178;
  wire tmp26179;
  wire tmp26180;
  wire tmp26181;
  wire tmp26182;
  wire tmp26183;
  wire tmp26184;
  wire tmp26185;
  wire tmp26186;
  wire tmp26187;
  wire tmp26188;
  wire tmp26189;
  wire tmp26190;
  wire tmp26191;
  wire tmp26192;
  wire tmp26193;
  wire tmp26194;
  wire tmp26195;
  wire tmp26196;
  wire tmp26197;
  wire tmp26198;
  wire tmp26199;
  wire tmp26200;
  wire tmp26201;
  wire tmp26202;
  wire tmp26203;
  wire tmp26204;
  wire tmp26205;
  wire tmp26206;
  wire tmp26207;
  wire tmp26208;
  wire tmp26209;
  wire tmp26210;
  wire tmp26211;
  wire tmp26212;
  wire tmp26213;
  wire tmp26214;
  wire tmp26215;
  wire tmp26216;
  wire tmp26217;
  wire tmp26218;
  wire tmp26219;
  wire tmp26220;
  wire tmp26221;
  wire tmp26222;
  wire tmp26223;
  wire tmp26224;
  wire tmp26225;
  wire tmp26226;
  wire tmp26227;
  wire tmp26228;
  wire tmp26229;
  wire tmp26230;
  wire tmp26231;
  wire tmp26232;
  wire tmp26233;
  wire tmp26234;
  wire tmp26235;
  wire tmp26236;
  wire tmp26237;
  wire tmp26238;
  wire tmp26239;
  wire tmp26240;
  wire tmp26241;
  wire tmp26242;
  wire tmp26243;
  wire tmp26244;
  wire tmp26245;
  wire tmp26246;
  wire tmp26247;
  wire tmp26248;
  wire tmp26249;
  wire tmp26250;
  wire tmp26251;
  wire tmp26252;
  wire tmp26253;
  wire tmp26254;
  wire tmp26255;
  wire tmp26256;
  wire tmp26257;
  wire tmp26258;
  wire tmp26259;
  wire tmp26260;
  wire tmp26261;
  wire tmp26262;
  wire tmp26263;
  wire tmp26264;
  wire tmp26265;
  wire tmp26266;
  wire tmp26267;
  wire tmp26268;
  wire tmp26269;
  wire tmp26270;
  wire tmp26271;
  wire tmp26272;
  wire tmp26273;
  wire tmp26274;
  wire tmp26275;
  wire tmp26276;
  wire tmp26277;
  wire tmp26278;
  wire tmp26279;
  wire tmp26280;
  wire tmp26281;
  wire tmp26282;
  wire tmp26283;
  wire tmp26284;
  wire tmp26285;
  wire tmp26286;
  wire tmp26287;
  wire tmp26288;
  wire tmp26289;
  wire tmp26290;
  wire tmp26291;
  wire tmp26292;
  wire tmp26293;
  wire tmp26294;
  wire tmp26295;
  wire tmp26296;
  wire tmp26297;
  wire tmp26298;
  wire tmp26299;
  wire tmp26300;
  wire tmp26301;
  wire tmp26302;
  wire tmp26303;
  wire tmp26304;
  wire tmp26305;
  wire tmp26306;
  wire tmp26307;
  wire tmp26308;
  wire tmp26309;
  wire tmp26310;
  wire tmp26311;
  wire tmp26312;
  wire tmp26313;
  wire tmp26314;
  wire tmp26315;
  wire tmp26316;
  wire tmp26317;
  wire tmp26318;
  wire tmp26319;
  wire tmp26320;
  wire tmp26321;
  wire tmp26322;
  wire tmp26323;
  wire tmp26324;
  wire tmp26325;
  wire tmp26326;
  wire tmp26327;
  wire tmp26328;
  wire tmp26329;
  wire tmp26330;
  wire tmp26331;
  wire tmp26332;
  wire tmp26333;
  wire tmp26334;
  wire tmp26335;
  wire tmp26336;
  wire tmp26337;
  wire tmp26338;
  wire tmp26339;
  wire tmp26340;
  wire tmp26341;
  wire tmp26342;
  wire tmp26343;
  wire tmp26344;
  wire tmp26345;
  wire tmp26346;
  wire tmp26347;
  wire tmp26348;
  wire tmp26349;
  wire tmp26350;
  wire tmp26351;
  wire tmp26352;
  wire tmp26353;
  wire tmp26354;
  wire tmp26355;
  wire tmp26356;
  wire tmp26357;
  wire tmp26358;
  wire tmp26359;
  wire tmp26360;
  wire tmp26361;
  wire tmp26362;
  wire tmp26363;
  wire tmp26364;
  wire tmp26365;
  wire tmp26366;
  wire tmp26367;
  wire tmp26368;
  wire tmp26369;
  wire tmp26370;
  wire tmp26371;
  wire tmp26372;
  wire tmp26373;
  wire tmp26374;
  wire tmp26375;
  wire tmp26376;
  wire tmp26377;
  wire tmp26378;
  wire tmp26379;
  wire tmp26380;
  wire tmp26381;
  wire tmp26382;
  wire tmp26383;
  wire tmp26384;
  wire tmp26385;
  wire tmp26386;
  wire tmp26387;
  wire tmp26388;
  wire tmp26389;
  wire tmp26390;
  wire tmp26391;
  wire tmp26392;
  wire tmp26393;
  wire tmp26394;
  wire tmp26395;
  wire tmp26396;
  wire tmp26397;
  wire tmp26398;
  wire tmp26399;
  wire tmp26400;
  wire tmp26401;
  wire tmp26402;
  wire tmp26403;
  wire tmp26404;
  wire tmp26405;
  wire tmp26406;
  wire tmp26407;
  wire tmp26408;
  wire tmp26409;
  wire tmp26410;
  wire tmp26411;
  wire tmp26412;
  wire tmp26413;
  wire tmp26414;
  wire tmp26415;
  wire tmp26416;
  wire tmp26417;
  wire tmp26418;
  wire tmp26419;
  wire tmp26420;
  wire tmp26421;
  wire tmp26422;
  wire tmp26423;
  wire tmp26424;
  wire tmp26425;
  wire tmp26426;
  wire tmp26427;
  wire tmp26428;
  wire tmp26429;
  wire tmp26430;
  wire tmp26431;
  wire tmp26432;
  wire tmp26433;
  wire tmp26434;
  wire tmp26435;
  wire tmp26436;
  wire tmp26437;
  wire tmp26438;
  wire tmp26439;
  wire tmp26440;
  wire tmp26441;
  wire tmp26442;
  wire tmp26443;
  wire tmp26444;
  wire tmp26445;
  wire tmp26446;
  wire tmp26447;
  wire tmp26448;
  wire tmp26449;
  wire tmp26450;
  wire tmp26451;
  wire tmp26452;
  wire tmp26453;
  wire tmp26454;
  wire tmp26455;
  wire tmp26456;
  wire tmp26457;
  wire tmp26458;
  wire tmp26459;
  wire tmp26460;
  wire tmp26461;
  wire tmp26462;
  wire tmp26463;
  wire tmp26464;
  wire tmp26465;
  wire tmp26466;
  wire tmp26467;
  wire tmp26468;
  wire tmp26469;
  wire tmp26470;
  wire tmp26471;
  wire tmp26472;
  wire tmp26473;
  wire tmp26474;
  wire tmp26475;
  wire tmp26476;
  wire tmp26477;
  wire tmp26478;
  wire tmp26479;
  wire tmp26480;
  wire tmp26481;
  wire tmp26482;
  wire tmp26483;
  wire tmp26484;
  wire tmp26485;
  wire tmp26486;
  wire tmp26487;
  wire tmp26488;
  wire tmp26489;
  wire tmp26490;
  wire tmp26491;
  wire tmp26492;
  wire tmp26493;
  wire tmp26494;
  wire tmp26495;
  wire tmp26496;
  wire tmp26497;
  wire tmp26498;
  wire tmp26499;
  wire tmp26500;
  wire tmp26501;
  wire tmp26502;
  wire tmp26503;
  wire tmp26504;
  wire tmp26505;
  wire tmp26506;
  wire tmp26507;
  wire tmp26508;
  wire tmp26509;
  wire tmp26510;
  wire tmp26511;
  wire tmp26512;
  wire tmp26513;
  wire tmp26514;
  wire tmp26515;
  wire tmp26516;
  wire tmp26517;
  wire tmp26518;
  wire tmp26519;
  wire tmp26520;
  wire tmp26521;
  wire tmp26522;
  wire tmp26523;
  wire tmp26524;
  wire tmp26525;
  wire tmp26526;
  wire tmp26527;
  wire tmp26528;
  wire tmp26529;
  wire tmp26530;
  wire tmp26531;
  wire tmp26532;
  wire tmp26533;
  wire tmp26534;
  wire tmp26535;
  wire tmp26536;
  wire tmp26537;
  wire tmp26538;
  wire tmp26539;
  wire tmp26540;
  wire tmp26541;
  wire tmp26542;
  wire tmp26543;
  wire tmp26544;
  wire tmp26545;
  wire tmp26546;
  wire tmp26547;
  wire tmp26548;
  wire tmp26549;
  wire tmp26550;
  wire tmp26551;
  wire tmp26552;
  wire tmp26553;
  wire tmp26554;
  wire tmp26555;
  wire tmp26556;
  wire tmp26557;
  wire tmp26558;
  wire tmp26559;
  wire tmp26560;
  wire tmp26561;
  wire tmp26562;
  wire tmp26563;
  wire tmp26564;
  wire tmp26565;
  wire tmp26566;
  wire tmp26567;
  wire tmp26568;
  wire tmp26569;
  wire tmp26570;
  wire tmp26571;
  wire tmp26572;
  wire tmp26573;
  wire tmp26574;
  wire tmp26575;
  wire tmp26576;
  wire tmp26577;
  wire tmp26578;
  wire tmp26579;
  wire tmp26580;
  wire tmp26581;
  wire tmp26582;
  wire tmp26583;
  wire tmp26584;
  wire tmp26585;
  wire tmp26586;
  wire tmp26587;
  wire tmp26588;
  wire tmp26589;
  wire tmp26590;
  wire tmp26591;
  wire tmp26592;
  wire tmp26593;
  wire tmp26594;
  wire tmp26595;
  wire tmp26596;
  wire tmp26597;
  wire tmp26598;
  wire tmp26599;
  wire tmp26600;
  wire tmp26601;
  wire tmp26602;
  wire tmp26603;
  wire tmp26604;
  wire tmp26605;
  wire tmp26606;
  wire tmp26607;
  wire tmp26608;
  wire tmp26609;
  wire tmp26610;
  wire tmp26611;
  wire tmp26612;
  wire tmp26613;
  wire tmp26614;
  wire tmp26615;
  wire tmp26616;
  wire tmp26617;
  wire tmp26618;
  wire tmp26619;
  wire tmp26620;
  wire tmp26621;
  wire tmp26622;
  wire tmp26623;
  wire tmp26624;
  wire tmp26625;
  wire tmp26626;
  wire tmp26627;
  wire tmp26628;
  wire tmp26629;
  wire tmp26630;
  wire tmp26631;
  wire tmp26632;
  wire tmp26633;
  wire tmp26634;
  wire tmp26635;
  wire tmp26636;
  wire tmp26637;
  wire tmp26638;
  wire tmp26639;
  wire tmp26640;
  wire tmp26641;
  wire tmp26642;
  wire tmp26643;
  wire tmp26644;
  wire tmp26645;
  wire tmp26646;
  wire tmp26647;
  wire tmp26648;
  wire tmp26649;
  wire tmp26650;
  wire tmp26651;
  wire tmp26652;
  wire tmp26653;
  wire tmp26654;
  wire tmp26655;
  wire tmp26656;
  wire tmp26657;
  wire tmp26658;
  wire tmp26659;
  wire tmp26660;
  wire tmp26661;
  wire tmp26662;
  wire tmp26663;
  wire tmp26664;
  wire tmp26665;
  wire tmp26666;
  wire tmp26667;
  wire tmp26668;
  wire tmp26669;
  wire tmp26670;
  wire tmp26671;
  wire tmp26672;
  wire tmp26673;
  wire tmp26674;
  wire tmp26675;
  wire tmp26676;
  wire tmp26677;
  wire tmp26678;
  wire tmp26679;
  wire tmp26680;
  wire tmp26681;
  wire tmp26682;
  wire tmp26683;
  wire tmp26684;
  wire tmp26685;
  wire tmp26686;
  wire tmp26687;
  wire tmp26688;
  wire tmp26689;
  wire tmp26690;
  wire tmp26691;
  wire tmp26692;
  wire tmp26693;
  wire tmp26694;
  wire tmp26695;
  wire tmp26696;
  wire tmp26697;
  wire tmp26698;
  wire tmp26699;
  wire tmp26700;
  wire tmp26701;
  wire tmp26702;
  wire tmp26703;
  wire tmp26704;
  wire tmp26705;
  wire tmp26706;
  wire tmp26707;
  wire tmp26708;
  wire tmp26709;
  wire tmp26710;
  wire tmp26711;
  wire tmp26712;
  wire tmp26713;
  wire tmp26714;
  wire tmp26715;
  wire tmp26716;
  wire tmp26717;
  wire tmp26718;
  wire tmp26719;
  wire tmp26720;
  wire tmp26721;
  wire tmp26722;
  wire tmp26723;
  wire tmp26724;
  wire tmp26725;
  wire tmp26726;
  wire tmp26727;
  wire tmp26728;
  wire tmp26729;
  wire tmp26730;
  wire tmp26731;
  wire tmp26732;
  wire tmp26733;
  wire tmp26734;
  wire tmp26735;
  wire tmp26736;
  wire tmp26737;
  wire tmp26738;
  wire tmp26739;
  wire tmp26740;
  wire tmp26741;
  wire tmp26742;
  wire tmp26743;
  wire tmp26744;
  wire tmp26745;
  wire tmp26746;
  wire tmp26747;
  wire tmp26748;
  wire tmp26749;
  wire tmp26750;
  wire tmp26751;
  wire tmp26752;
  wire tmp26753;
  wire tmp26754;
  wire tmp26755;
  wire tmp26756;
  wire tmp26757;
  wire tmp26758;
  wire tmp26759;
  wire tmp26760;
  wire tmp26761;
  wire tmp26762;
  wire tmp26763;
  wire tmp26764;
  wire tmp26765;
  wire tmp26766;
  wire tmp26767;
  wire tmp26768;
  wire tmp26769;
  wire tmp26770;
  wire tmp26771;
  wire tmp26772;
  wire tmp26773;
  wire tmp26774;
  wire tmp26775;
  wire tmp26776;
  wire tmp26777;
  wire tmp26778;
  wire tmp26779;
  wire tmp26780;
  wire tmp26781;
  wire tmp26782;
  wire tmp26783;
  wire tmp26784;
  wire tmp26785;
  wire tmp26786;
  wire tmp26787;
  wire tmp26788;
  wire tmp26789;
  wire tmp26790;
  wire tmp26791;
  wire tmp26792;
  wire tmp26793;
  wire tmp26794;
  wire tmp26795;
  wire tmp26796;
  wire tmp26797;
  wire tmp26798;
  wire tmp26799;
  wire tmp26800;
  wire tmp26801;
  wire tmp26802;
  wire tmp26803;
  wire tmp26804;
  wire tmp26805;
  wire tmp26806;
  wire tmp26807;
  wire tmp26808;
  wire tmp26809;
  wire tmp26810;
  wire tmp26811;
  wire tmp26812;
  wire tmp26813;
  wire tmp26814;
  wire tmp26815;
  wire tmp26816;
  wire tmp26817;
  wire tmp26818;
  wire tmp26819;
  wire tmp26820;
  wire tmp26821;
  wire tmp26822;
  wire tmp26823;
  wire tmp26824;
  wire tmp26825;
  wire tmp26826;
  wire tmp26827;
  wire tmp26828;
  wire tmp26829;
  wire tmp26830;
  wire tmp26831;
  wire tmp26832;
  wire tmp26833;
  wire tmp26834;
  wire tmp26835;
  wire tmp26836;
  wire tmp26837;
  wire tmp26838;
  wire tmp26839;
  wire tmp26840;
  wire tmp26841;
  wire tmp26842;
  wire tmp26843;
  wire tmp26844;
  wire tmp26845;
  wire tmp26846;
  wire tmp26847;
  wire tmp26848;
  wire tmp26849;
  wire tmp26850;
  wire tmp26851;
  wire tmp26852;
  wire tmp26853;
  wire tmp26854;
  wire tmp26855;
  wire tmp26856;
  wire tmp26857;
  wire tmp26858;
  wire tmp26859;
  wire tmp26860;
  wire tmp26861;
  wire tmp26862;
  wire tmp26863;
  wire tmp26864;
  wire tmp26865;
  wire tmp26866;
  wire tmp26867;
  wire tmp26868;
  wire tmp26869;
  wire tmp26870;
  wire tmp26871;
  wire tmp26872;
  wire tmp26873;
  wire tmp26874;
  wire tmp26875;
  wire tmp26876;
  wire tmp26877;
  wire tmp26878;
  wire tmp26879;
  wire tmp26880;
  wire tmp26881;
  wire tmp26882;
  wire tmp26883;
  wire tmp26884;
  wire tmp26885;
  wire tmp26886;
  wire tmp26887;
  wire tmp26888;
  wire tmp26889;
  wire tmp26890;
  wire tmp26891;
  wire tmp26892;
  wire tmp26893;
  wire tmp26894;
  wire tmp26895;
  wire tmp26896;
  wire tmp26897;
  wire tmp26898;
  wire tmp26899;
  wire tmp26900;
  wire tmp26901;
  wire tmp26902;
  wire tmp26903;
  wire tmp26904;
  wire tmp26905;
  wire tmp26906;
  wire tmp26907;
  wire tmp26908;
  wire tmp26909;
  wire tmp26910;
  wire tmp26911;
  wire tmp26912;
  wire tmp26913;
  wire tmp26914;
  wire tmp26915;
  wire tmp26916;
  wire tmp26917;
  wire tmp26918;
  wire tmp26919;
  wire tmp26920;
  wire tmp26921;
  wire tmp26922;
  wire tmp26923;
  wire tmp26924;
  wire tmp26925;
  wire tmp26926;
  wire tmp26927;
  wire tmp26928;
  wire tmp26929;
  wire tmp26930;
  wire tmp26931;
  wire tmp26932;
  wire tmp26933;
  wire tmp26934;
  wire tmp26935;
  wire tmp26936;
  wire tmp26937;
  wire tmp26938;
  wire tmp26939;
  wire tmp26940;
  wire tmp26941;
  wire tmp26942;
  wire tmp26943;
  wire tmp26944;
  wire tmp26945;
  wire tmp26946;
  wire tmp26947;
  wire tmp26948;
  wire tmp26949;
  wire tmp26950;
  wire tmp26951;
  wire tmp26952;
  wire tmp26953;
  wire tmp26954;
  wire tmp26955;
  wire tmp26956;
  wire tmp26957;
  wire tmp26958;
  wire tmp26959;
  wire tmp26960;
  wire tmp26961;
  wire tmp26962;
  wire tmp26963;
  wire tmp26964;
  wire tmp26965;
  wire tmp26966;
  wire tmp26967;
  wire tmp26968;
  wire tmp26969;
  wire tmp26970;
  wire tmp26971;
  wire tmp26972;
  wire tmp26973;
  wire tmp26974;
  wire tmp26975;
  wire tmp26976;
  wire tmp26977;
  wire tmp26978;
  wire tmp26979;
  wire tmp26980;
  wire tmp26981;
  wire tmp26982;
  wire tmp26983;
  wire tmp26984;
  wire tmp26985;
  wire tmp26986;
  wire tmp26987;
  wire tmp26988;
  wire tmp26989;
  wire tmp26990;
  wire tmp26991;
  wire tmp26992;
  wire tmp26993;
  wire tmp26994;
  wire tmp26995;
  wire tmp26996;
  wire tmp26997;
  wire tmp26998;
  wire tmp26999;
  wire tmp27000;
  wire tmp27001;
  wire tmp27002;
  wire tmp27003;
  wire tmp27004;
  wire tmp27005;
  wire tmp27006;
  wire tmp27007;
  wire tmp27008;
  wire tmp27009;
  wire tmp27010;
  wire tmp27011;
  wire tmp27012;
  wire tmp27013;
  wire tmp27014;
  wire tmp27015;
  wire tmp27016;
  wire tmp27017;
  wire tmp27018;
  wire tmp27019;
  wire tmp27020;
  wire tmp27021;
  wire tmp27022;
  wire tmp27023;
  wire tmp27024;
  wire tmp27025;
  wire tmp27026;
  wire tmp27027;
  wire tmp27028;
  wire tmp27029;
  wire tmp27030;
  wire tmp27031;
  wire tmp27032;
  wire tmp27033;
  wire tmp27034;
  wire tmp27035;
  wire tmp27036;
  wire tmp27037;
  wire tmp27038;
  wire tmp27039;
  wire tmp27040;
  wire tmp27041;
  wire tmp27042;
  wire tmp27043;
  wire tmp27044;
  wire tmp27045;
  wire tmp27046;
  wire tmp27047;
  wire tmp27048;
  wire tmp27049;
  wire tmp27050;
  wire tmp27051;
  wire tmp27052;
  wire tmp27053;
  wire tmp27054;
  wire tmp27055;
  wire tmp27056;
  wire tmp27057;
  wire tmp27058;
  wire tmp27059;
  wire tmp27060;
  wire tmp27061;
  wire tmp27062;
  wire tmp27063;
  wire tmp27064;
  wire tmp27065;
  wire tmp27066;
  wire tmp27067;
  wire tmp27068;
  wire tmp27069;
  wire tmp27070;
  wire tmp27071;
  wire tmp27072;
  wire tmp27073;
  wire tmp27074;
  wire tmp27075;
  wire tmp27076;
  wire tmp27077;
  wire tmp27078;
  wire tmp27079;
  wire tmp27080;
  wire tmp27081;
  wire tmp27082;
  wire tmp27083;
  wire tmp27084;
  wire tmp27085;
  wire tmp27086;
  wire tmp27087;
  wire tmp27088;
  wire tmp27089;
  wire tmp27090;
  wire tmp27091;
  wire tmp27092;
  wire tmp27093;
  wire tmp27094;
  wire tmp27095;
  wire tmp27096;
  wire tmp27097;
  wire tmp27098;
  wire tmp27099;
  wire tmp27100;
  wire tmp27101;
  wire tmp27102;
  wire tmp27103;
  wire tmp27104;
  wire tmp27105;
  wire tmp27106;
  wire tmp27107;
  wire tmp27108;
  wire tmp27109;
  wire tmp27110;
  wire tmp27111;
  wire tmp27112;
  wire tmp27113;
  wire tmp27114;
  wire tmp27115;
  wire tmp27116;
  wire tmp27117;
  wire tmp27118;
  wire tmp27119;
  wire tmp27120;
  wire tmp27121;
  wire tmp27122;
  wire tmp27123;
  wire tmp27124;
  wire tmp27125;
  wire tmp27126;
  wire tmp27127;
  wire tmp27128;
  wire tmp27129;
  wire tmp27130;
  wire tmp27131;
  wire tmp27132;
  wire tmp27133;
  wire tmp27134;
  wire tmp27135;
  wire tmp27136;
  wire tmp27137;
  wire tmp27138;
  wire tmp27139;
  wire tmp27140;
  wire tmp27141;
  wire tmp27142;
  wire tmp27143;
  wire tmp27144;
  wire tmp27145;
  wire tmp27146;
  wire tmp27147;
  wire tmp27148;
  wire tmp27149;
  wire tmp27150;
  wire tmp27151;
  wire tmp27152;
  wire tmp27153;
  wire tmp27154;
  wire tmp27155;
  wire tmp27156;
  wire tmp27157;
  wire tmp27158;
  wire tmp27159;
  wire tmp27160;
  wire tmp27161;
  wire tmp27162;
  wire tmp27163;
  wire tmp27164;
  wire tmp27165;
  wire tmp27166;
  wire tmp27167;
  wire tmp27168;
  wire tmp27169;
  wire tmp27170;
  wire tmp27171;
  wire tmp27172;
  wire tmp27173;
  wire tmp27174;
  wire tmp27175;
  wire tmp27176;
  wire tmp27177;
  wire tmp27178;
  wire tmp27179;
  wire tmp27180;
  wire tmp27181;
  wire tmp27182;
  wire tmp27183;
  wire tmp27184;
  wire tmp27185;
  wire tmp27186;
  wire tmp27187;
  wire tmp27188;
  wire tmp27189;
  wire tmp27190;
  wire tmp27191;
  wire tmp27192;
  wire tmp27193;
  wire tmp27194;
  wire tmp27195;
  wire tmp27196;
  wire tmp27197;
  wire tmp27198;
  wire tmp27199;
  wire tmp27200;
  wire tmp27201;
  wire tmp27202;
  wire tmp27203;
  wire tmp27204;
  wire tmp27205;
  wire tmp27206;
  wire tmp27207;
  wire tmp27208;
  wire tmp27209;
  wire tmp27210;
  wire tmp27211;
  wire tmp27212;
  wire tmp27213;
  wire tmp27214;
  wire tmp27215;
  wire tmp27216;
  wire tmp27217;
  wire tmp27218;
  wire tmp27219;
  wire tmp27220;
  wire tmp27221;
  wire tmp27222;
  wire tmp27223;
  wire tmp27224;
  wire tmp27225;
  wire tmp27226;
  wire tmp27227;
  wire tmp27228;
  wire tmp27229;
  wire tmp27230;
  wire tmp27231;
  wire tmp27232;
  wire tmp27233;
  wire tmp27234;
  wire tmp27235;
  wire tmp27236;
  wire tmp27237;
  wire tmp27238;
  wire tmp27239;
  wire tmp27240;
  wire tmp27241;
  wire tmp27242;
  wire tmp27243;
  wire tmp27244;
  wire tmp27245;
  wire tmp27246;
  wire tmp27247;
  wire tmp27248;
  wire tmp27249;
  wire tmp27250;
  wire tmp27251;
  wire tmp27252;
  wire tmp27253;
  wire tmp27254;
  wire tmp27255;
  wire tmp27256;
  wire tmp27257;
  wire tmp27258;
  wire tmp27259;
  wire tmp27260;
  wire tmp27261;
  wire tmp27262;
  wire tmp27263;
  wire tmp27264;
  wire tmp27265;
  wire tmp27266;
  wire tmp27267;
  wire tmp27268;
  wire tmp27269;
  wire tmp27270;
  wire tmp27271;
  wire tmp27272;
  wire tmp27273;
  wire tmp27274;
  wire tmp27275;
  wire tmp27276;
  wire tmp27277;
  wire tmp27278;
  wire tmp27279;
  wire tmp27280;
  wire tmp27281;
  wire tmp27282;
  wire tmp27283;
  wire tmp27284;
  wire tmp27285;
  wire tmp27286;
  wire tmp27287;
  wire tmp27288;
  wire tmp27289;
  wire tmp27290;
  wire tmp27291;
  wire tmp27292;
  wire tmp27293;
  wire tmp27294;
  wire tmp27295;
  wire tmp27296;
  wire tmp27297;
  wire tmp27298;
  wire tmp27299;
  wire tmp27300;
  wire tmp27301;
  wire tmp27302;
  wire tmp27303;
  wire tmp27304;
  wire tmp27305;
  wire tmp27306;
  wire tmp27307;
  wire tmp27308;
  wire tmp27309;
  wire tmp27310;
  wire tmp27311;
  wire tmp27312;
  wire tmp27313;
  wire tmp27314;
  wire tmp27315;
  wire tmp27316;
  wire tmp27317;
  wire tmp27318;
  wire tmp27319;
  wire tmp27320;
  wire tmp27321;
  wire tmp27322;
  wire tmp27323;
  wire tmp27324;
  wire tmp27325;
  wire tmp27326;
  wire tmp27327;
  wire tmp27328;
  wire tmp27329;
  wire tmp27330;
  wire tmp27331;
  wire tmp27332;
  wire tmp27333;
  wire tmp27334;
  wire tmp27335;
  wire tmp27336;
  wire tmp27337;
  wire tmp27338;
  wire tmp27339;
  wire tmp27340;
  wire tmp27341;
  wire tmp27342;
  wire tmp27343;
  wire tmp27344;
  wire tmp27345;
  wire tmp27346;
  wire tmp27347;
  wire tmp27348;
  wire tmp27349;
  wire tmp27350;
  wire tmp27351;
  wire tmp27352;
  wire tmp27353;
  wire tmp27354;
  wire tmp27355;
  wire tmp27356;
  wire tmp27357;
  wire tmp27358;
  wire tmp27359;
  wire tmp27360;
  wire tmp27361;
  wire tmp27362;
  wire tmp27363;
  wire tmp27364;
  wire tmp27365;
  wire tmp27366;
  wire tmp27367;
  wire tmp27368;
  wire tmp27369;
  wire tmp27370;
  wire tmp27371;
  wire tmp27372;
  wire tmp27373;
  wire tmp27374;
  wire tmp27375;
  wire tmp27376;
  wire tmp27377;
  wire tmp27378;
  wire tmp27379;
  wire tmp27380;
  wire tmp27381;
  wire tmp27382;
  wire tmp27383;
  wire tmp27384;
  wire tmp27385;
  wire tmp27386;
  wire tmp27387;
  wire tmp27388;
  wire tmp27389;
  wire tmp27390;
  wire tmp27391;
  wire tmp27392;
  wire tmp27393;
  wire tmp27394;
  wire tmp27395;
  wire tmp27396;
  wire tmp27397;
  wire tmp27398;
  wire tmp27399;
  wire tmp27400;
  wire tmp27401;
  wire tmp27402;
  wire tmp27403;
  wire tmp27404;
  wire tmp27405;
  wire tmp27406;
  wire tmp27407;
  wire tmp27408;
  wire tmp27409;
  wire tmp27410;
  wire tmp27411;
  wire tmp27412;
  wire tmp27413;
  wire tmp27414;
  wire tmp27415;
  wire tmp27416;
  wire tmp27417;
  wire tmp27418;
  wire tmp27419;
  wire tmp27420;
  wire tmp27421;
  wire tmp27422;
  wire tmp27423;
  wire tmp27424;
  wire tmp27425;
  wire tmp27426;
  wire tmp27427;
  wire tmp27428;
  wire tmp27429;
  wire tmp27430;
  wire tmp27431;
  wire tmp27432;
  wire tmp27433;
  wire tmp27434;
  wire tmp27435;
  wire tmp27436;
  wire tmp27437;
  wire tmp27438;
  wire tmp27439;
  wire tmp27440;
  wire tmp27441;
  wire tmp27442;
  wire tmp27443;
  wire tmp27444;
  wire tmp27445;
  wire tmp27446;
  wire tmp27447;
  wire tmp27448;
  wire tmp27449;
  wire tmp27450;
  wire tmp27451;
  wire tmp27452;
  wire tmp27453;
  wire tmp27454;
  wire tmp27455;
  wire tmp27456;
  wire tmp27457;
  wire tmp27458;
  wire tmp27459;
  wire tmp27460;
  wire tmp27461;
  wire tmp27462;
  wire tmp27463;
  wire tmp27464;
  wire tmp27465;
  wire tmp27466;
  wire tmp27467;
  wire tmp27468;
  wire tmp27469;
  wire tmp27470;
  wire tmp27471;
  wire tmp27472;
  wire tmp27473;
  wire tmp27474;
  wire tmp27475;
  wire tmp27476;
  wire tmp27477;
  wire tmp27478;
  wire tmp27479;
  wire tmp27480;
  wire tmp27481;
  wire tmp27482;
  wire tmp27483;
  wire tmp27484;
  wire tmp27485;
  wire tmp27486;
  wire tmp27487;
  wire tmp27488;
  wire tmp27489;
  wire tmp27490;
  wire tmp27491;
  wire tmp27492;
  wire tmp27493;
  wire tmp27494;
  wire tmp27495;
  wire tmp27496;
  wire tmp27497;
  wire tmp27498;
  wire tmp27499;
  wire tmp27500;
  wire tmp27501;
  wire tmp27502;
  wire tmp27503;
  wire tmp27504;
  wire tmp27505;
  wire tmp27506;
  wire tmp27507;
  wire tmp27508;
  wire tmp27509;
  wire tmp27510;
  wire tmp27511;
  wire tmp27512;
  wire tmp27513;
  wire tmp27514;
  wire tmp27515;
  wire tmp27516;
  wire tmp27517;
  wire tmp27518;
  wire tmp27519;
  wire tmp27520;
  wire tmp27521;
  wire tmp27522;
  wire tmp27523;
  wire tmp27524;
  wire tmp27525;
  wire tmp27526;
  wire tmp27527;
  wire tmp27528;
  wire tmp27529;
  wire tmp27530;
  wire tmp27531;
  wire tmp27532;
  wire tmp27533;
  wire tmp27534;
  wire tmp27535;
  wire tmp27536;
  wire tmp27537;
  wire tmp27538;
  wire tmp27539;
  wire tmp27540;
  wire tmp27541;
  wire tmp27542;
  wire tmp27543;
  wire tmp27544;
  wire tmp27545;
  wire tmp27546;
  wire tmp27547;
  wire tmp27548;
  wire tmp27549;
  wire tmp27550;
  wire tmp27551;
  wire tmp27552;
  wire tmp27553;
  wire tmp27554;
  wire tmp27555;
  wire tmp27556;
  wire tmp27557;
  wire tmp27558;
  wire tmp27559;
  wire tmp27560;
  wire tmp27561;
  wire tmp27562;
  wire tmp27563;
  wire tmp27564;
  wire tmp27565;
  wire tmp27566;
  wire tmp27567;
  wire tmp27568;
  wire tmp27569;
  wire tmp27570;
  wire tmp27571;
  wire tmp27572;
  wire tmp27573;
  wire tmp27574;
  wire tmp27575;
  wire tmp27576;
  wire tmp27577;
  wire tmp27578;
  wire tmp27579;
  wire tmp27580;
  wire tmp27581;
  wire tmp27582;
  wire tmp27583;
  wire tmp27584;
  wire tmp27585;
  wire tmp27586;
  wire tmp27587;
  wire tmp27588;
  wire tmp27589;
  wire tmp27590;
  wire tmp27591;
  wire tmp27592;
  wire tmp27593;
  wire tmp27594;
  wire tmp27595;
  wire tmp27596;
  wire tmp27597;
  wire tmp27598;
  wire tmp27599;
  wire tmp27600;
  wire tmp27601;
  wire tmp27602;
  wire tmp27603;
  wire tmp27604;
  wire tmp27605;
  wire tmp27606;
  wire tmp27607;
  wire tmp27608;
  wire tmp27609;
  wire tmp27610;
  wire tmp27611;
  wire tmp27612;
  wire tmp27613;
  wire tmp27614;
  wire tmp27615;
  wire tmp27616;
  wire tmp27617;
  wire tmp27618;
  wire tmp27619;
  wire tmp27620;
  wire tmp27621;
  wire tmp27622;
  wire tmp27623;
  wire tmp27624;
  wire tmp27625;
  wire tmp27626;
  wire tmp27627;
  wire tmp27628;
  wire tmp27629;
  wire tmp27630;
  wire tmp27631;
  wire tmp27632;
  wire tmp27633;
  wire tmp27634;
  wire tmp27635;
  wire tmp27636;
  wire tmp27637;
  wire tmp27638;
  wire tmp27639;
  wire tmp27640;
  wire tmp27641;
  wire tmp27642;
  wire tmp27643;
  wire tmp27644;
  wire tmp27645;
  wire tmp27646;
  wire tmp27647;
  wire tmp27648;
  wire tmp27649;
  wire tmp27650;
  wire tmp27651;
  wire tmp27652;
  wire tmp27653;
  wire tmp27654;
  wire tmp27655;
  wire tmp27656;
  wire tmp27657;
  wire tmp27658;
  wire tmp27659;
  wire tmp27660;
  wire tmp27661;
  wire tmp27662;
  wire tmp27663;
  wire tmp27664;
  wire tmp27665;
  wire tmp27666;
  wire tmp27667;
  wire tmp27668;
  wire tmp27669;
  wire tmp27670;
  wire tmp27671;
  wire tmp27672;
  wire tmp27673;
  wire tmp27674;
  wire tmp27675;
  wire tmp27676;
  wire tmp27677;
  wire tmp27678;
  wire tmp27679;
  wire tmp27680;
  wire tmp27681;
  wire tmp27682;
  wire tmp27683;
  wire tmp27684;
  wire tmp27685;
  wire tmp27686;
  wire tmp27687;
  wire tmp27688;
  wire tmp27689;
  wire tmp27690;
  wire tmp27691;
  wire tmp27692;
  wire tmp27693;
  wire tmp27694;
  wire tmp27695;
  wire tmp27696;
  wire tmp27697;
  wire tmp27698;
  wire tmp27699;
  wire tmp27700;
  wire tmp27701;
  wire tmp27702;
  wire tmp27703;
  wire tmp27704;
  wire tmp27705;
  wire tmp27706;
  wire tmp27707;
  wire tmp27708;
  wire tmp27709;
  wire tmp27710;
  wire tmp27711;
  wire tmp27712;
  wire tmp27713;
  wire tmp27714;
  wire tmp27715;
  wire tmp27716;
  wire tmp27717;
  wire tmp27718;
  wire tmp27719;
  wire tmp27720;
  wire tmp27721;
  wire tmp27722;
  wire tmp27723;
  wire tmp27724;
  wire tmp27725;
  wire tmp27726;
  wire tmp27727;
  wire tmp27728;
  wire tmp27729;
  wire tmp27730;
  wire tmp27731;
  wire tmp27732;
  wire tmp27733;
  wire tmp27734;
  wire tmp27735;
  wire tmp27736;
  wire tmp27737;
  wire tmp27738;
  wire tmp27739;
  wire tmp27740;
  wire tmp27741;
  wire tmp27742;
  wire tmp27743;
  wire tmp27744;
  wire tmp27745;
  wire tmp27746;
  wire tmp27747;
  wire tmp27748;
  wire tmp27749;
  wire tmp27750;
  wire tmp27751;
  wire tmp27752;
  wire tmp27753;
  wire tmp27754;
  wire tmp27755;
  wire tmp27756;
  wire tmp27757;
  wire tmp27758;
  wire tmp27759;
  wire tmp27760;
  wire tmp27761;
  wire tmp27762;
  wire tmp27763;
  wire tmp27764;
  wire tmp27765;
  wire tmp27766;
  wire tmp27767;
  wire tmp27768;
  wire tmp27769;
  wire tmp27770;
  wire tmp27771;
  wire tmp27772;
  wire tmp27773;
  wire tmp27774;
  wire tmp27775;
  wire tmp27776;
  wire tmp27777;
  wire tmp27778;
  wire tmp27779;
  wire tmp27780;
  wire tmp27781;
  wire tmp27782;
  wire tmp27783;
  wire tmp27784;
  wire tmp27785;
  wire tmp27786;
  wire tmp27787;
  wire tmp27788;
  wire tmp27789;
  wire tmp27790;
  wire tmp27791;
  wire tmp27792;
  wire tmp27793;
  wire tmp27794;
  wire tmp27795;
  wire tmp27796;
  wire tmp27797;
  wire tmp27798;
  wire tmp27799;
  wire tmp27800;
  wire tmp27801;
  wire tmp27802;
  wire tmp27803;
  wire tmp27804;
  wire tmp27805;
  wire tmp27806;
  wire tmp27807;
  wire tmp27808;
  wire tmp27809;
  wire tmp27810;
  wire tmp27811;
  wire tmp27812;
  wire tmp27813;
  wire tmp27814;
  wire tmp27815;
  wire tmp27816;
  wire tmp27817;
  wire tmp27818;
  wire tmp27819;
  wire tmp27820;
  wire tmp27821;
  wire tmp27822;
  wire tmp27823;
  wire tmp27824;
  wire tmp27825;
  wire tmp27826;
  wire tmp27827;
  wire tmp27828;
  wire tmp27829;
  wire tmp27830;
  wire tmp27831;
  wire tmp27832;
  wire tmp27833;
  wire tmp27834;
  wire tmp27835;
  wire tmp27836;
  wire tmp27837;
  wire tmp27838;
  wire tmp27839;
  wire tmp27840;
  wire tmp27841;
  wire tmp27842;
  wire tmp27843;
  wire tmp27844;
  wire tmp27845;
  wire tmp27846;
  wire tmp27847;
  wire tmp27848;
  wire tmp27849;
  wire tmp27850;
  wire tmp27851;
  wire tmp27852;
  wire tmp27853;
  wire tmp27854;
  wire tmp27855;
  wire tmp27856;
  wire tmp27857;
  wire tmp27858;
  wire tmp27859;
  wire tmp27860;
  wire tmp27861;
  wire tmp27862;
  wire tmp27863;
  wire tmp27864;
  wire tmp27865;
  wire tmp27866;
  wire tmp27867;
  wire tmp27868;
  wire tmp27869;
  wire tmp27870;
  wire tmp27871;
  wire tmp27872;
  wire tmp27873;
  wire tmp27874;
  wire tmp27875;
  wire tmp27876;
  wire tmp27877;
  wire tmp27878;
  wire tmp27879;
  wire tmp27880;
  wire tmp27881;
  wire tmp27882;
  wire tmp27883;
  wire tmp27884;
  wire tmp27885;
  wire tmp27886;
  wire tmp27887;
  wire tmp27888;
  wire tmp27889;
  wire tmp27890;
  wire tmp27891;
  wire tmp27892;
  wire tmp27893;
  wire tmp27894;
  wire tmp27895;
  wire tmp27896;
  wire tmp27897;
  wire tmp27898;
  wire tmp27899;
  wire tmp27900;
  wire tmp27901;
  wire tmp27902;
  wire tmp27903;
  wire tmp27904;
  wire tmp27905;
  wire tmp27906;
  wire tmp27907;
  wire tmp27908;
  wire tmp27909;
  wire tmp27910;
  wire tmp27911;
  wire tmp27912;
  wire tmp27913;
  wire tmp27914;
  wire tmp27915;
  wire tmp27916;
  wire tmp27917;
  wire tmp27918;
  wire tmp27919;
  wire tmp27920;
  wire tmp27921;
  wire tmp27922;
  wire tmp27923;
  wire tmp27924;
  wire tmp27925;
  wire tmp27926;
  wire tmp27927;
  wire tmp27928;
  wire tmp27929;
  wire tmp27930;
  wire tmp27931;
  wire tmp27932;
  wire tmp27933;
  wire tmp27934;
  wire tmp27935;
  wire tmp27936;
  wire tmp27937;
  wire tmp27938;
  wire tmp27939;
  wire tmp27940;
  wire tmp27941;
  wire tmp27942;
  wire tmp27943;
  wire tmp27944;
  wire tmp27945;
  wire tmp27946;
  wire tmp27947;
  wire tmp27948;
  wire tmp27949;
  wire tmp27950;
  wire tmp27951;
  wire tmp27952;
  wire tmp27953;
  wire tmp27954;
  wire tmp27955;
  wire tmp27956;
  wire tmp27957;
  wire tmp27958;
  wire tmp27959;
  wire tmp27960;
  wire tmp27961;
  wire tmp27962;
  wire tmp27963;
  wire tmp27964;
  wire tmp27965;
  wire tmp27966;
  wire tmp27967;
  wire tmp27968;
  wire tmp27969;
  wire tmp27970;
  wire tmp27971;
  wire tmp27972;
  wire tmp27973;
  wire tmp27974;
  wire tmp27975;
  wire tmp27976;
  wire tmp27977;
  wire tmp27978;
  wire tmp27979;
  wire tmp27980;
  wire tmp27981;
  wire tmp27982;
  wire tmp27983;
  wire tmp27984;
  wire tmp27985;
  wire tmp27986;
  wire tmp27987;
  wire tmp27988;
  wire tmp27989;
  wire tmp27990;
  wire tmp27991;
  wire tmp27992;
  wire tmp27993;
  wire tmp27994;
  wire tmp27995;
  wire tmp27996;
  wire tmp27997;
  wire tmp27998;
  wire tmp27999;
  wire tmp28000;
  wire tmp28001;
  wire tmp28002;
  wire tmp28003;
  wire tmp28004;
  wire tmp28005;
  wire tmp28006;
  wire tmp28007;
  wire tmp28008;
  wire tmp28009;
  wire tmp28010;
  wire tmp28011;
  wire tmp28012;
  wire tmp28013;
  wire tmp28014;
  wire tmp28015;
  wire tmp28016;
  wire tmp28017;
  wire tmp28018;
  wire tmp28019;
  wire tmp28020;
  wire tmp28021;
  wire tmp28022;
  wire tmp28023;
  wire tmp28024;
  wire tmp28025;
  wire tmp28026;
  wire tmp28027;
  wire tmp28028;
  wire tmp28029;
  wire tmp28030;
  wire tmp28031;
  wire tmp28032;
  wire tmp28033;
  wire tmp28034;
  wire tmp28035;
  wire tmp28036;
  wire tmp28037;
  wire tmp28038;
  wire tmp28039;
  wire tmp28040;
  wire tmp28041;
  wire tmp28042;
  wire tmp28043;
  wire tmp28044;
  wire tmp28045;
  wire tmp28046;
  wire tmp28047;
  wire tmp28048;
  wire tmp28049;
  wire tmp28050;
  wire tmp28051;
  wire tmp28052;
  wire tmp28053;
  wire tmp28054;
  wire tmp28055;
  wire tmp28056;
  wire tmp28057;
  wire tmp28058;
  wire tmp28059;
  wire tmp28060;
  wire tmp28061;
  wire tmp28062;
  wire tmp28063;
  wire tmp28064;
  wire tmp28065;
  wire tmp28066;
  wire tmp28067;
  wire tmp28068;
  wire tmp28069;
  wire tmp28070;
  wire tmp28071;
  wire tmp28072;
  wire tmp28073;
  wire tmp28074;
  wire tmp28075;
  wire tmp28076;
  wire tmp28077;
  wire tmp28078;
  wire tmp28079;
  wire tmp28080;
  wire tmp28081;
  wire tmp28082;
  wire tmp28083;
  wire tmp28084;
  wire tmp28085;
  wire tmp28086;
  wire tmp28087;
  wire tmp28088;
  wire tmp28089;
  wire tmp28090;
  wire tmp28091;
  wire tmp28092;
  wire tmp28093;
  wire tmp28094;
  wire tmp28095;
  wire tmp28096;
  wire tmp28097;
  wire tmp28098;
  wire tmp28099;
  wire tmp28100;
  wire tmp28101;
  wire tmp28102;
  wire tmp28103;
  wire tmp28104;
  wire tmp28105;
  wire tmp28106;
  wire tmp28107;
  wire tmp28108;
  wire tmp28109;
  wire tmp28110;
  wire tmp28111;
  wire tmp28112;
  wire tmp28113;
  wire tmp28114;
  wire tmp28115;
  wire tmp28116;
  wire tmp28117;
  wire tmp28118;
  wire tmp28119;
  wire tmp28120;
  wire tmp28121;
  wire tmp28122;
  wire tmp28123;
  wire tmp28124;
  wire tmp28125;
  wire tmp28126;
  wire tmp28127;
  wire tmp28128;
  wire tmp28129;
  wire tmp28130;
  wire tmp28131;
  wire tmp28132;
  wire tmp28133;
  wire tmp28134;
  wire tmp28135;
  wire tmp28136;
  wire tmp28137;
  wire tmp28138;
  wire tmp28139;
  wire tmp28140;
  wire tmp28141;
  wire tmp28142;
  wire tmp28143;
  wire tmp28144;
  wire tmp28145;
  wire tmp28146;
  wire tmp28147;
  wire tmp28148;
  wire tmp28149;
  wire tmp28150;
  wire tmp28151;
  wire tmp28152;
  wire tmp28153;
  wire tmp28154;
  wire tmp28155;
  wire tmp28156;
  wire tmp28157;
  wire tmp28158;
  wire tmp28159;
  wire tmp28160;
  wire tmp28161;
  wire tmp28162;
  wire tmp28163;
  wire tmp28164;
  wire tmp28165;
  wire tmp28166;
  wire tmp28167;
  wire tmp28168;
  wire tmp28169;
  wire tmp28170;
  wire tmp28171;
  wire tmp28172;
  wire tmp28173;
  wire tmp28174;
  wire tmp28175;
  wire tmp28176;
  wire tmp28177;
  wire tmp28178;
  wire tmp28179;
  wire tmp28180;
  wire tmp28181;
  wire tmp28182;
  wire tmp28183;
  wire tmp28184;
  wire tmp28185;
  wire tmp28186;
  wire tmp28187;
  wire tmp28188;
  wire tmp28189;
  wire tmp28190;
  wire tmp28191;
  wire tmp28192;
  wire tmp28193;
  wire tmp28194;
  wire tmp28195;
  wire tmp28196;
  wire tmp28197;
  wire tmp28198;
  wire tmp28199;
  wire tmp28200;
  wire tmp28201;
  wire tmp28202;
  wire tmp28203;
  wire tmp28204;
  wire tmp28205;
  wire tmp28206;
  wire tmp28207;
  wire tmp28208;
  wire tmp28209;
  wire tmp28210;
  wire tmp28211;
  wire tmp28212;
  wire tmp28213;
  wire tmp28214;
  wire tmp28215;
  wire tmp28216;
  wire tmp28217;
  wire tmp28218;
  wire tmp28219;
  wire tmp28220;
  wire tmp28221;
  wire tmp28222;
  wire tmp28223;
  wire tmp28224;
  wire tmp28225;
  wire tmp28226;
  wire tmp28227;
  wire tmp28228;
  wire tmp28229;
  wire tmp28230;
  wire tmp28231;
  wire tmp28232;
  wire tmp28233;
  wire tmp28234;
  wire tmp28235;
  wire tmp28236;
  wire tmp28237;
  wire tmp28238;
  wire tmp28239;
  wire tmp28240;
  wire tmp28241;
  wire tmp28242;
  wire tmp28243;
  wire tmp28244;
  wire tmp28245;
  wire tmp28246;
  wire tmp28247;
  wire tmp28248;
  wire tmp28249;
  wire tmp28250;
  wire tmp28251;
  wire tmp28252;
  wire tmp28253;
  wire tmp28254;
  wire tmp28255;
  wire tmp28256;
  wire tmp28257;
  wire tmp28258;
  wire tmp28259;
  wire tmp28260;
  wire tmp28261;
  wire tmp28262;
  wire tmp28263;
  wire tmp28264;
  wire tmp28265;
  wire tmp28266;
  wire tmp28267;
  wire tmp28268;
  wire tmp28269;
  wire tmp28270;
  wire tmp28271;
  wire tmp28272;
  wire tmp28273;
  wire tmp28274;
  wire tmp28275;
  wire tmp28276;
  wire tmp28277;
  wire tmp28278;
  wire tmp28279;
  wire tmp28280;
  wire tmp28281;
  wire tmp28282;
  wire tmp28283;
  wire tmp28284;
  wire tmp28285;
  wire tmp28286;
  wire tmp28287;
  wire tmp28288;
  wire tmp28289;
  wire tmp28290;
  wire tmp28291;
  wire tmp28292;
  wire tmp28293;
  wire tmp28294;
  wire tmp28295;
  wire tmp28296;
  wire tmp28297;
  wire tmp28298;
  wire tmp28299;
  wire tmp28300;
  wire tmp28301;
  wire tmp28302;
  wire tmp28303;
  wire tmp28304;
  wire tmp28305;
  wire tmp28306;
  wire tmp28307;
  wire tmp28308;
  wire tmp28309;
  wire tmp28310;
  wire tmp28311;
  wire tmp28312;
  wire tmp28313;
  wire tmp28314;
  wire tmp28315;
  wire tmp28316;
  wire tmp28317;
  wire tmp28318;
  wire tmp28319;
  wire tmp28320;
  wire tmp28321;
  wire tmp28322;
  wire tmp28323;
  wire tmp28324;
  wire tmp28325;
  wire tmp28326;
  wire tmp28327;
  wire tmp28328;
  wire tmp28329;
  wire tmp28330;
  wire tmp28331;
  wire tmp28332;
  wire tmp28333;
  wire tmp28334;
  wire tmp28335;
  wire tmp28336;
  wire tmp28337;
  wire tmp28338;
  wire tmp28339;
  wire tmp28340;
  wire tmp28341;
  wire tmp28342;
  wire tmp28343;
  wire tmp28344;
  wire tmp28345;
  wire tmp28346;
  wire tmp28347;
  wire tmp28348;
  wire tmp28349;
  wire tmp28350;
  wire tmp28351;
  wire tmp28352;
  wire tmp28353;
  wire tmp28354;
  wire tmp28355;
  wire tmp28356;
  wire tmp28357;
  wire tmp28358;
  wire tmp28359;
  wire tmp28360;
  wire tmp28361;
  wire tmp28362;
  wire tmp28363;
  wire tmp28364;
  wire tmp28365;
  wire tmp28366;
  wire tmp28367;
  wire tmp28368;
  wire tmp28369;
  wire tmp28370;
  wire tmp28371;
  wire tmp28372;
  wire tmp28373;
  wire tmp28374;
  wire tmp28375;
  wire tmp28376;
  wire tmp28377;
  wire tmp28378;
  wire tmp28379;
  wire tmp28380;
  wire tmp28381;
  wire tmp28382;
  wire tmp28383;
  wire tmp28384;
  wire tmp28385;
  wire tmp28386;
  wire tmp28387;
  wire tmp28388;
  wire tmp28389;
  wire tmp28390;
  wire tmp28391;
  wire tmp28392;
  wire tmp28393;
  wire tmp28394;
  wire tmp28395;
  wire tmp28396;
  wire tmp28397;
  wire tmp28398;
  wire tmp28399;
  wire tmp28400;
  wire tmp28401;
  wire tmp28402;
  wire tmp28403;
  wire tmp28404;
  wire tmp28405;
  wire tmp28406;
  wire tmp28407;
  wire tmp28408;
  wire tmp28409;
  wire tmp28410;
  wire tmp28411;
  wire tmp28412;
  wire tmp28413;
  wire tmp28414;
  wire tmp28415;
  wire tmp28416;
  wire tmp28417;
  wire tmp28418;
  wire tmp28419;
  wire tmp28420;
  wire tmp28421;
  wire tmp28422;
  wire tmp28423;
  wire tmp28424;
  wire tmp28425;
  wire tmp28426;
  wire tmp28427;
  wire tmp28428;
  wire tmp28429;
  wire tmp28430;
  wire tmp28431;
  wire tmp28432;
  wire tmp28433;
  wire tmp28434;
  wire tmp28435;
  wire tmp28436;
  wire tmp28437;
  wire tmp28438;
  wire tmp28439;
  wire tmp28440;
  wire tmp28441;
  wire tmp28442;
  wire tmp28443;
  wire tmp28444;
  wire tmp28445;
  wire tmp28446;
  wire tmp28447;
  wire tmp28448;
  wire tmp28449;
  wire tmp28450;
  wire tmp28451;
  wire tmp28452;
  wire tmp28453;
  wire tmp28454;
  wire tmp28455;
  wire tmp28456;
  wire tmp28457;
  wire tmp28458;
  wire tmp28459;
  wire tmp28460;
  wire tmp28461;
  wire tmp28462;
  wire tmp28463;
  wire tmp28464;
  wire tmp28465;
  wire tmp28466;
  wire tmp28467;
  wire tmp28468;
  wire tmp28469;
  wire tmp28470;
  wire tmp28471;
  wire tmp28472;
  wire tmp28473;
  wire tmp28474;
  wire tmp28475;
  wire tmp28476;
  wire tmp28477;
  wire tmp28478;
  wire tmp28479;
  wire tmp28480;
  wire tmp28481;
  wire tmp28482;
  wire tmp28483;
  wire tmp28484;
  wire tmp28485;
  wire tmp28486;
  wire tmp28487;
  wire tmp28488;
  wire tmp28489;
  wire tmp28490;
  wire tmp28491;
  wire tmp28492;
  wire tmp28493;
  wire tmp28494;
  wire tmp28495;
  wire tmp28496;
  wire tmp28497;
  wire tmp28498;
  wire tmp28499;
  wire tmp28500;
  wire tmp28501;
  wire tmp28502;
  wire tmp28503;
  wire tmp28504;
  wire tmp28505;
  wire tmp28506;
  wire tmp28507;
  wire tmp28508;
  wire tmp28509;
  wire tmp28510;
  wire tmp28511;
  wire tmp28512;
  wire tmp28513;
  wire tmp28514;
  wire tmp28515;
  wire tmp28516;
  wire tmp28517;
  wire tmp28518;
  wire tmp28519;
  wire tmp28520;
  wire tmp28521;
  wire tmp28522;
  wire tmp28523;
  wire tmp28524;
  wire tmp28525;
  wire tmp28526;
  wire tmp28527;
  wire tmp28528;
  wire tmp28529;
  wire tmp28530;
  wire tmp28531;
  wire tmp28532;
  wire tmp28533;
  wire tmp28534;
  wire tmp28535;
  wire tmp28536;
  wire tmp28537;
  wire tmp28538;
  wire tmp28539;
  wire tmp28540;
  wire tmp28541;
  wire tmp28542;
  wire tmp28543;
  wire tmp28544;
  wire tmp28545;
  wire tmp28546;
  wire tmp28547;
  wire tmp28548;
  wire tmp28549;
  wire tmp28550;
  wire tmp28551;
  wire tmp28552;
  wire tmp28553;
  wire tmp28554;
  wire tmp28555;
  wire tmp28556;
  wire tmp28557;
  wire tmp28558;
  wire tmp28559;
  wire tmp28560;
  wire tmp28561;
  wire tmp28562;
  wire tmp28563;
  wire tmp28564;
  wire tmp28565;
  wire tmp28566;
  wire tmp28567;
  wire tmp28568;
  wire tmp28569;
  wire tmp28570;
  wire tmp28571;
  wire tmp28572;
  wire tmp28573;
  wire tmp28574;
  wire tmp28575;
  wire tmp28576;
  wire tmp28577;
  wire tmp28578;
  wire tmp28579;
  wire tmp28580;
  wire tmp28581;
  wire tmp28582;
  wire tmp28583;
  wire tmp28584;
  wire tmp28585;
  wire tmp28586;
  wire tmp28587;
  wire tmp28588;
  wire tmp28589;
  wire tmp28590;
  wire tmp28591;
  wire tmp28592;
  wire tmp28593;
  wire tmp28594;
  wire tmp28595;
  wire tmp28596;
  wire tmp28597;
  wire tmp28598;
  wire tmp28599;
  wire tmp28600;
  wire tmp28601;
  wire tmp28602;
  wire tmp28603;
  wire tmp28604;
  wire tmp28605;
  wire tmp28606;
  wire tmp28607;
  wire tmp28608;
  wire tmp28609;
  wire tmp28610;
  wire tmp28611;
  wire tmp28612;
  wire tmp28613;
  wire tmp28614;
  wire tmp28615;
  wire tmp28616;
  wire tmp28617;
  wire tmp28618;
  wire tmp28619;
  wire tmp28620;
  wire tmp28621;
  wire tmp28622;
  wire tmp28623;
  wire tmp28624;
  wire tmp28625;
  wire tmp28626;
  wire tmp28627;
  wire tmp28628;
  wire tmp28629;
  wire tmp28630;
  wire tmp28631;
  wire tmp28632;
  wire tmp28633;
  wire tmp28634;
  wire tmp28635;
  wire tmp28636;
  wire tmp28637;
  wire tmp28638;
  wire tmp28639;
  wire tmp28640;
  wire tmp28641;
  wire tmp28642;
  wire tmp28643;
  wire tmp28644;
  wire tmp28645;
  wire tmp28646;
  wire tmp28647;
  wire tmp28648;
  wire tmp28649;
  wire tmp28650;
  wire tmp28651;
  wire tmp28652;
  wire tmp28653;
  wire tmp28654;
  wire tmp28655;
  wire tmp28656;
  wire tmp28657;
  wire tmp28658;
  wire tmp28659;
  wire tmp28660;
  wire tmp28661;
  wire tmp28662;
  wire tmp28663;
  wire tmp28664;
  wire tmp28665;
  wire tmp28666;
  wire tmp28667;
  wire tmp28668;
  wire tmp28669;
  wire tmp28670;
  wire tmp28671;
  wire tmp28672;
  wire tmp28673;
  wire tmp28674;
  wire tmp28675;
  wire tmp28676;
  wire tmp28677;
  wire tmp28678;
  wire tmp28679;
  wire tmp28680;
  wire tmp28681;
  wire tmp28682;
  wire tmp28683;
  wire tmp28684;
  wire tmp28685;
  wire tmp28686;
  wire tmp28687;
  wire tmp28688;
  wire tmp28689;
  wire tmp28690;
  wire tmp28691;
  wire tmp28692;
  wire tmp28693;
  wire tmp28694;
  wire tmp28695;
  wire tmp28696;
  wire tmp28697;
  wire tmp28698;
  wire tmp28699;
  wire tmp28700;
  wire tmp28701;
  wire tmp28702;
  wire tmp28703;
  wire tmp28704;
  wire tmp28705;
  wire tmp28706;
  wire tmp28707;
  wire tmp28708;
  wire tmp28709;
  wire tmp28710;
  wire tmp28711;
  wire tmp28712;
  wire tmp28713;
  wire tmp28714;
  wire tmp28715;
  wire tmp28716;
  wire tmp28717;
  wire tmp28718;
  wire tmp28719;
  wire tmp28720;
  wire tmp28721;
  wire tmp28722;
  wire tmp28723;
  wire tmp28724;
  wire tmp28725;
  wire tmp28726;
  wire tmp28727;
  wire tmp28728;
  wire tmp28729;
  wire tmp28730;
  wire tmp28731;
  wire tmp28732;
  wire tmp28733;
  wire tmp28734;
  wire tmp28735;
  wire tmp28736;
  wire tmp28737;
  wire tmp28738;
  wire tmp28739;
  wire tmp28740;
  wire tmp28741;
  wire tmp28742;
  wire tmp28743;
  wire tmp28744;
  wire tmp28745;
  wire tmp28746;
  wire tmp28747;
  wire tmp28748;
  wire tmp28749;
  wire tmp28750;
  wire tmp28751;
  wire tmp28752;
  wire tmp28753;
  wire tmp28754;
  wire tmp28755;
  wire tmp28756;
  wire tmp28757;
  wire tmp28758;
  wire tmp28759;
  wire tmp28760;
  wire tmp28761;
  wire tmp28762;
  wire tmp28763;
  wire tmp28764;
  wire tmp28765;
  wire tmp28766;
  wire tmp28767;
  wire tmp28768;
  wire tmp28769;
  wire tmp28770;
  wire tmp28771;
  wire tmp28772;
  wire tmp28773;
  wire tmp28774;
  wire tmp28775;
  wire tmp28776;
  wire tmp28777;
  wire tmp28778;
  wire tmp28779;
  wire tmp28780;
  wire tmp28781;
  wire tmp28782;
  wire tmp28783;
  wire tmp28784;
  wire tmp28785;
  wire tmp28786;
  wire tmp28787;
  wire tmp28788;
  wire tmp28789;
  wire tmp28790;
  wire tmp28791;
  wire tmp28792;
  wire tmp28793;
  wire tmp28794;
  wire tmp28795;
  wire tmp28796;
  wire tmp28797;
  wire tmp28798;
  wire tmp28799;
  wire tmp28800;
  wire tmp28801;
  wire tmp28802;
  wire tmp28803;
  wire tmp28804;
  wire tmp28805;
  wire tmp28806;
  wire tmp28807;
  wire tmp28808;
  wire tmp28809;
  wire tmp28810;
  wire tmp28811;
  wire tmp28812;
  wire tmp28813;
  wire tmp28814;
  wire tmp28815;
  wire tmp28816;
  wire tmp28817;
  wire tmp28818;
  wire tmp28819;
  wire tmp28820;
  wire tmp28821;
  wire tmp28822;
  wire tmp28823;
  wire tmp28824;
  wire tmp28825;
  wire tmp28826;
  wire tmp28827;
  wire tmp28828;
  wire tmp28829;
  wire tmp28830;
  wire tmp28831;
  wire tmp28832;
  wire tmp28833;
  wire tmp28834;
  wire tmp28835;
  wire tmp28836;
  wire tmp28837;
  wire tmp28838;
  wire tmp28839;
  wire tmp28840;
  wire tmp28841;
  wire tmp28842;
  wire tmp28843;
  wire tmp28844;
  wire tmp28845;
  wire tmp28846;
  wire tmp28847;
  wire tmp28848;
  wire tmp28849;
  wire tmp28850;
  wire tmp28851;
  wire tmp28852;
  wire tmp28853;
  wire tmp28854;
  wire tmp28855;
  wire tmp28856;
  wire tmp28857;
  wire tmp28858;
  wire tmp28859;
  wire tmp28860;
  wire tmp28861;
  wire tmp28862;
  wire tmp28863;
  wire tmp28864;
  wire tmp28865;
  wire tmp28866;
  wire tmp28867;
  wire tmp28868;
  wire tmp28869;
  wire tmp28870;
  wire tmp28871;
  wire tmp28872;
  wire tmp28873;
  wire tmp28874;
  wire tmp28875;
  wire tmp28876;
  wire tmp28877;
  wire tmp28878;
  wire tmp28879;
  wire tmp28880;
  wire tmp28881;
  wire tmp28882;
  wire tmp28883;
  wire tmp28884;
  wire tmp28885;
  wire tmp28886;
  wire tmp28887;
  wire tmp28888;
  wire tmp28889;
  wire tmp28890;
  wire tmp28891;
  wire tmp28892;
  wire tmp28893;
  wire tmp28894;
  wire tmp28895;
  wire tmp28896;
  wire tmp28897;
  wire tmp28898;
  wire tmp28899;
  wire tmp28900;
  wire tmp28901;
  wire tmp28902;
  wire tmp28903;
  wire tmp28904;
  wire tmp28905;
  wire tmp28906;
  wire tmp28907;
  wire tmp28908;
  wire tmp28909;
  wire tmp28910;
  wire tmp28911;
  wire tmp28912;
  wire tmp28913;
  wire tmp28914;
  wire tmp28915;
  wire tmp28916;
  wire tmp28917;
  wire tmp28918;
  wire tmp28919;
  wire tmp28920;
  wire tmp28921;
  wire tmp28922;
  wire tmp28923;
  wire tmp28924;
  wire tmp28925;
  wire tmp28926;
  wire tmp28927;
  wire tmp28928;
  wire tmp28929;
  wire tmp28930;
  wire tmp28931;
  wire tmp28932;
  wire tmp28933;
  wire tmp28934;
  wire tmp28935;
  wire tmp28936;
  wire tmp28937;
  wire tmp28938;
  wire tmp28939;
  wire tmp28940;
  wire tmp28941;
  wire tmp28942;
  wire tmp28943;
  wire tmp28944;
  wire tmp28945;
  wire tmp28946;
  wire tmp28947;
  wire tmp28948;
  wire tmp28949;
  wire tmp28950;
  wire tmp28951;
  wire tmp28952;
  wire tmp28953;
  wire tmp28954;
  wire tmp28955;
  wire tmp28956;
  wire tmp28957;
  wire tmp28958;
  wire tmp28959;
  wire tmp28960;
  wire tmp28961;
  wire tmp28962;
  wire tmp28963;
  wire tmp28964;
  wire tmp28965;
  wire tmp28966;
  wire tmp28967;
  wire tmp28968;
  wire tmp28969;
  wire tmp28970;
  wire tmp28971;
  wire tmp28972;
  wire tmp28973;
  wire tmp28974;
  wire tmp28975;
  wire tmp28976;
  wire tmp28977;
  wire tmp28978;
  wire tmp28979;
  wire tmp28980;
  wire tmp28981;
  wire tmp28982;
  wire tmp28983;
  wire tmp28984;
  wire tmp28985;
  wire tmp28986;
  wire tmp28987;
  wire tmp28988;
  wire tmp28989;
  wire tmp28990;
  wire tmp28991;
  wire tmp28992;
  wire tmp28993;
  wire tmp28994;
  wire tmp28995;
  wire tmp28996;
  wire tmp28997;
  wire tmp28998;
  wire tmp28999;
  wire tmp29000;
  wire tmp29001;
  wire tmp29002;
  wire tmp29003;
  wire tmp29004;
  wire tmp29005;
  wire tmp29006;
  wire tmp29007;
  wire tmp29008;
  wire tmp29009;
  wire tmp29010;
  wire tmp29011;
  wire tmp29012;
  wire tmp29013;
  wire tmp29014;
  wire tmp29015;
  wire tmp29016;
  wire tmp29017;
  wire tmp29018;
  wire tmp29019;
  wire tmp29020;
  wire tmp29021;
  wire tmp29022;
  wire tmp29023;
  wire tmp29024;
  wire tmp29025;
  wire tmp29026;
  wire tmp29027;
  wire tmp29028;
  wire tmp29029;
  wire tmp29030;
  wire tmp29031;
  wire tmp29032;
  wire tmp29033;
  wire tmp29034;
  wire tmp29035;
  wire tmp29036;
  wire tmp29037;
  wire tmp29038;
  wire tmp29039;
  wire tmp29040;
  wire tmp29041;
  wire tmp29042;
  wire tmp29043;
  wire tmp29044;
  wire tmp29045;
  wire tmp29046;
  wire tmp29047;
  wire tmp29048;
  wire tmp29049;
  wire tmp29050;
  wire tmp29051;
  wire tmp29052;
  wire tmp29053;
  wire tmp29054;
  wire tmp29055;
  wire tmp29056;
  wire tmp29057;
  wire tmp29058;
  wire tmp29059;
  wire tmp29060;
  wire tmp29061;
  wire tmp29062;
  wire tmp29063;
  wire tmp29064;
  wire tmp29065;
  wire tmp29066;
  wire tmp29067;
  wire tmp29068;
  wire tmp29069;
  wire tmp29070;
  wire tmp29071;
  wire tmp29072;
  wire tmp29073;
  wire tmp29074;
  wire tmp29075;
  wire tmp29076;
  wire tmp29077;
  wire tmp29078;
  wire tmp29079;
  wire tmp29080;
  wire tmp29081;
  wire tmp29082;
  wire tmp29083;
  wire tmp29084;
  wire tmp29085;
  wire tmp29086;
  wire tmp29087;
  wire tmp29088;
  wire tmp29089;
  wire tmp29090;
  wire tmp29091;
  wire tmp29092;
  wire tmp29093;
  wire tmp29094;
  wire tmp29095;
  wire tmp29096;
  wire tmp29097;
  wire tmp29098;
  wire tmp29099;
  wire tmp29100;
  wire tmp29101;
  wire tmp29102;
  wire tmp29103;
  wire tmp29104;
  wire tmp29105;
  wire tmp29106;
  wire tmp29107;
  wire tmp29108;
  wire tmp29109;
  wire tmp29110;
  wire tmp29111;
  wire tmp29112;
  wire tmp29113;
  wire tmp29114;
  wire tmp29115;
  wire tmp29116;
  wire tmp29117;
  wire tmp29118;
  wire tmp29119;
  wire tmp29120;
  wire tmp29121;
  wire tmp29122;
  wire tmp29123;
  wire tmp29124;
  wire tmp29125;
  wire tmp29126;
  wire tmp29127;
  wire tmp29128;
  wire tmp29129;
  wire tmp29130;
  wire tmp29131;
  wire tmp29132;
  wire tmp29133;
  wire tmp29134;
  wire tmp29135;
  wire tmp29136;
  wire tmp29137;
  wire tmp29138;
  wire tmp29139;
  wire tmp29140;
  wire tmp29141;
  wire tmp29142;
  wire tmp29143;
  wire tmp29144;
  wire tmp29145;
  wire tmp29146;
  wire tmp29147;
  wire tmp29148;
  wire tmp29149;
  wire tmp29150;
  wire tmp29151;
  wire tmp29152;
  wire tmp29153;
  wire tmp29154;
  wire tmp29155;
  wire tmp29156;
  wire tmp29157;
  wire tmp29158;
  wire tmp29159;
  wire tmp29160;
  wire tmp29161;
  wire tmp29162;
  wire tmp29163;
  wire tmp29164;
  wire tmp29165;
  wire tmp29166;
  wire tmp29167;
  wire tmp29168;
  wire tmp29169;
  wire tmp29170;
  wire tmp29171;
  wire tmp29172;
  wire tmp29173;
  wire tmp29174;
  wire tmp29175;
  wire tmp29176;
  wire tmp29177;
  wire tmp29178;
  wire tmp29179;
  wire tmp29180;
  wire tmp29181;
  wire tmp29182;
  wire tmp29183;
  wire tmp29184;
  wire tmp29185;
  wire tmp29186;
  wire tmp29187;
  wire tmp29188;
  wire tmp29189;
  wire tmp29190;
  wire tmp29191;
  wire tmp29192;
  wire tmp29193;
  wire tmp29194;
  wire tmp29195;
  wire tmp29196;
  wire tmp29197;
  wire tmp29198;
  wire tmp29199;
  wire tmp29200;
  wire tmp29201;
  wire tmp29202;
  wire tmp29203;
  wire tmp29204;
  wire tmp29205;
  wire tmp29206;
  wire tmp29207;
  wire tmp29208;
  wire tmp29209;
  wire tmp29210;
  wire tmp29211;
  wire tmp29212;
  wire tmp29213;
  wire tmp29214;
  wire tmp29215;
  wire tmp29216;
  wire tmp29217;
  wire tmp29218;
  wire tmp29219;
  wire tmp29220;
  wire tmp29221;
  wire tmp29222;
  wire tmp29223;
  wire tmp29224;
  wire tmp29225;
  wire tmp29226;
  wire tmp29227;
  wire tmp29228;
  wire tmp29229;
  wire tmp29230;
  wire tmp29231;
  wire tmp29232;
  wire tmp29233;
  wire tmp29234;
  wire tmp29235;
  wire tmp29236;
  wire tmp29237;
  wire tmp29238;
  wire tmp29239;
  wire tmp29240;
  wire tmp29241;
  wire tmp29242;
  wire tmp29243;
  wire tmp29244;
  wire tmp29245;
  wire tmp29246;
  wire tmp29247;
  wire tmp29248;
  wire tmp29249;
  wire tmp29250;
  wire tmp29251;
  wire tmp29252;
  wire tmp29253;
  wire tmp29254;
  wire tmp29255;
  wire tmp29256;
  wire tmp29257;
  wire tmp29258;
  wire tmp29259;
  wire tmp29260;
  wire tmp29261;
  wire tmp29262;
  wire tmp29263;
  wire tmp29264;
  wire tmp29265;
  wire tmp29266;
  wire tmp29267;
  wire tmp29268;
  wire tmp29269;
  wire tmp29270;
  wire tmp29271;
  wire tmp29272;
  wire tmp29273;
  wire tmp29274;
  wire tmp29275;
  wire tmp29276;
  wire tmp29277;
  wire tmp29278;
  wire tmp29279;
  wire tmp29280;
  wire tmp29281;
  wire tmp29282;
  wire tmp29283;
  wire tmp29284;
  wire tmp29285;
  wire tmp29286;
  wire tmp29287;
  wire tmp29288;
  wire tmp29289;
  wire tmp29290;
  wire tmp29291;
  wire tmp29292;
  wire tmp29293;
  wire tmp29294;
  wire tmp29295;
  wire tmp29296;
  wire tmp29297;
  wire tmp29298;
  wire tmp29299;
  wire tmp29300;
  wire tmp29301;
  wire tmp29302;
  wire tmp29303;
  wire tmp29304;
  wire tmp29305;
  wire tmp29306;
  wire tmp29307;
  wire tmp29308;
  wire tmp29309;
  wire tmp29310;
  wire tmp29311;
  wire tmp29312;
  wire tmp29313;
  wire tmp29314;
  wire tmp29315;
  wire tmp29316;
  wire tmp29317;
  wire tmp29318;
  wire tmp29319;
  wire tmp29320;
  wire tmp29321;
  wire tmp29322;
  wire tmp29323;
  wire tmp29324;
  wire tmp29325;
  wire tmp29326;
  wire tmp29327;
  wire tmp29328;
  wire tmp29329;
  wire tmp29330;
  wire tmp29331;
  wire tmp29332;
  wire tmp29333;
  wire tmp29334;
  wire tmp29335;
  wire tmp29336;
  wire tmp29337;
  wire tmp29338;
  wire tmp29339;
  wire tmp29340;
  wire tmp29341;
  wire tmp29342;
  wire tmp29343;
  wire tmp29344;
  wire tmp29345;
  wire tmp29346;
  wire tmp29347;
  wire tmp29348;
  wire tmp29349;
  wire tmp29350;
  wire tmp29351;
  wire tmp29352;
  wire tmp29353;
  wire tmp29354;
  wire tmp29355;
  wire tmp29356;
  wire tmp29357;
  wire tmp29358;
  wire tmp29359;
  wire tmp29360;
  wire tmp29361;
  wire tmp29362;
  wire tmp29363;
  wire tmp29364;
  wire tmp29365;
  wire tmp29366;
  wire tmp29367;
  wire tmp29368;
  wire tmp29369;
  wire tmp29370;
  wire tmp29371;
  wire tmp29372;
  wire tmp29373;
  wire tmp29374;
  wire tmp29375;
  wire tmp29376;
  wire tmp29377;
  wire tmp29378;
  wire tmp29379;
  wire tmp29380;
  wire tmp29381;
  wire tmp29382;
  wire tmp29383;
  wire tmp29384;
  wire tmp29385;
  wire tmp29386;
  wire tmp29387;
  wire tmp29388;
  wire tmp29389;
  wire tmp29390;
  wire tmp29391;
  wire tmp29392;
  wire tmp29393;
  wire tmp29394;
  wire tmp29395;
  wire tmp29396;
  wire tmp29397;
  wire tmp29398;
  wire tmp29399;
  wire tmp29400;
  wire tmp29401;
  wire tmp29402;
  wire tmp29403;
  wire tmp29404;
  wire tmp29405;
  wire tmp29406;
  wire tmp29407;
  wire tmp29408;
  wire tmp29409;
  wire tmp29410;
  wire tmp29411;
  wire tmp29412;
  wire tmp29413;
  wire tmp29414;
  wire tmp29415;
  wire tmp29416;
  wire tmp29417;
  wire tmp29418;
  wire tmp29419;
  wire tmp29420;
  wire tmp29421;
  wire tmp29422;
  wire tmp29423;
  wire tmp29424;
  wire tmp29425;
  wire tmp29426;
  wire tmp29427;
  wire tmp29428;
  wire tmp29429;
  wire tmp29430;
  wire tmp29431;
  wire tmp29432;
  wire tmp29433;
  wire tmp29434;
  wire tmp29435;
  wire tmp29436;
  wire tmp29437;
  wire tmp29438;
  wire tmp29439;
  wire tmp29440;
  wire tmp29441;
  wire tmp29442;
  wire tmp29443;
  wire tmp29444;
  wire tmp29445;
  wire tmp29446;
  wire tmp29447;
  wire tmp29448;
  wire tmp29449;
  wire tmp29450;
  wire tmp29451;
  wire tmp29452;
  wire tmp29453;
  wire tmp29454;
  wire tmp29455;
  wire tmp29456;
  wire tmp29457;
  wire tmp29458;
  wire tmp29459;
  wire tmp29460;
  wire tmp29461;
  wire tmp29462;
  wire tmp29463;
  wire tmp29464;
  wire tmp29465;
  wire tmp29466;
  wire tmp29467;
  wire tmp29468;
  wire tmp29469;
  wire tmp29470;
  wire tmp29471;
  wire tmp29472;
  wire tmp29473;
  wire tmp29474;
  wire tmp29475;
  wire tmp29476;
  wire tmp29477;
  wire tmp29478;
  wire tmp29479;
  wire tmp29480;
  wire tmp29481;
  wire tmp29482;
  wire tmp29483;
  wire tmp29484;
  wire tmp29485;
  wire tmp29486;
  wire tmp29487;
  wire tmp29488;
  wire tmp29489;
  wire tmp29490;
  wire tmp29491;
  wire tmp29492;
  wire tmp29493;
  wire tmp29494;
  wire tmp29495;
  wire tmp29496;
  wire tmp29497;
  wire tmp29498;
  wire tmp29499;
  wire tmp29500;
  wire tmp29501;
  wire tmp29502;
  wire tmp29503;
  wire tmp29504;
  wire tmp29505;
  wire tmp29506;
  wire tmp29507;
  wire tmp29508;
  wire tmp29509;
  wire tmp29510;
  wire tmp29511;
  wire tmp29512;
  wire tmp29513;
  wire tmp29514;
  wire tmp29515;
  wire tmp29516;
  wire tmp29517;
  wire tmp29518;
  wire tmp29519;
  wire tmp29520;
  wire tmp29521;
  wire tmp29522;
  wire tmp29523;
  wire tmp29524;
  wire tmp29525;
  wire tmp29526;
  wire tmp29527;
  wire tmp29528;
  wire tmp29529;
  wire tmp29530;
  wire tmp29531;
  wire tmp29532;
  wire tmp29533;
  wire tmp29534;
  wire tmp29535;
  wire tmp29536;
  wire tmp29537;
  wire tmp29538;
  wire tmp29539;
  wire tmp29540;
  wire tmp29541;
  wire tmp29542;
  wire tmp29543;
  wire tmp29544;
  wire tmp29545;
  wire tmp29546;
  wire tmp29547;
  wire tmp29548;
  wire tmp29549;
  wire tmp29550;
  wire tmp29551;
  wire tmp29552;
  wire tmp29553;
  wire tmp29554;
  wire tmp29555;
  wire tmp29556;
  wire tmp29557;
  wire tmp29558;
  wire tmp29559;
  wire tmp29560;
  wire tmp29561;
  wire tmp29562;
  wire tmp29563;
  wire tmp29564;
  wire tmp29565;
  wire tmp29566;
  wire tmp29567;
  wire tmp29568;
  wire tmp29569;
  wire tmp29570;
  wire tmp29571;
  wire tmp29572;
  wire tmp29573;
  wire tmp29574;
  wire tmp29575;
  wire tmp29576;
  wire tmp29577;
  wire tmp29578;
  wire tmp29579;
  wire tmp29580;
  wire tmp29581;
  wire tmp29582;
  wire tmp29583;
  wire tmp29584;
  wire tmp29585;
  wire tmp29586;
  wire tmp29587;
  wire tmp29588;
  wire tmp29589;
  wire tmp29590;
  wire tmp29591;
  wire tmp29592;
  wire tmp29593;
  wire tmp29594;
  wire tmp29595;
  wire tmp29596;
  wire tmp29597;
  wire tmp29598;
  wire tmp29599;
  wire tmp29600;
  wire tmp29601;
  wire tmp29602;
  wire tmp29603;
  wire tmp29604;
  wire tmp29605;
  wire tmp29606;
  wire tmp29607;
  wire tmp29608;
  wire tmp29609;
  wire tmp29610;
  wire tmp29611;
  wire tmp29612;
  wire tmp29613;
  wire tmp29614;
  wire tmp29615;
  wire tmp29616;
  wire tmp29617;
  wire tmp29618;
  wire tmp29619;
  wire tmp29620;
  wire tmp29621;
  wire tmp29622;
  wire tmp29623;
  wire tmp29624;
  wire tmp29625;
  wire tmp29626;
  wire tmp29627;
  wire tmp29628;
  wire tmp29629;
  wire tmp29630;
  wire tmp29631;
  wire tmp29632;
  wire tmp29633;
  wire tmp29634;
  wire tmp29635;
  wire tmp29636;
  wire tmp29637;
  wire tmp29638;
  wire tmp29639;
  wire tmp29640;
  wire tmp29641;
  wire tmp29642;
  wire tmp29643;
  wire tmp29644;
  wire tmp29645;
  wire tmp29646;
  wire tmp29647;
  wire tmp29648;
  wire tmp29649;
  wire tmp29650;
  wire tmp29651;
  wire tmp29652;
  wire tmp29653;
  wire tmp29654;
  wire tmp29655;
  wire tmp29656;
  wire tmp29657;
  wire tmp29658;
  wire tmp29659;
  wire tmp29660;
  wire tmp29661;
  wire tmp29662;
  wire tmp29663;
  wire tmp29664;
  wire tmp29665;
  wire tmp29666;
  wire tmp29667;
  wire tmp29668;
  wire tmp29669;
  wire tmp29670;
  wire tmp29671;
  wire tmp29672;
  wire tmp29673;
  wire tmp29674;
  wire tmp29675;
  wire tmp29676;
  wire tmp29677;
  wire tmp29678;
  wire tmp29679;
  wire tmp29680;
  wire tmp29681;
  wire tmp29682;
  wire tmp29683;
  wire tmp29684;
  wire tmp29685;
  wire tmp29686;
  wire tmp29687;
  wire tmp29688;
  wire tmp29689;
  wire tmp29690;
  wire tmp29691;
  wire tmp29692;
  wire tmp29693;
  wire tmp29694;
  wire tmp29695;
  wire tmp29696;
  wire tmp29697;
  wire tmp29698;
  wire tmp29699;
  wire tmp29700;
  wire tmp29701;
  wire tmp29702;
  wire tmp29703;
  wire tmp29704;
  wire tmp29705;
  wire tmp29706;
  wire tmp29707;
  wire tmp29708;
  wire tmp29709;
  wire tmp29710;
  wire tmp29711;
  wire tmp29712;
  wire tmp29713;
  wire tmp29714;
  wire tmp29715;
  wire tmp29716;
  wire tmp29717;
  wire tmp29718;
  wire tmp29719;
  wire tmp29720;
  wire tmp29721;
  wire tmp29722;
  wire tmp29723;
  wire tmp29724;
  wire tmp29725;
  wire tmp29726;
  wire tmp29727;
  wire tmp29728;
  wire tmp29729;
  wire tmp29730;
  wire tmp29731;
  wire tmp29732;
  wire tmp29733;
  wire tmp29734;
  wire tmp29735;
  wire tmp29736;
  wire tmp29737;
  wire tmp29738;
  wire tmp29739;
  wire tmp29740;
  wire tmp29741;
  wire tmp29742;
  wire tmp29743;
  wire tmp29744;
  wire tmp29745;
  wire tmp29746;
  wire tmp29747;
  wire tmp29748;
  wire tmp29749;
  wire tmp29750;
  wire tmp29751;
  wire tmp29752;
  wire tmp29753;
  wire tmp29754;
  wire tmp29755;
  wire tmp29756;
  wire tmp29757;
  wire tmp29758;
  wire tmp29759;
  wire tmp29760;
  wire tmp29761;
  wire tmp29762;
  wire tmp29763;
  wire tmp29764;
  wire tmp29765;
  wire tmp29766;
  wire tmp29767;
  wire tmp29768;
  wire tmp29769;
  wire tmp29770;
  wire tmp29771;
  wire tmp29772;
  wire tmp29773;
  wire tmp29774;
  wire tmp29775;
  wire tmp29776;
  wire tmp29777;
  wire tmp29778;
  wire tmp29779;
  wire tmp29780;
  wire tmp29781;
  wire tmp29782;
  wire tmp29783;
  wire tmp29784;
  wire tmp29785;
  wire tmp29786;
  wire tmp29787;
  wire tmp29788;
  wire tmp29789;
  wire tmp29790;
  wire tmp29791;
  wire tmp29792;
  wire tmp29793;
  wire tmp29794;
  wire tmp29795;
  wire tmp29796;
  wire tmp29797;
  wire tmp29798;
  wire tmp29799;
  wire tmp29800;
  wire tmp29801;
  wire tmp29802;
  wire tmp29803;
  wire tmp29804;
  wire tmp29805;
  wire tmp29806;
  wire tmp29807;
  wire tmp29808;
  wire tmp29809;
  wire tmp29810;
  wire tmp29811;
  wire tmp29812;
  wire tmp29813;
  wire tmp29814;
  wire tmp29815;
  wire tmp29816;
  wire tmp29817;
  wire tmp29818;
  wire tmp29819;
  wire tmp29820;
  wire tmp29821;
  wire tmp29822;
  wire tmp29823;
  wire tmp29824;
  wire tmp29825;
  wire tmp29826;
  wire tmp29827;
  wire tmp29828;
  wire tmp29829;
  wire tmp29830;
  wire tmp29831;
  wire tmp29832;
  wire tmp29833;
  wire tmp29834;
  wire tmp29835;
  wire tmp29836;
  wire tmp29837;
  wire tmp29838;
  wire tmp29839;
  wire tmp29840;
  wire tmp29841;
  wire tmp29842;
  wire tmp29843;
  wire tmp29844;
  wire tmp29845;
  wire tmp29846;
  wire tmp29847;
  wire tmp29848;
  wire tmp29849;
  wire tmp29850;
  wire tmp29851;
  wire tmp29852;
  wire tmp29853;
  wire tmp29854;
  wire tmp29855;
  wire tmp29856;
  wire tmp29857;
  wire tmp29858;
  wire tmp29859;
  wire tmp29860;
  wire tmp29861;
  wire tmp29862;
  wire tmp29863;
  wire tmp29864;
  wire tmp29865;
  wire tmp29866;
  wire tmp29867;
  wire tmp29868;
  wire tmp29869;
  wire tmp29870;
  wire tmp29871;
  wire tmp29872;
  wire tmp29873;
  wire tmp29874;
  wire tmp29875;
  wire tmp29876;
  wire tmp29877;
  wire tmp29878;
  wire tmp29879;
  wire tmp29880;
  wire tmp29881;
  wire tmp29882;
  wire tmp29883;
  wire tmp29884;
  wire tmp29885;
  wire tmp29886;
  wire tmp29887;
  wire tmp29888;
  wire tmp29889;
  wire tmp29890;
  wire tmp29891;
  wire tmp29892;
  wire tmp29893;
  wire tmp29894;
  wire tmp29895;
  wire tmp29896;
  wire tmp29897;
  wire tmp29898;
  wire tmp29899;
  wire tmp29900;
  wire tmp29901;
  wire tmp29902;
  wire tmp29903;
  wire tmp29904;
  wire tmp29905;
  wire tmp29906;
  wire tmp29907;
  wire tmp29908;
  wire tmp29909;
  wire tmp29910;
  wire tmp29911;
  wire tmp29912;
  wire tmp29913;
  wire tmp29914;
  wire tmp29915;
  wire tmp29916;
  wire tmp29917;
  wire tmp29918;
  wire tmp29919;
  wire tmp29920;
  wire tmp29921;
  wire tmp29922;
  wire tmp29923;
  wire tmp29924;
  wire tmp29925;
  wire tmp29926;
  wire tmp29927;
  wire tmp29928;
  wire tmp29929;
  wire tmp29930;
  wire tmp29931;
  wire tmp29932;
  wire tmp29933;
  wire tmp29934;
  wire tmp29935;
  wire tmp29936;
  wire tmp29937;
  wire tmp29938;
  wire tmp29939;
  wire tmp29940;
  wire tmp29941;
  wire tmp29942;
  wire tmp29943;
  wire tmp29944;
  wire tmp29945;
  wire tmp29946;
  wire tmp29947;
  wire tmp29948;
  wire tmp29949;
  wire tmp29950;
  wire tmp29951;
  wire tmp29952;
  wire tmp29953;
  wire tmp29954;
  wire tmp29955;
  wire tmp29956;
  wire tmp29957;
  wire tmp29958;
  wire tmp29959;
  wire tmp29960;
  wire tmp29961;
  wire tmp29962;
  wire tmp29963;
  wire tmp29964;
  wire tmp29965;
  wire tmp29966;
  wire tmp29967;
  wire tmp29968;
  wire tmp29969;
  wire tmp29970;
  wire tmp29971;
  wire tmp29972;
  wire tmp29973;
  wire tmp29974;
  wire tmp29975;
  wire tmp29976;
  wire tmp29977;
  wire tmp29978;
  wire tmp29979;
  wire tmp29980;
  wire tmp29981;
  wire tmp29982;
  wire tmp29983;
  wire tmp29984;
  wire tmp29985;
  wire tmp29986;
  wire tmp29987;
  wire tmp29988;
  wire tmp29989;
  wire tmp29990;
  wire tmp29991;
  wire tmp29992;
  wire tmp29993;
  wire tmp29994;
  wire tmp29995;
  wire tmp29996;
  wire tmp29997;
  wire tmp29998;
  wire tmp29999;
  wire tmp30000;
  wire tmp30001;
  wire tmp30002;
  wire tmp30003;
  wire tmp30004;
  wire tmp30005;
  wire tmp30006;
  wire tmp30007;
  wire tmp30008;
  wire tmp30009;
  wire tmp30010;
  wire tmp30011;
  wire tmp30012;
  wire tmp30013;
  wire tmp30014;
  wire tmp30015;
  wire tmp30016;
  wire tmp30017;
  wire tmp30018;
  wire tmp30019;
  wire tmp30020;
  wire tmp30021;
  wire tmp30022;
  wire tmp30023;
  wire tmp30024;
  wire tmp30025;
  wire tmp30026;
  wire tmp30027;
  wire tmp30028;
  wire tmp30029;
  wire tmp30030;
  wire tmp30031;
  wire tmp30032;
  wire tmp30033;
  wire tmp30034;
  wire tmp30035;
  wire tmp30036;
  wire tmp30037;
  wire tmp30038;
  wire tmp30039;
  wire tmp30040;
  wire tmp30041;
  wire tmp30042;
  wire tmp30043;
  wire tmp30044;
  wire tmp30045;
  wire tmp30046;
  wire tmp30047;
  wire tmp30048;
  wire tmp30049;
  wire tmp30050;
  wire tmp30051;
  wire tmp30052;
  wire tmp30053;
  wire tmp30054;
  wire tmp30055;
  wire tmp30056;
  wire tmp30057;
  wire tmp30058;
  wire tmp30059;
  wire tmp30060;
  wire tmp30061;
  wire tmp30062;
  wire tmp30063;
  wire tmp30064;
  wire tmp30065;
  wire tmp30066;
  wire tmp30067;
  wire tmp30068;
  wire tmp30069;
  wire tmp30070;
  wire tmp30071;
  wire tmp30072;
  wire tmp30073;
  wire tmp30074;
  wire tmp30075;
  wire tmp30076;
  wire tmp30077;
  wire tmp30078;
  wire tmp30079;
  wire tmp30080;
  wire tmp30081;
  wire tmp30082;
  wire tmp30083;
  wire tmp30084;
  wire tmp30085;
  wire tmp30086;
  wire tmp30087;
  wire tmp30088;
  wire tmp30089;
  wire tmp30090;
  wire tmp30091;
  wire tmp30092;
  wire tmp30093;
  wire tmp30094;
  wire tmp30095;
  wire tmp30096;
  wire tmp30097;
  wire tmp30098;
  wire tmp30099;
  wire tmp30100;
  wire tmp30101;
  wire tmp30102;
  wire tmp30103;
  wire tmp30104;
  wire tmp30105;
  wire tmp30106;
  wire tmp30107;
  wire tmp30108;
  wire tmp30109;
  wire tmp30110;
  wire tmp30111;
  wire tmp30112;
  wire tmp30113;
  wire tmp30114;
  wire tmp30115;
  wire tmp30116;
  wire tmp30117;
  wire tmp30118;
  wire tmp30119;
  wire tmp30120;
  wire tmp30121;
  wire tmp30122;
  wire tmp30123;
  wire tmp30124;
  wire tmp30125;
  wire tmp30126;
  wire tmp30127;
  wire tmp30128;
  wire tmp30129;
  wire tmp30130;
  wire tmp30131;
  wire tmp30132;
  wire tmp30133;
  wire tmp30134;
  wire tmp30135;
  wire tmp30136;
  wire tmp30137;
  wire tmp30138;
  wire tmp30139;
  wire tmp30140;
  wire tmp30141;
  wire tmp30142;
  wire tmp30143;
  wire tmp30144;
  wire tmp30145;
  wire tmp30146;
  wire tmp30147;
  wire tmp30148;
  wire tmp30149;
  wire tmp30150;
  wire tmp30151;
  wire tmp30152;
  wire tmp30153;
  wire tmp30154;
  wire tmp30155;
  wire tmp30156;
  wire tmp30157;
  wire tmp30158;
  wire tmp30159;
  wire tmp30160;
  wire tmp30161;
  wire tmp30162;
  wire tmp30163;
  wire tmp30164;
  wire tmp30165;
  wire tmp30166;
  wire tmp30167;
  wire tmp30168;
  wire tmp30169;
  wire tmp30170;
  wire tmp30171;
  wire tmp30172;
  wire tmp30173;
  wire tmp30174;
  wire tmp30175;
  wire tmp30176;
  wire tmp30177;
  wire tmp30178;
  wire tmp30179;
  wire tmp30180;
  wire tmp30181;
  wire tmp30182;
  wire tmp30183;
  wire tmp30184;
  wire tmp30185;
  wire tmp30186;
  wire tmp30187;
  wire tmp30188;
  wire tmp30189;
  wire tmp30190;
  wire tmp30191;
  wire tmp30192;
  wire tmp30193;
  wire tmp30194;
  wire tmp30195;
  wire tmp30196;
  wire tmp30197;
  wire tmp30198;
  wire tmp30199;
  wire tmp30200;
  wire tmp30201;
  wire tmp30202;
  wire tmp30203;
  wire tmp30204;
  wire tmp30205;
  wire tmp30206;
  wire tmp30207;
  wire tmp30208;
  wire tmp30209;
  wire tmp30210;
  wire tmp30211;
  wire tmp30212;
  wire tmp30213;
  wire tmp30214;
  wire tmp30215;
  wire tmp30216;
  wire tmp30217;
  wire tmp30218;
  wire tmp30219;
  wire tmp30220;
  wire tmp30221;
  wire tmp30222;
  wire tmp30223;
  wire tmp30224;
  wire tmp30225;
  wire tmp30226;
  wire tmp30227;
  wire tmp30228;
  wire tmp30229;
  wire tmp30230;
  wire tmp30231;
  wire tmp30232;
  wire tmp30233;
  wire tmp30234;
  wire tmp30235;
  wire tmp30236;
  wire tmp30237;
  wire tmp30238;
  wire tmp30239;
  wire tmp30240;
  wire tmp30241;
  wire tmp30242;
  wire tmp30243;
  wire tmp30244;
  wire tmp30245;
  wire tmp30246;
  wire tmp30247;
  wire tmp30248;
  wire tmp30249;
  wire tmp30250;
  wire tmp30251;
  wire tmp30252;
  wire tmp30253;
  wire tmp30254;
  wire tmp30255;
  wire tmp30256;
  wire tmp30257;
  wire tmp30258;
  wire tmp30259;
  wire tmp30260;
  wire tmp30261;
  wire tmp30262;
  wire tmp30263;
  wire tmp30264;
  wire tmp30265;
  wire tmp30266;
  wire tmp30267;
  wire tmp30268;
  wire tmp30269;
  wire tmp30270;
  wire tmp30271;
  wire tmp30272;
  wire tmp30273;
  wire tmp30274;
  wire tmp30275;
  wire tmp30276;
  wire tmp30277;
  wire tmp30278;
  wire tmp30279;
  wire tmp30280;
  wire tmp30281;
  wire tmp30282;
  wire tmp30283;
  wire tmp30284;
  wire tmp30285;
  wire tmp30286;
  wire tmp30287;
  wire tmp30288;
  wire tmp30289;
  wire tmp30290;
  wire tmp30291;
  wire tmp30292;
  wire tmp30293;
  wire tmp30294;
  wire tmp30295;
  wire tmp30296;
  wire tmp30297;
  wire tmp30298;
  wire tmp30299;
  wire tmp30300;
  wire tmp30301;
  wire tmp30302;
  wire tmp30303;
  wire tmp30304;
  wire tmp30305;
  wire tmp30306;
  wire tmp30307;
  wire tmp30308;
  wire tmp30309;
  wire tmp30310;
  wire tmp30311;
  wire tmp30312;
  wire tmp30313;
  wire tmp30314;
  wire tmp30315;
  wire tmp30316;
  wire tmp30317;
  wire tmp30318;
  wire tmp30319;
  wire tmp30320;
  wire tmp30321;
  wire tmp30322;
  wire tmp30323;
  wire tmp30324;
  wire tmp30325;
  wire tmp30326;
  wire tmp30327;
  wire tmp30328;
  wire tmp30329;
  wire tmp30330;
  wire tmp30331;
  wire tmp30332;
  wire tmp30333;
  wire tmp30334;
  wire tmp30335;
  wire tmp30336;
  wire tmp30337;
  wire tmp30338;
  wire tmp30339;
  wire tmp30340;
  wire tmp30341;
  wire tmp30342;
  wire tmp30343;
  wire tmp30344;
  wire tmp30345;
  wire tmp30346;
  wire tmp30347;
  wire tmp30348;
  wire tmp30349;
  wire tmp30350;
  wire tmp30351;
  wire tmp30352;
  wire tmp30353;
  wire tmp30354;
  wire tmp30355;
  wire tmp30356;
  wire tmp30357;
  wire tmp30358;
  wire tmp30359;
  wire tmp30360;
  wire tmp30361;
  wire tmp30362;
  wire tmp30363;
  wire tmp30364;
  wire tmp30365;
  wire tmp30366;
  wire tmp30367;
  wire tmp30368;
  wire tmp30369;
  wire tmp30370;
  wire tmp30371;
  wire tmp30372;
  wire tmp30373;
  wire tmp30374;
  wire tmp30375;
  wire tmp30376;
  wire tmp30377;
  wire tmp30378;
  wire tmp30379;
  wire tmp30380;
  wire tmp30381;
  wire tmp30382;
  wire tmp30383;
  wire tmp30384;
  wire tmp30385;
  wire tmp30386;
  wire tmp30387;
  wire tmp30388;
  wire tmp30389;
  wire tmp30390;
  wire tmp30391;
  wire tmp30392;
  wire tmp30393;
  wire tmp30394;
  wire tmp30395;
  wire tmp30396;
  wire tmp30397;
  wire tmp30398;
  wire tmp30399;
  wire tmp30400;
  wire tmp30401;
  wire tmp30402;
  wire tmp30403;
  wire tmp30404;
  wire tmp30405;
  wire tmp30406;
  wire tmp30407;
  wire tmp30408;
  wire tmp30409;
  wire tmp30410;
  wire tmp30411;
  wire tmp30412;
  wire tmp30413;
  wire tmp30414;
  wire tmp30415;
  wire tmp30416;
  wire tmp30417;
  wire tmp30418;
  wire tmp30419;
  wire tmp30420;
  wire tmp30421;
  wire tmp30422;
  wire tmp30423;
  wire tmp30424;
  wire tmp30425;
  wire tmp30426;
  wire tmp30427;
  wire tmp30428;
  wire tmp30429;
  wire tmp30430;
  wire tmp30431;
  wire tmp30432;
  wire tmp30433;
  wire tmp30434;
  wire tmp30435;
  wire tmp30436;
  wire tmp30437;
  wire tmp30438;
  wire tmp30439;
  wire tmp30440;
  wire tmp30441;
  wire tmp30442;
  wire tmp30443;
  wire tmp30444;
  wire tmp30445;
  wire tmp30446;
  wire tmp30447;
  wire tmp30448;
  wire tmp30449;
  wire tmp30450;
  wire tmp30451;
  wire tmp30452;
  wire tmp30453;
  wire tmp30454;
  wire tmp30455;
  wire tmp30456;
  wire tmp30457;
  wire tmp30458;
  wire tmp30459;
  wire tmp30460;
  wire tmp30461;
  wire tmp30462;
  wire tmp30463;
  wire tmp30464;
  wire tmp30465;
  wire tmp30466;
  wire tmp30467;
  wire tmp30468;
  wire tmp30469;
  wire tmp30470;
  wire tmp30471;
  wire tmp30472;
  wire tmp30473;
  wire tmp30474;
  wire tmp30475;
  wire tmp30476;
  wire tmp30477;
  wire tmp30478;
  wire tmp30479;
  wire tmp30480;
  wire tmp30481;
  wire tmp30482;
  wire tmp30483;
  wire tmp30484;
  wire tmp30485;
  wire tmp30486;
  wire tmp30487;
  wire tmp30488;
  wire tmp30489;
  wire tmp30490;
  wire tmp30491;
  wire tmp30492;
  wire tmp30493;
  wire tmp30494;
  wire tmp30495;
  wire tmp30496;
  wire tmp30497;
  wire tmp30498;
  wire tmp30499;
  wire tmp30500;
  wire tmp30501;
  wire tmp30502;
  wire tmp30503;
  wire tmp30504;
  wire tmp30505;
  wire tmp30506;
  wire tmp30507;
  wire tmp30508;
  wire tmp30509;
  wire tmp30510;
  wire tmp30511;
  wire tmp30512;
  wire tmp30513;
  wire tmp30514;
  wire tmp30515;
  wire tmp30516;
  wire tmp30517;
  wire tmp30518;
  wire tmp30519;
  wire tmp30520;
  wire tmp30521;
  wire tmp30522;
  wire tmp30523;
  wire tmp30524;
  wire tmp30525;
  wire tmp30526;
  wire tmp30527;
  wire tmp30528;
  wire tmp30529;
  wire tmp30530;
  wire tmp30531;
  wire tmp30532;
  wire tmp30533;
  wire tmp30534;
  wire tmp30535;
  wire tmp30536;
  wire tmp30537;
  wire tmp30538;
  wire tmp30539;
  wire tmp30540;
  wire tmp30541;
  wire tmp30542;
  wire tmp30543;
  wire tmp30544;
  wire tmp30545;
  wire tmp30546;
  wire tmp30547;
  wire tmp30548;
  wire tmp30549;
  wire tmp30550;
  wire tmp30551;
  wire tmp30552;
  wire tmp30553;
  wire tmp30554;
  wire tmp30555;
  wire tmp30556;
  wire tmp30557;
  wire tmp30558;
  wire tmp30559;
  wire tmp30560;
  wire tmp30561;
  wire tmp30562;
  wire tmp30563;
  wire tmp30564;
  wire tmp30565;
  wire tmp30566;
  wire tmp30567;
  wire tmp30568;
  wire tmp30569;
  wire tmp30570;
  wire tmp30571;
  wire tmp30572;
  wire tmp30573;
  wire tmp30574;
  wire tmp30575;
  wire tmp30576;
  wire tmp30577;
  wire tmp30578;
  wire tmp30579;
  wire tmp30580;
  wire tmp30581;
  wire tmp30582;
  wire tmp30583;
  wire tmp30584;
  wire tmp30585;
  wire tmp30586;
  wire tmp30587;
  wire tmp30588;
  wire tmp30589;
  wire tmp30590;
  wire tmp30591;
  wire tmp30592;
  wire tmp30593;
  wire tmp30594;
  wire tmp30595;
  wire tmp30596;
  wire tmp30597;
  wire tmp30598;
  wire tmp30599;
  wire tmp30600;
  wire tmp30601;
  wire tmp30602;
  wire tmp30603;
  wire tmp30604;
  wire tmp30605;
  wire tmp30606;
  wire tmp30607;
  wire tmp30608;
  wire tmp30609;
  wire tmp30610;
  wire tmp30611;
  wire tmp30612;
  wire tmp30613;
  wire tmp30614;
  wire tmp30615;
  wire tmp30616;
  wire tmp30617;
  wire tmp30618;
  wire tmp30619;
  wire tmp30620;
  wire tmp30621;
  wire tmp30622;
  wire tmp30623;
  wire tmp30624;
  wire tmp30625;
  wire tmp30626;
  wire tmp30627;
  wire tmp30628;
  wire tmp30629;
  wire tmp30630;
  wire tmp30631;
  wire tmp30632;
  wire tmp30633;
  wire tmp30634;
  wire tmp30635;
  wire tmp30636;
  wire tmp30637;
  wire tmp30638;
  wire tmp30639;
  wire tmp30640;
  wire tmp30641;
  wire tmp30642;
  wire tmp30643;
  wire tmp30644;
  wire tmp30645;
  wire tmp30646;
  wire tmp30647;
  wire tmp30648;
  wire tmp30649;
  wire tmp30650;
  wire tmp30651;
  wire tmp30652;
  wire tmp30653;
  wire tmp30654;
  wire tmp30655;
  wire tmp30656;
  wire tmp30657;
  wire tmp30658;
  wire tmp30659;
  wire tmp30660;
  wire tmp30661;
  wire tmp30662;
  wire tmp30663;
  wire tmp30664;
  wire tmp30665;
  wire tmp30666;
  wire tmp30667;
  wire tmp30668;
  wire tmp30669;
  wire tmp30670;
  wire tmp30671;
  wire tmp30672;
  wire tmp30673;
  wire tmp30674;
  wire tmp30675;
  wire tmp30676;
  wire tmp30677;
  wire tmp30678;
  wire tmp30679;
  wire tmp30680;
  wire tmp30681;
  wire tmp30682;
  wire tmp30683;
  wire tmp30684;
  wire tmp30685;
  wire tmp30686;
  wire tmp30687;
  wire tmp30688;
  wire tmp30689;
  wire tmp30690;
  wire tmp30691;
  wire tmp30692;
  wire tmp30693;
  wire tmp30694;
  wire tmp30695;
  wire tmp30696;
  wire tmp30697;
  wire tmp30698;
  wire tmp30699;
  wire tmp30700;
  wire tmp30701;
  wire tmp30702;
  wire tmp30703;
  wire tmp30704;
  wire tmp30705;
  wire tmp30706;
  wire tmp30707;
  wire tmp30708;
  wire tmp30709;
  wire tmp30710;
  wire tmp30711;
  wire tmp30712;
  wire tmp30713;
  wire tmp30714;
  wire tmp30715;
  wire tmp30716;
  wire tmp30717;
  wire tmp30718;
  wire tmp30719;
  wire tmp30720;
  wire tmp30721;
  wire tmp30722;
  wire tmp30723;
  wire tmp30724;
  wire tmp30725;
  wire tmp30726;
  wire tmp30727;
  wire tmp30728;
  wire tmp30729;
  wire tmp30730;
  wire tmp30731;
  wire tmp30732;
  wire tmp30733;
  wire tmp30734;
  wire tmp30735;
  wire tmp30736;
  wire tmp30737;
  wire tmp30738;
  wire tmp30739;
  wire tmp30740;
  wire tmp30741;
  wire tmp30742;
  wire tmp30743;
  wire tmp30744;
  wire tmp30745;
  wire tmp30746;
  wire tmp30747;
  wire tmp30748;
  wire tmp30749;
  wire tmp30750;
  wire tmp30751;
  wire tmp30752;
  wire tmp30753;
  wire tmp30754;
  wire tmp30755;
  wire tmp30756;
  wire tmp30757;
  wire tmp30758;
  wire tmp30759;
  wire tmp30760;
  wire tmp30761;
  wire tmp30762;
  wire tmp30763;
  wire tmp30764;
  wire tmp30765;
  wire tmp30766;
  wire tmp30767;
  wire tmp30768;
  wire tmp30769;
  wire tmp30770;
  wire tmp30771;
  wire tmp30772;
  wire tmp30773;
  wire tmp30774;
  wire tmp30775;
  wire tmp30776;
  wire tmp30777;
  wire tmp30778;
  wire tmp30779;
  wire tmp30780;
  wire tmp30781;
  wire tmp30782;
  wire tmp30783;
  wire tmp30784;
  wire tmp30785;
  wire tmp30786;
  wire tmp30787;
  wire tmp30788;
  wire tmp30789;
  wire tmp30790;
  wire tmp30791;
  wire tmp30792;
  wire tmp30793;
  wire tmp30794;
  wire tmp30795;
  wire tmp30796;
  wire tmp30797;
  wire tmp30798;
  wire tmp30799;
  wire tmp30800;
  wire tmp30801;
  wire tmp30802;
  wire tmp30803;
  wire tmp30804;
  wire tmp30805;
  wire tmp30806;
  wire tmp30807;
  wire tmp30808;
  wire tmp30809;
  wire tmp30810;
  wire tmp30811;
  wire tmp30812;
  wire tmp30813;
  wire tmp30814;
  wire tmp30815;
  wire tmp30816;
  wire tmp30817;
  wire tmp30818;
  wire tmp30819;
  wire tmp30820;
  wire tmp30821;
  wire tmp30822;
  wire tmp30823;
  wire tmp30824;
  wire tmp30825;
  wire tmp30826;
  wire tmp30827;
  wire tmp30828;
  wire tmp30829;
  wire tmp30830;
  wire tmp30831;
  wire tmp30832;
  wire tmp30833;
  wire tmp30834;
  wire tmp30835;
  wire tmp30836;
  wire tmp30837;
  wire tmp30838;
  wire tmp30839;
  wire tmp30840;
  wire tmp30841;
  wire tmp30842;
  wire tmp30843;
  wire tmp30844;
  wire tmp30845;
  wire tmp30846;
  wire tmp30847;
  wire tmp30848;
  wire tmp30849;
  wire tmp30850;
  wire tmp30851;
  wire tmp30852;
  wire tmp30853;
  wire tmp30854;
  wire tmp30855;
  wire tmp30856;
  wire tmp30857;
  wire tmp30858;
  wire tmp30859;
  wire tmp30860;
  wire tmp30861;
  wire tmp30862;
  wire tmp30863;
  wire tmp30864;
  wire tmp30865;
  wire tmp30866;
  wire tmp30867;
  wire tmp30868;
  wire tmp30869;
  wire tmp30870;
  wire tmp30871;
  wire tmp30872;
  wire tmp30873;
  wire tmp30874;
  wire tmp30875;
  wire tmp30876;
  wire tmp30877;
  wire tmp30878;
  wire tmp30879;
  wire tmp30880;
  wire tmp30881;
  wire tmp30882;
  wire tmp30883;
  wire tmp30884;
  wire tmp30885;
  wire tmp30886;
  wire tmp30887;
  wire tmp30888;
  wire tmp30889;
  wire tmp30890;
  wire tmp30891;
  wire tmp30892;
  wire tmp30893;
  wire tmp30894;
  wire tmp30895;
  wire tmp30896;
  wire tmp30897;
  wire tmp30898;
  wire tmp30899;
  wire tmp30900;
  wire tmp30901;
  wire tmp30902;
  wire tmp30903;
  wire tmp30904;
  wire tmp30905;
  wire tmp30906;
  wire tmp30907;
  wire tmp30908;
  wire tmp30909;
  wire tmp30910;
  wire tmp30911;
  wire tmp30912;
  wire tmp30913;
  wire tmp30914;
  wire tmp30915;
  wire tmp30916;
  wire tmp30917;
  wire tmp30918;
  wire tmp30919;
  wire tmp30920;
  wire tmp30921;
  wire tmp30922;
  wire tmp30923;
  wire tmp30924;
  wire tmp30925;
  wire tmp30926;
  wire tmp30927;
  wire tmp30928;
  wire tmp30929;
  wire tmp30930;
  wire tmp30931;
  wire tmp30932;
  wire tmp30933;
  wire tmp30934;
  wire tmp30935;
  wire tmp30936;
  wire tmp30937;
  wire tmp30938;
  wire tmp30939;
  wire tmp30940;
  wire tmp30941;
  wire tmp30942;
  wire tmp30943;
  wire tmp30944;
  wire tmp30945;
  wire tmp30946;
  wire tmp30947;
  wire tmp30948;
  wire tmp30949;
  wire tmp30950;
  wire tmp30951;
  wire tmp30952;
  wire tmp30953;
  wire tmp30954;
  wire tmp30955;
  wire tmp30956;
  wire tmp30957;
  wire tmp30958;
  wire tmp30959;
  wire tmp30960;
  wire tmp30961;
  wire tmp30962;
  wire tmp30963;
  wire tmp30964;
  wire tmp30965;
  wire tmp30966;
  wire tmp30967;
  wire tmp30968;
  wire tmp30969;
  wire tmp30970;
  wire tmp30971;
  wire tmp30972;
  wire tmp30973;
  wire tmp30974;
  wire tmp30975;
  wire tmp30976;
  wire tmp30977;
  wire tmp30978;
  wire tmp30979;
  wire tmp30980;
  wire tmp30981;
  wire tmp30982;
  wire tmp30983;
  wire tmp30984;
  wire tmp30985;
  wire tmp30986;
  wire tmp30987;
  wire tmp30988;
  wire tmp30989;
  wire tmp30990;
  wire tmp30991;
  wire tmp30992;
  wire tmp30993;
  wire tmp30994;
  wire tmp30995;
  wire tmp30996;
  wire tmp30997;
  wire tmp30998;
  wire tmp30999;
  wire tmp31000;
  wire tmp31001;
  wire tmp31002;
  wire tmp31003;
  wire tmp31004;
  wire tmp31005;
  wire tmp31006;
  wire tmp31007;
  wire tmp31008;
  wire tmp31009;
  wire tmp31010;
  wire tmp31011;
  wire tmp31012;
  wire tmp31013;
  wire tmp31014;
  wire tmp31015;
  wire tmp31016;
  wire tmp31017;
  wire tmp31018;
  wire tmp31019;
  wire tmp31020;
  wire tmp31021;
  wire tmp31022;
  wire tmp31023;
  wire tmp31024;
  wire tmp31025;
  wire tmp31026;
  wire tmp31027;
  wire tmp31028;
  wire tmp31029;
  wire tmp31030;
  wire tmp31031;
  wire tmp31032;
  wire tmp31033;
  wire tmp31034;
  wire tmp31035;
  wire tmp31036;
  wire tmp31037;
  wire tmp31038;
  wire tmp31039;
  wire tmp31040;
  wire tmp31041;
  wire tmp31042;
  wire tmp31043;
  wire tmp31044;
  wire tmp31045;
  wire tmp31046;
  wire tmp31047;
  wire tmp31048;
  wire tmp31049;
  wire tmp31050;
  wire tmp31051;
  wire tmp31052;
  wire tmp31053;
  wire tmp31054;
  wire tmp31055;
  wire tmp31056;
  wire tmp31057;
  wire tmp31058;
  wire tmp31059;
  wire tmp31060;
  wire tmp31061;
  wire tmp31062;
  wire tmp31063;
  wire tmp31064;
  wire tmp31065;
  wire tmp31066;
  wire tmp31067;
  wire tmp31068;
  wire tmp31069;
  wire tmp31070;
  wire tmp31071;
  wire tmp31072;
  wire tmp31073;
  wire tmp31074;
  wire tmp31075;
  wire tmp31076;
  wire tmp31077;
  wire tmp31078;
  wire tmp31079;
  wire tmp31080;
  wire tmp31081;
  wire tmp31082;
  wire tmp31083;
  wire tmp31084;
  wire tmp31085;
  wire tmp31086;
  wire tmp31087;
  wire tmp31088;
  wire tmp31089;
  wire tmp31090;
  wire tmp31091;
  wire tmp31092;
  wire tmp31093;
  wire tmp31094;
  wire tmp31095;
  wire tmp31096;
  wire tmp31097;
  wire tmp31098;
  wire tmp31099;
  wire tmp31100;
  wire tmp31101;
  wire tmp31102;
  wire tmp31103;
  wire tmp31104;
  wire tmp31105;
  wire tmp31106;
  wire tmp31107;
  wire tmp31108;
  wire tmp31109;
  wire tmp31110;
  wire tmp31111;
  wire tmp31112;
  wire tmp31113;
  wire tmp31114;
  wire tmp31115;
  wire tmp31116;
  wire tmp31117;
  wire tmp31118;
  wire tmp31119;
  wire tmp31120;
  wire tmp31121;
  wire tmp31122;
  wire tmp31123;
  wire tmp31124;
  wire tmp31125;
  wire tmp31126;
  wire tmp31127;
  wire tmp31128;
  wire tmp31129;
  wire tmp31130;
  wire tmp31131;
  wire tmp31132;
  wire tmp31133;
  wire tmp31134;
  wire tmp31135;
  wire tmp31136;
  wire tmp31137;
  wire tmp31138;
  wire tmp31139;
  wire tmp31140;
  wire tmp31141;
  wire tmp31142;
  wire tmp31143;
  wire tmp31144;
  wire tmp31145;
  wire tmp31146;
  wire tmp31147;
  wire tmp31148;
  wire tmp31149;
  wire tmp31150;
  wire tmp31151;
  wire tmp31152;
  wire tmp31153;
  wire tmp31154;
  wire tmp31155;
  wire tmp31156;
  wire tmp31157;
  wire tmp31158;
  wire tmp31159;
  wire tmp31160;
  wire tmp31161;
  wire tmp31162;
  wire tmp31163;
  wire tmp31164;
  wire tmp31165;
  wire tmp31166;
  wire tmp31167;
  wire tmp31168;
  wire tmp31169;
  wire tmp31170;
  wire tmp31171;
  wire tmp31172;
  wire tmp31173;
  wire tmp31174;
  wire tmp31175;
  wire tmp31176;
  wire tmp31177;
  wire tmp31178;
  wire tmp31179;
  wire tmp31180;
  wire tmp31181;
  wire tmp31182;
  wire tmp31183;
  wire tmp31184;
  wire tmp31185;
  wire tmp31186;
  wire tmp31187;
  wire tmp31188;
  wire tmp31189;
  wire tmp31190;
  wire tmp31191;
  wire tmp31192;
  wire tmp31193;
  wire tmp31194;
  wire tmp31195;
  wire tmp31196;
  wire tmp31197;
  wire tmp31198;
  wire tmp31199;
  wire tmp31200;
  wire tmp31201;
  wire tmp31202;
  wire tmp31203;
  wire tmp31204;
  wire tmp31205;
  wire tmp31206;
  wire tmp31207;
  wire tmp31208;
  wire tmp31209;
  wire tmp31210;
  wire tmp31211;
  wire tmp31212;
  wire tmp31213;
  wire tmp31214;
  wire tmp31215;
  wire tmp31216;
  wire tmp31217;
  wire tmp31218;
  wire tmp31219;
  wire tmp31220;
  wire tmp31221;
  wire tmp31222;
  wire tmp31223;
  wire tmp31224;
  wire tmp31225;
  wire tmp31226;
  wire tmp31227;
  wire tmp31228;
  wire tmp31229;
  wire tmp31230;
  wire tmp31231;
  wire tmp31232;
  wire tmp31233;
  wire tmp31234;
  wire tmp31235;
  wire tmp31236;
  wire tmp31237;
  wire tmp31238;
  wire tmp31239;
  wire tmp31240;
  wire tmp31241;
  wire tmp31242;
  wire tmp31243;
  wire tmp31244;
  wire tmp31245;
  wire tmp31246;
  wire tmp31247;
  wire tmp31248;
  wire tmp31249;
  wire tmp31250;
  wire tmp31251;
  wire tmp31252;
  wire tmp31253;
  wire tmp31254;
  wire tmp31255;
  wire tmp31256;
  wire tmp31257;
  wire tmp31258;
  wire tmp31259;
  wire tmp31260;
  wire tmp31261;
  wire tmp31262;
  wire tmp31263;
  wire tmp31264;
  wire tmp31265;
  wire tmp31266;
  wire tmp31267;
  wire tmp31268;
  wire tmp31269;
  wire tmp31270;
  wire tmp31271;
  wire tmp31272;
  wire tmp31273;
  wire tmp31274;
  wire tmp31275;
  wire tmp31276;
  wire tmp31277;
  wire tmp31278;
  wire tmp31279;
  wire tmp31280;
  wire tmp31281;
  wire tmp31282;
  wire tmp31283;
  wire tmp31284;
  wire tmp31285;
  wire tmp31286;
  wire tmp31287;
  wire tmp31288;
  wire tmp31289;
  wire tmp31290;
  wire tmp31291;
  wire tmp31292;
  wire tmp31293;
  wire tmp31294;
  wire tmp31295;
  wire tmp31296;
  wire tmp31297;
  wire tmp31298;
  wire tmp31299;
  wire tmp31300;
  wire tmp31301;
  wire tmp31302;
  wire tmp31303;
  wire tmp31304;
  wire tmp31305;
  wire tmp31306;
  wire tmp31307;
  wire tmp31308;
  wire tmp31309;
  wire tmp31310;
  wire tmp31311;
  wire tmp31312;
  wire tmp31313;
  wire tmp31314;
  wire tmp31315;
  wire tmp31316;
  wire tmp31317;
  wire tmp31318;
  wire tmp31319;
  wire tmp31320;
  wire tmp31321;
  wire tmp31322;
  wire tmp31323;
  wire tmp31324;
  wire tmp31325;
  wire tmp31326;
  wire tmp31327;
  wire tmp31328;
  wire tmp31329;
  wire tmp31330;
  wire tmp31331;
  wire tmp31332;
  wire tmp31333;
  wire tmp31334;
  wire tmp31335;
  wire tmp31336;
  wire tmp31337;
  wire tmp31338;
  wire tmp31339;
  wire tmp31340;
  wire tmp31341;
  wire tmp31342;
  wire tmp31343;
  wire tmp31344;
  wire tmp31345;
  wire tmp31346;
  wire tmp31347;
  wire tmp31348;
  wire tmp31349;
  wire tmp31350;
  wire tmp31351;
  wire tmp31352;
  wire tmp31353;
  wire tmp31354;
  wire tmp31355;
  wire tmp31356;
  wire tmp31357;
  wire tmp31358;
  wire tmp31359;
  wire tmp31360;
  wire tmp31361;
  wire tmp31362;
  wire tmp31363;
  wire tmp31364;
  wire tmp31365;
  wire tmp31366;
  wire tmp31367;
  wire tmp31368;
  wire tmp31369;
  wire tmp31370;
  wire tmp31371;
  wire tmp31372;
  wire tmp31373;
  wire tmp31374;
  wire tmp31375;
  wire tmp31376;
  wire tmp31377;
  wire tmp31378;
  wire tmp31379;
  wire tmp31380;
  wire tmp31381;
  wire tmp31382;
  wire tmp31383;
  wire tmp31384;
  wire tmp31385;
  wire tmp31386;
  wire tmp31387;
  wire tmp31388;
  wire tmp31389;
  wire tmp31390;
  wire tmp31391;
  wire tmp31392;
  wire tmp31393;
  wire tmp31394;
  wire tmp31395;
  wire tmp31396;
  wire tmp31397;
  wire tmp31398;
  wire tmp31399;
  wire tmp31400;
  wire tmp31401;
  wire tmp31402;
  wire tmp31403;
  wire tmp31404;
  wire tmp31405;
  wire tmp31406;
  wire tmp31407;
  wire tmp31408;
  wire tmp31409;
  wire tmp31410;
  wire tmp31411;
  wire tmp31412;
  wire tmp31413;
  wire tmp31414;
  wire tmp31415;
  wire tmp31416;
  wire tmp31417;
  wire tmp31418;
  wire tmp31419;
  wire tmp31420;
  wire tmp31421;
  wire tmp31422;
  wire tmp31423;
  wire tmp31424;
  wire tmp31425;
  wire tmp31426;
  wire tmp31427;
  wire tmp31428;
  wire tmp31429;
  wire tmp31430;
  wire tmp31431;
  wire tmp31432;
  wire tmp31433;
  wire tmp31434;
  wire tmp31435;
  wire tmp31436;
  wire tmp31437;
  wire tmp31438;
  wire tmp31439;
  wire tmp31440;
  wire tmp31441;
  wire tmp31442;
  wire tmp31443;
  wire tmp31444;
  wire tmp31445;
  wire tmp31446;
  wire tmp31447;
  wire tmp31448;
  wire tmp31449;
  wire tmp31450;
  wire tmp31451;
  wire tmp31452;
  wire tmp31453;
  wire tmp31454;
  wire tmp31455;
  wire tmp31456;
  wire tmp31457;
  wire tmp31458;
  wire tmp31459;
  wire tmp31460;
  wire tmp31461;
  wire tmp31462;
  wire tmp31463;
  wire tmp31464;
  wire tmp31465;
  wire tmp31466;
  wire tmp31467;
  wire tmp31468;
  wire tmp31469;
  wire tmp31470;
  wire tmp31471;
  wire tmp31472;
  wire tmp31473;
  wire tmp31474;
  wire tmp31475;
  wire tmp31476;
  wire tmp31477;
  wire tmp31478;
  wire tmp31479;
  wire tmp31480;
  wire tmp31481;
  wire tmp31482;
  wire tmp31483;
  wire tmp31484;
  wire tmp31485;
  wire tmp31486;
  wire tmp31487;
  wire tmp31488;
  wire tmp31489;
  wire tmp31490;
  wire tmp31491;
  wire tmp31492;
  wire tmp31493;
  wire tmp31494;
  wire tmp31495;
  wire tmp31496;
  wire tmp31497;
  wire tmp31498;
  wire tmp31499;
  wire tmp31500;
  wire tmp31501;
  wire tmp31502;
  wire tmp31503;
  wire tmp31504;
  wire tmp31505;
  wire tmp31506;
  wire tmp31507;
  wire tmp31508;
  wire tmp31509;
  wire tmp31510;
  wire tmp31511;
  wire tmp31512;
  wire tmp31513;
  wire tmp31514;
  wire tmp31515;
  wire tmp31516;
  wire tmp31517;
  wire tmp31518;
  wire tmp31519;
  wire tmp31520;
  wire tmp31521;
  wire tmp31522;
  wire tmp31523;
  wire tmp31524;
  wire tmp31525;
  wire tmp31526;
  wire tmp31527;
  wire tmp31528;
  wire tmp31529;
  wire tmp31530;
  wire tmp31531;
  wire tmp31532;
  wire tmp31533;
  wire tmp31534;
  wire tmp31535;
  wire tmp31536;
  wire tmp31537;
  wire tmp31538;
  wire tmp31539;
  wire tmp31540;
  wire tmp31541;
  wire tmp31542;
  wire tmp31543;
  wire tmp31544;
  wire tmp31545;
  wire tmp31546;
  wire tmp31547;
  wire tmp31548;
  wire tmp31549;
  wire tmp31550;
  wire tmp31551;
  wire tmp31552;
  wire tmp31553;
  wire tmp31554;
  wire tmp31555;
  wire tmp31556;
  wire tmp31557;
  wire tmp31558;
  wire tmp31559;
  wire tmp31560;
  wire tmp31561;
  wire tmp31562;
  wire tmp31563;
  wire tmp31564;
  wire tmp31565;
  wire tmp31566;
  wire tmp31567;
  wire tmp31568;
  wire tmp31569;
  wire tmp31570;
  wire tmp31571;
  wire tmp31572;
  wire tmp31573;
  wire tmp31574;
  wire tmp31575;
  wire tmp31576;
  wire tmp31577;
  wire tmp31578;
  wire tmp31579;
  wire tmp31580;
  wire tmp31581;
  wire tmp31582;
  wire tmp31583;
  wire tmp31584;
  wire tmp31585;
  wire tmp31586;
  wire tmp31587;
  wire tmp31588;
  wire tmp31589;
  wire tmp31590;
  wire tmp31591;
  wire tmp31592;
  wire tmp31593;
  wire tmp31594;
  wire tmp31595;
  wire tmp31596;
  wire tmp31597;
  wire tmp31598;
  wire tmp31599;
  wire tmp31600;
  wire tmp31601;
  wire tmp31602;
  wire tmp31603;
  wire tmp31604;
  wire tmp31605;
  wire tmp31606;
  wire tmp31607;
  wire tmp31608;
  wire tmp31609;
  wire tmp31610;
  wire tmp31611;
  wire tmp31612;
  wire tmp31613;
  wire tmp31614;
  wire tmp31615;
  wire tmp31616;
  wire tmp31617;
  wire tmp31618;
  wire tmp31619;
  wire tmp31620;
  wire tmp31621;
  wire tmp31622;
  wire tmp31623;
  wire tmp31624;
  wire tmp31625;
  wire tmp31626;
  wire tmp31627;
  wire tmp31628;
  wire tmp31629;
  wire tmp31630;
  wire tmp31631;
  wire tmp31632;
  wire tmp31633;
  wire tmp31634;
  wire tmp31635;
  wire tmp31636;
  wire tmp31637;
  wire tmp31638;
  wire tmp31639;
  wire tmp31640;
  wire tmp31641;
  wire tmp31642;
  wire tmp31643;
  wire tmp31644;
  wire tmp31645;
  wire tmp31646;
  wire tmp31647;
  wire tmp31648;
  wire tmp31649;
  wire tmp31650;
  wire tmp31651;
  wire tmp31652;
  wire tmp31653;
  wire tmp31654;
  wire tmp31655;
  wire tmp31656;
  wire tmp31657;
  wire tmp31658;
  wire tmp31659;
  wire tmp31660;
  wire tmp31661;
  wire tmp31662;
  wire tmp31663;
  wire tmp31664;
  wire tmp31665;
  wire tmp31666;
  wire tmp31667;
  wire tmp31668;
  wire tmp31669;
  wire tmp31670;
  wire tmp31671;
  wire tmp31672;
  wire tmp31673;
  wire tmp31674;
  wire tmp31675;
  wire tmp31676;
  wire tmp31677;
  wire tmp31678;
  wire tmp31679;
  wire tmp31680;
  wire tmp31681;
  wire tmp31682;
  wire tmp31683;
  wire tmp31684;
  wire tmp31685;
  wire tmp31686;
  wire tmp31687;
  wire tmp31688;
  wire tmp31689;
  wire tmp31690;
  wire tmp31691;
  wire tmp31692;
  wire tmp31693;
  wire tmp31694;
  wire tmp31695;
  wire tmp31696;
  wire tmp31697;
  wire tmp31698;
  wire tmp31699;
  wire tmp31700;
  wire tmp31701;
  wire tmp31702;
  wire tmp31703;
  wire tmp31704;
  wire tmp31705;
  wire tmp31706;
  wire tmp31707;
  wire tmp31708;
  wire tmp31709;
  wire tmp31710;
  wire tmp31711;
  wire tmp31712;
  wire tmp31713;
  wire tmp31714;
  wire tmp31715;
  wire tmp31716;
  wire tmp31717;
  wire tmp31718;
  wire tmp31719;
  wire tmp31720;
  wire tmp31721;
  wire tmp31722;
  wire tmp31723;
  wire tmp31724;
  wire tmp31725;
  wire tmp31726;
  wire tmp31727;
  wire tmp31728;
  wire tmp31729;
  wire tmp31730;
  wire tmp31731;
  wire tmp31732;
  wire tmp31733;
  wire tmp31734;
  wire tmp31735;
  wire tmp31736;
  wire tmp31737;
  wire tmp31738;
  wire tmp31739;
  wire tmp31740;
  wire tmp31741;
  wire tmp31742;
  wire tmp31743;
  wire tmp31744;
  wire tmp31745;
  wire tmp31746;
  wire tmp31747;
  wire tmp31748;
  wire tmp31749;
  wire tmp31750;
  wire tmp31751;
  wire tmp31752;
  wire tmp31753;
  wire tmp31754;
  wire tmp31755;
  wire tmp31756;
  wire tmp31757;
  wire tmp31758;
  wire tmp31759;
  wire tmp31760;
  wire tmp31761;
  wire tmp31762;
  wire tmp31763;
  wire tmp31764;
  wire tmp31765;
  wire tmp31766;
  wire tmp31767;
  wire tmp31768;
  wire tmp31769;
  wire tmp31770;
  wire tmp31771;
  wire tmp31772;
  wire tmp31773;
  wire tmp31774;
  wire tmp31775;
  wire tmp31776;
  wire tmp31777;
  wire tmp31778;
  wire tmp31779;
  wire tmp31780;
  wire tmp31781;
  wire tmp31782;
  wire tmp31783;
  wire tmp31784;
  wire tmp31785;
  wire tmp31786;
  wire tmp31787;
  wire tmp31788;
  wire tmp31789;
  wire tmp31790;
  wire tmp31791;
  wire tmp31792;
  wire tmp31793;
  wire tmp31794;
  wire tmp31795;
  wire tmp31796;
  wire tmp31797;
  wire tmp31798;
  wire tmp31799;
  wire tmp31800;
  wire tmp31801;
  wire tmp31802;
  wire tmp31803;
  wire tmp31804;
  wire tmp31805;
  wire tmp31806;
  wire tmp31807;
  wire tmp31808;
  wire tmp31809;
  wire tmp31810;
  wire tmp31811;
  wire tmp31812;
  wire tmp31813;
  wire tmp31814;
  wire tmp31815;
  wire tmp31816;
  wire tmp31817;
  wire tmp31818;
  wire tmp31819;
  wire tmp31820;
  wire tmp31821;
  wire tmp31822;
  wire tmp31823;
  wire tmp31824;
  wire tmp31825;
  wire tmp31826;
  wire tmp31827;
  wire tmp31828;
  wire tmp31829;
  wire tmp31830;
  wire tmp31831;
  wire tmp31832;
  wire tmp31833;
  wire tmp31834;
  wire tmp31835;
  wire tmp31836;
  wire tmp31837;
  wire tmp31838;
  wire tmp31839;
  wire tmp31840;
  wire tmp31841;
  wire tmp31842;
  wire tmp31843;
  wire tmp31844;
  wire tmp31845;
  wire tmp31846;
  wire tmp31847;
  wire tmp31848;
  wire tmp31849;
  wire tmp31850;
  wire tmp31851;
  wire tmp31852;
  wire tmp31853;
  wire tmp31854;
  wire tmp31855;
  wire tmp31856;
  wire tmp31857;
  wire tmp31858;
  wire tmp31859;
  wire tmp31860;
  wire tmp31861;
  wire tmp31862;
  wire tmp31863;
  wire tmp31864;
  wire tmp31865;
  wire tmp31866;
  wire tmp31867;
  wire tmp31868;
  wire tmp31869;
  wire tmp31870;
  wire tmp31871;
  wire tmp31872;
  wire tmp31873;
  wire tmp31874;
  wire tmp31875;
  wire tmp31876;
  wire tmp31877;
  wire tmp31878;
  wire tmp31879;
  wire tmp31880;
  wire tmp31881;
  wire tmp31882;
  wire tmp31883;
  wire tmp31884;
  wire tmp31885;
  wire tmp31886;
  wire tmp31887;
  wire tmp31888;
  wire tmp31889;
  wire tmp31890;
  wire tmp31891;
  wire tmp31892;
  wire tmp31893;
  wire tmp31894;
  wire tmp31895;
  wire tmp31896;
  wire tmp31897;
  wire tmp31898;
  wire tmp31899;
  wire tmp31900;
  wire tmp31901;
  wire tmp31902;
  wire tmp31903;
  wire tmp31904;
  wire tmp31905;
  wire tmp31906;
  wire tmp31907;
  wire tmp31908;
  wire tmp31909;
  wire tmp31910;
  wire tmp31911;
  wire tmp31912;
  wire tmp31913;
  wire tmp31914;
  wire tmp31915;
  wire tmp31916;
  wire tmp31917;
  wire tmp31918;
  wire tmp31919;
  wire tmp31920;
  wire tmp31921;
  wire tmp31922;
  wire tmp31923;
  wire tmp31924;
  wire tmp31925;
  wire tmp31926;
  wire tmp31927;
  wire tmp31928;
  wire tmp31929;
  wire tmp31930;
  wire tmp31931;
  wire tmp31932;
  wire tmp31933;
  wire tmp31934;
  wire tmp31935;
  wire tmp31936;
  wire tmp31937;
  wire tmp31938;
  wire tmp31939;
  wire tmp31940;
  wire tmp31941;
  wire tmp31942;
  wire tmp31943;
  wire tmp31944;
  wire tmp31945;
  wire tmp31946;
  wire tmp31947;
  wire tmp31948;
  wire tmp31949;
  wire tmp31950;
  wire tmp31951;
  wire tmp31952;
  wire tmp31953;
  wire tmp31954;
  wire tmp31955;
  wire tmp31956;
  wire tmp31957;
  wire tmp31958;
  wire tmp31959;
  wire tmp31960;
  wire tmp31961;
  wire tmp31962;
  wire tmp31963;
  wire tmp31964;
  wire tmp31965;
  wire tmp31966;
  wire tmp31967;
  wire tmp31968;
  wire tmp31969;
  wire tmp31970;
  wire tmp31971;
  wire tmp31972;
  wire tmp31973;
  wire tmp31974;
  wire tmp31975;
  wire tmp31976;
  wire tmp31977;
  wire tmp31978;
  wire tmp31979;
  wire tmp31980;
  wire tmp31981;
  wire tmp31982;
  wire tmp31983;
  wire tmp31984;
  wire tmp31985;
  wire tmp31986;
  wire tmp31987;
  wire tmp31988;
  wire tmp31989;
  wire tmp31990;
  wire tmp31991;
  wire tmp31992;
  wire tmp31993;
  wire tmp31994;
  wire tmp31995;
  wire tmp31996;
  wire tmp31997;
  wire tmp31998;
  wire tmp31999;
  wire tmp32000;
  wire tmp32001;
  wire tmp32002;
  wire tmp32003;
  wire tmp32004;
  wire tmp32005;
  wire tmp32006;
  wire tmp32007;
  wire tmp32008;
  wire tmp32009;
  wire tmp32010;
  wire tmp32011;
  wire tmp32012;
  wire tmp32013;
  wire tmp32014;
  wire tmp32015;
  wire tmp32016;
  wire tmp32017;
  wire tmp32018;
  wire tmp32019;
  wire tmp32020;
  wire tmp32021;
  wire tmp32022;
  wire tmp32023;
  wire tmp32024;
  wire tmp32025;
  wire tmp32026;
  wire tmp32027;
  wire tmp32028;
  wire tmp32029;
  wire tmp32030;
  wire tmp32031;
  wire tmp32032;
  wire tmp32033;
  wire tmp32034;
  wire tmp32035;
  wire tmp32036;
  wire tmp32037;
  wire tmp32038;
  wire tmp32039;
  wire tmp32040;
  wire tmp32041;
  wire tmp32042;
  wire tmp32043;
  wire tmp32044;
  wire tmp32045;
  wire tmp32046;
  wire tmp32047;
  wire tmp32048;
  wire tmp32049;
  wire tmp32050;
  wire tmp32051;
  wire tmp32052;
  wire tmp32053;
  wire tmp32054;
  wire tmp32055;
  wire tmp32056;
  wire tmp32057;
  wire tmp32058;
  wire tmp32059;
  wire tmp32060;
  wire tmp32061;
  wire tmp32062;
  wire tmp32063;
  wire tmp32064;
  wire tmp32065;
  wire tmp32066;
  wire tmp32067;
  wire tmp32068;
  wire tmp32069;
  wire tmp32070;
  wire tmp32071;
  wire tmp32072;
  wire tmp32073;
  wire tmp32074;
  wire tmp32075;
  wire tmp32076;
  wire tmp32077;
  wire tmp32078;
  wire tmp32079;
  wire tmp32080;
  wire tmp32081;
  wire tmp32082;
  wire tmp32083;
  wire tmp32084;
  wire tmp32085;
  wire tmp32086;
  wire tmp32087;
  wire tmp32088;
  wire tmp32089;
  wire tmp32090;
  wire tmp32091;
  wire tmp32092;
  wire tmp32093;
  wire tmp32094;
  wire tmp32095;
  wire tmp32096;
  wire tmp32097;
  wire tmp32098;
  wire tmp32099;
  wire tmp32100;
  wire tmp32101;
  wire tmp32102;
  wire tmp32103;
  wire tmp32104;
  wire tmp32105;
  wire tmp32106;
  wire tmp32107;
  wire tmp32108;
  wire tmp32109;
  wire tmp32110;
  wire tmp32111;
  wire tmp32112;
  wire tmp32113;
  wire tmp32114;
  wire tmp32115;
  wire tmp32116;
  wire tmp32117;
  wire tmp32118;
  wire tmp32119;
  wire tmp32120;
  wire tmp32121;
  wire tmp32122;
  wire tmp32123;
  wire tmp32124;
  wire tmp32125;
  wire tmp32126;
  wire tmp32127;
  wire tmp32128;
  wire tmp32129;
  wire tmp32130;
  wire tmp32131;
  wire tmp32132;
  wire tmp32133;
  wire tmp32134;
  wire tmp32135;
  wire tmp32136;
  wire tmp32137;
  wire tmp32138;
  wire tmp32139;
  wire tmp32140;
  wire tmp32141;
  wire tmp32142;
  wire tmp32143;
  wire tmp32144;
  wire tmp32145;
  wire tmp32146;
  wire tmp32147;
  wire tmp32148;
  wire tmp32149;
  wire tmp32150;
  wire tmp32151;
  wire tmp32152;
  wire tmp32153;
  wire tmp32154;
  wire tmp32155;
  wire tmp32156;
  wire tmp32157;
  wire tmp32158;
  wire tmp32159;
  wire tmp32160;
  wire tmp32161;
  wire tmp32162;
  wire tmp32163;
  wire tmp32164;
  wire tmp32165;
  wire tmp32166;
  wire tmp32167;
  wire tmp32168;
  wire tmp32169;
  wire tmp32170;
  wire tmp32171;
  wire tmp32172;
  wire tmp32173;
  wire tmp32174;
  wire tmp32175;
  wire tmp32176;
  wire tmp32177;
  wire tmp32178;
  wire tmp32179;
  wire tmp32180;
  wire tmp32181;
  wire tmp32182;
  wire tmp32183;
  wire tmp32184;
  wire tmp32185;
  wire tmp32186;
  wire tmp32187;
  wire tmp32188;
  wire tmp32189;
  wire tmp32190;
  wire tmp32191;
  wire tmp32192;
  wire tmp32193;
  wire tmp32194;
  wire tmp32195;
  wire tmp32196;
  wire tmp32197;
  wire tmp32198;
  wire tmp32199;
  wire tmp32200;
  wire tmp32201;
  wire tmp32202;
  wire tmp32203;
  wire tmp32204;
  wire tmp32205;
  wire tmp32206;
  wire tmp32207;
  wire tmp32208;
  wire tmp32209;
  wire tmp32210;
  wire tmp32211;
  wire tmp32212;
  wire tmp32213;
  wire tmp32214;
  wire tmp32215;
  wire tmp32216;
  wire tmp32217;
  wire tmp32218;
  wire tmp32219;
  wire tmp32220;
  wire tmp32221;
  wire tmp32222;
  wire tmp32223;
  wire tmp32224;
  wire tmp32225;
  wire tmp32226;
  wire tmp32227;
  wire tmp32228;
  wire tmp32229;
  wire tmp32230;
  wire tmp32231;
  wire tmp32232;
  wire tmp32233;
  wire tmp32234;
  wire tmp32235;
  wire tmp32236;
  wire tmp32237;
  wire tmp32238;
  wire tmp32239;
  wire tmp32240;
  wire tmp32241;
  wire tmp32242;
  wire tmp32243;
  wire tmp32244;
  wire tmp32245;
  wire tmp32246;
  wire tmp32247;
  wire tmp32248;
  wire tmp32249;
  wire tmp32250;
  wire tmp32251;
  wire tmp32252;
  wire tmp32253;
  wire tmp32254;
  wire tmp32255;
  wire tmp32256;
  wire tmp32257;
  wire tmp32258;
  wire tmp32259;
  wire tmp32260;
  wire tmp32261;
  wire tmp32262;
  wire tmp32263;
  wire tmp32264;
  wire tmp32265;
  wire tmp32266;
  wire tmp32267;
  wire tmp32268;
  wire tmp32269;
  wire tmp32270;
  wire tmp32271;
  wire tmp32272;
  wire tmp32273;
  wire tmp32274;
  wire tmp32275;
  wire tmp32276;
  wire tmp32277;
  wire tmp32278;
  wire tmp32279;
  wire tmp32280;
  wire tmp32281;
  wire tmp32282;
  wire tmp32283;
  wire tmp32284;
  wire tmp32285;
  wire tmp32286;
  wire tmp32287;
  wire tmp32288;
  wire tmp32289;
  wire tmp32290;
  wire tmp32291;
  wire tmp32292;
  wire tmp32293;
  wire tmp32294;
  wire tmp32295;
  wire tmp32296;
  wire tmp32297;
  wire tmp32298;
  wire tmp32299;
  wire tmp32300;
  wire tmp32301;
  wire tmp32302;
  wire tmp32303;
  wire tmp32304;
  wire tmp32305;
  wire tmp32306;
  wire tmp32307;
  wire tmp32308;
  wire tmp32309;
  wire tmp32310;
  wire tmp32311;
  wire tmp32312;
  wire tmp32313;
  wire tmp32314;
  wire tmp32315;
  wire tmp32316;
  wire tmp32317;
  wire tmp32318;
  wire tmp32319;
  wire tmp32320;
  wire tmp32321;
  wire tmp32322;
  wire tmp32323;
  wire tmp32324;
  wire tmp32325;
  wire tmp32326;
  wire tmp32327;
  wire tmp32328;
  wire tmp32329;
  wire tmp32330;
  wire tmp32331;
  wire tmp32332;
  wire tmp32333;
  wire tmp32334;
  wire tmp32335;
  wire tmp32336;
  wire tmp32337;
  wire tmp32338;
  wire tmp32339;
  wire tmp32340;
  wire tmp32341;
  wire tmp32342;
  wire tmp32343;
  wire tmp32344;
  wire tmp32345;
  wire tmp32346;
  wire tmp32347;
  wire tmp32348;
  wire tmp32349;
  wire tmp32350;
  wire tmp32351;
  wire tmp32352;
  wire tmp32353;
  wire tmp32354;
  wire tmp32355;
  wire tmp32356;
  wire tmp32357;
  wire tmp32358;
  wire tmp32359;
  wire tmp32360;
  wire tmp32361;
  wire tmp32362;
  wire tmp32363;
  wire tmp32364;
  wire tmp32365;
  wire tmp32366;
  wire tmp32367;
  wire tmp32368;
  wire tmp32369;
  wire tmp32370;
  wire tmp32371;
  wire tmp32372;
  wire tmp32373;
  wire tmp32374;
  wire tmp32375;
  wire tmp32376;
  wire tmp32377;
  wire tmp32378;
  wire tmp32379;
  wire tmp32380;
  wire tmp32381;
  wire tmp32382;
  wire tmp32383;
  wire tmp32384;
  wire tmp32385;
  wire tmp32386;
  wire tmp32387;
  wire tmp32388;
  wire tmp32389;
  wire tmp32390;
  wire tmp32391;
  wire tmp32392;
  wire tmp32393;
  wire tmp32394;
  wire tmp32395;
  wire tmp32396;
  wire tmp32397;
  wire tmp32398;
  wire tmp32399;
  wire tmp32400;
  wire tmp32401;
  wire tmp32402;
  wire tmp32403;
  wire tmp32404;
  wire tmp32405;
  wire tmp32406;
  wire tmp32407;
  wire tmp32408;
  wire tmp32409;
  wire tmp32410;
  wire tmp32411;
  wire tmp32412;
  wire tmp32413;
  wire tmp32414;
  wire tmp32415;
  wire tmp32416;
  wire tmp32417;
  wire tmp32418;
  wire tmp32419;
  wire tmp32420;
  wire tmp32421;
  wire tmp32422;
  wire tmp32423;
  wire tmp32424;
  wire tmp32425;
  wire tmp32426;
  wire tmp32427;
  wire tmp32428;
  wire tmp32429;
  wire tmp32430;
  wire tmp32431;
  wire tmp32432;
  wire tmp32433;
  wire tmp32434;
  wire tmp32435;
  wire tmp32436;
  wire tmp32437;
  wire tmp32438;
  wire tmp32439;
  wire tmp32440;
  wire tmp32441;
  wire tmp32442;
  wire tmp32443;
  wire tmp32444;
  wire tmp32445;
  wire tmp32446;
  wire tmp32447;
  wire tmp32448;
  wire tmp32449;
  wire tmp32450;
  wire tmp32451;
  wire tmp32452;
  wire tmp32453;
  wire tmp32454;
  wire tmp32455;
  wire tmp32456;
  wire tmp32457;
  wire tmp32458;
  wire tmp32459;
  wire tmp32460;
  wire tmp32461;
  wire tmp32462;
  wire tmp32463;
  wire tmp32464;
  wire tmp32465;
  wire tmp32466;
  wire tmp32467;
  wire tmp32468;
  wire tmp32469;
  wire tmp32470;
  wire tmp32471;
  wire tmp32472;
  wire tmp32473;
  wire tmp32474;
  wire tmp32475;
  wire tmp32476;
  wire tmp32477;
  wire tmp32478;
  wire tmp32479;
  wire tmp32480;
  wire tmp32481;
  wire tmp32482;
  wire tmp32483;
  wire tmp32484;
  wire tmp32485;
  wire tmp32486;
  wire tmp32487;
  wire tmp32488;
  wire tmp32489;
  wire tmp32490;
  wire tmp32491;
  wire tmp32492;
  wire tmp32493;
  wire tmp32494;
  wire tmp32495;
  wire tmp32496;
  wire tmp32497;
  wire tmp32498;
  wire tmp32499;
  wire tmp32500;
  wire tmp32501;
  wire tmp32502;
  wire tmp32503;
  wire tmp32504;
  wire tmp32505;
  wire tmp32506;
  wire tmp32507;
  wire tmp32508;
  wire tmp32509;
  wire tmp32510;
  wire tmp32511;
  wire tmp32512;
  wire tmp32513;
  wire tmp32514;
  wire tmp32515;
  wire tmp32516;
  wire tmp32517;
  wire tmp32518;
  wire tmp32519;
  wire tmp32520;
  wire tmp32521;
  wire tmp32522;
  wire tmp32523;
  wire tmp32524;
  wire tmp32525;
  wire tmp32526;
  wire tmp32527;
  wire tmp32528;
  wire tmp32529;
  wire tmp32530;
  wire tmp32531;
  wire tmp32532;
  wire tmp32533;
  wire tmp32534;
  wire tmp32535;
  wire tmp32536;
  wire tmp32537;
  wire tmp32538;
  wire tmp32539;
  wire tmp32540;
  wire tmp32541;
  wire tmp32542;
  wire tmp32543;
  wire tmp32544;
  wire tmp32545;
  wire tmp32546;
  wire tmp32547;
  wire tmp32548;
  wire tmp32549;
  wire tmp32550;
  wire tmp32551;
  wire tmp32552;
  wire tmp32553;
  wire tmp32554;
  wire tmp32555;
  wire tmp32556;
  wire tmp32557;
  wire tmp32558;
  wire tmp32559;
  wire tmp32560;
  wire tmp32561;
  wire tmp32562;
  wire tmp32563;
  wire tmp32564;
  wire tmp32565;
  wire tmp32566;
  wire tmp32567;
  wire tmp32568;
  wire tmp32569;
  wire tmp32570;
  wire tmp32571;
  wire tmp32572;
  wire tmp32573;
  wire tmp32574;
  wire tmp32575;
  wire tmp32576;
  wire tmp32577;
  wire tmp32578;
  wire tmp32579;
  wire tmp32580;
  wire tmp32581;
  wire tmp32582;
  wire tmp32583;
  wire tmp32584;
  wire tmp32585;
  wire tmp32586;
  wire tmp32587;
  wire tmp32588;
  wire tmp32589;
  wire tmp32590;
  wire tmp32591;
  wire tmp32592;
  wire tmp32593;
  wire tmp32594;
  wire tmp32595;
  wire tmp32596;
  wire tmp32597;
  wire tmp32598;
  wire tmp32599;
  wire tmp32600;
  wire tmp32601;
  wire tmp32602;
  wire tmp32603;
  wire tmp32604;
  wire tmp32605;
  wire tmp32606;
  wire tmp32607;
  wire tmp32608;
  wire tmp32609;
  wire tmp32610;
  wire tmp32611;
  wire tmp32612;
  wire tmp32613;
  wire tmp32614;
  wire tmp32615;
  wire tmp32616;
  wire tmp32617;
  wire tmp32618;
  wire tmp32619;
  wire tmp32620;
  wire tmp32621;
  wire tmp32622;
  wire tmp32623;
  wire tmp32624;
  wire tmp32625;
  wire tmp32626;
  wire tmp32627;
  wire tmp32628;
  wire tmp32629;
  wire tmp32630;
  wire tmp32631;
  wire tmp32632;
  wire tmp32633;
  wire tmp32634;
  wire tmp32635;
  wire tmp32636;
  wire tmp32637;
  wire tmp32638;
  wire tmp32639;
  wire tmp32640;
  wire tmp32641;
  wire tmp32642;
  wire tmp32643;
  wire tmp32644;
  wire tmp32645;
  wire tmp32646;
  wire tmp32647;
  wire tmp32648;
  wire tmp32649;
  wire tmp32650;
  wire tmp32651;
  wire tmp32652;
  wire tmp32653;
  wire tmp32654;
  wire tmp32655;
  wire tmp32656;
  wire tmp32657;
  wire tmp32658;
  wire tmp32659;
  wire tmp32660;
  wire tmp32661;
  wire tmp32662;
  wire tmp32663;
  wire tmp32664;
  wire tmp32665;
  wire tmp32666;
  wire tmp32667;
  wire tmp32668;
  wire tmp32669;
  wire tmp32670;
  wire tmp32671;
  wire tmp32672;
  wire tmp32673;
  wire tmp32674;
  wire tmp32675;
  wire tmp32676;
  wire tmp32677;
  wire tmp32678;
  wire tmp32679;
  wire tmp32680;
  wire tmp32681;
  wire tmp32682;
  wire tmp32683;
  wire tmp32684;
  wire tmp32685;
  wire tmp32686;
  wire tmp32687;
  wire tmp32688;
  wire tmp32689;
  wire tmp32690;
  wire tmp32691;
  wire tmp32692;
  wire tmp32693;
  wire tmp32694;
  wire tmp32695;
  wire tmp32696;
  wire tmp32697;
  wire tmp32698;
  wire tmp32699;
  wire tmp32700;
  wire tmp32701;
  wire tmp32702;
  wire tmp32703;
  wire tmp32704;
  wire tmp32705;
  wire tmp32706;
  wire tmp32707;
  wire tmp32708;
  wire tmp32709;
  wire tmp32710;
  wire tmp32711;
  wire tmp32712;
  wire tmp32713;
  wire tmp32714;
  wire tmp32715;
  wire tmp32716;
  wire tmp32717;
  wire tmp32718;
  wire tmp32719;
  wire tmp32720;
  wire tmp32721;
  wire tmp32722;
  wire tmp32723;
  wire tmp32724;
  wire tmp32725;
  wire tmp32726;
  wire tmp32727;
  wire tmp32728;
  wire tmp32729;
  wire tmp32730;
  wire tmp32731;
  wire tmp32732;
  wire tmp32733;
  wire tmp32734;
  wire tmp32735;
  wire tmp32736;
  wire tmp32737;
  wire tmp32738;
  wire tmp32739;
  wire tmp32740;
  wire tmp32741;
  wire tmp32742;
  wire tmp32743;
  wire tmp32744;
  wire tmp32745;
  wire tmp32746;
  wire tmp32747;
  wire tmp32748;
  wire tmp32749;
  wire tmp32750;
  wire tmp32751;
  wire tmp32752;
  wire tmp32753;
  wire tmp32754;
  wire tmp32755;
  wire tmp32756;
  wire tmp32757;
  wire tmp32758;
  wire tmp32759;
  wire tmp32760;
  wire tmp32761;
  wire tmp32762;
  wire tmp32763;
  wire tmp32764;
  wire tmp32765;
  wire tmp32766;
  wire tmp32767;
  wire tmp32768;
  wire tmp32769;
  wire tmp32770;
  wire tmp32771;
  wire tmp32772;
  wire tmp32773;
  wire tmp32774;
  wire tmp32775;
  wire tmp32776;
  wire tmp32777;
  wire tmp32778;
  wire tmp32779;
  wire tmp32780;
  wire tmp32781;
  wire tmp32782;
  wire tmp32783;
  wire tmp32784;
  wire tmp32785;
  wire tmp32786;
  wire tmp32787;
  wire tmp32788;
  wire tmp32789;
  wire tmp32790;
  wire tmp32791;
  wire tmp32792;
  wire tmp32793;
  wire tmp32794;
  wire tmp32795;
  wire tmp32796;
  wire tmp32797;
  wire tmp32798;
  wire tmp32799;
  wire tmp32800;
  wire tmp32801;
  wire tmp32802;
  wire tmp32803;
  wire tmp32804;
  wire tmp32805;
  wire tmp32806;
  wire tmp32807;
  wire tmp32808;
  wire tmp32809;
  wire tmp32810;
  wire tmp32811;
  wire tmp32812;
  wire tmp32813;
  wire tmp32814;
  wire tmp32815;
  wire tmp32816;
  wire tmp32817;
  wire tmp32818;
  wire tmp32819;
  wire tmp32820;
  wire tmp32821;
  wire tmp32822;
  wire tmp32823;
  wire tmp32824;
  wire tmp32825;
  wire tmp32826;
  wire tmp32827;
  wire tmp32828;
  wire tmp32829;
  wire tmp32830;
  wire tmp32831;
  wire tmp32832;
  wire tmp32833;
  wire tmp32834;
  wire tmp32835;
  wire tmp32836;
  wire tmp32837;
  wire tmp32838;
  wire tmp32839;
  wire tmp32840;
  wire tmp32841;
  wire tmp32842;
  wire tmp32843;
  wire tmp32844;
  wire tmp32845;
  wire tmp32846;
  wire tmp32847;
  wire tmp32848;
  wire tmp32849;
  wire tmp32850;
  wire tmp32851;
  wire tmp32852;
  wire tmp32853;
  wire tmp32854;
  wire tmp32855;
  wire tmp32856;
  wire tmp32857;
  wire tmp32858;
  wire tmp32859;
  wire tmp32860;
  wire tmp32861;
  wire tmp32862;
  wire tmp32863;
  wire tmp32864;
  wire tmp32865;
  wire tmp32866;
  wire tmp32867;
  wire tmp32868;
  wire tmp32869;
  wire tmp32870;
  wire tmp32871;
  wire tmp32872;
  wire tmp32873;
  wire tmp32874;
  wire tmp32875;
  wire tmp32876;
  wire tmp32877;
  wire tmp32878;
  wire tmp32879;
  wire tmp32880;
  wire tmp32881;
  wire tmp32882;
  wire tmp32883;
  wire tmp32884;
  wire tmp32885;
  wire tmp32886;
  wire tmp32887;
  wire tmp32888;
  wire tmp32889;
  wire tmp32890;
  wire tmp32891;
  wire tmp32892;
  wire tmp32893;
  wire tmp32894;
  wire tmp32895;
  wire tmp32896;
  wire tmp32897;
  wire tmp32898;
  wire tmp32899;
  wire tmp32900;
  wire tmp32901;
  wire tmp32902;
  wire tmp32903;
  wire tmp32904;
  wire tmp32905;
  wire tmp32906;
  wire tmp32907;
  wire tmp32908;
  wire tmp32909;
  wire tmp32910;
  wire tmp32911;
  wire tmp32912;
  wire tmp32913;
  wire tmp32914;
  wire tmp32915;
  wire tmp32916;
  wire tmp32917;
  wire tmp32918;
  wire tmp32919;
  wire tmp32920;
  wire tmp32921;
  wire tmp32922;
  wire tmp32923;
  wire tmp32924;
  wire tmp32925;
  wire tmp32926;
  wire tmp32927;
  wire tmp32928;
  wire tmp32929;
  wire tmp32930;
  wire tmp32931;
  wire tmp32932;
  wire tmp32933;
  wire tmp32934;
  wire tmp32935;
  wire tmp32936;
  wire tmp32937;
  wire tmp32938;
  wire tmp32939;
  wire tmp32940;
  wire tmp32941;
  wire tmp32942;
  wire tmp32943;
  wire tmp32944;
  wire tmp32945;
  wire tmp32946;
  wire tmp32947;
  wire tmp32948;
  wire tmp32949;
  wire tmp32950;
  wire tmp32951;
  wire tmp32952;
  wire tmp32953;
  wire tmp32954;
  wire tmp32955;
  wire tmp32956;
  wire tmp32957;
  wire tmp32958;
  wire tmp32959;
  wire tmp32960;
  wire tmp32961;
  wire tmp32962;
  wire tmp32963;
  wire tmp32964;
  wire tmp32965;
  wire tmp32966;
  wire tmp32967;
  wire tmp32968;
  wire tmp32969;
  wire tmp32970;
  wire tmp32971;
  wire tmp32972;
  wire tmp32973;
  wire tmp32974;
  wire tmp32975;
  wire tmp32976;
  wire tmp32977;
  wire tmp32978;
  wire tmp32979;
  wire tmp32980;
  wire tmp32981;
  wire tmp32982;
  wire tmp32983;
  wire tmp32984;
  wire tmp32985;
  wire tmp32986;
  wire tmp32987;
  wire tmp32988;
  wire tmp32989;
  wire tmp32990;
  wire tmp32991;
  wire tmp32992;
  wire tmp32993;
  wire tmp32994;
  wire tmp32995;
  wire tmp32996;
  wire tmp32997;
  wire tmp32998;
  wire tmp32999;
  wire tmp33000;
  wire tmp33001;
  wire tmp33002;
  wire tmp33003;
  wire tmp33004;
  wire tmp33005;
  wire tmp33006;
  wire tmp33007;
  wire tmp33008;
  wire tmp33009;
  wire tmp33010;
  wire tmp33011;
  wire tmp33012;
  wire tmp33013;
  wire tmp33014;
  wire tmp33015;
  wire tmp33016;
  wire tmp33017;
  wire tmp33018;
  wire tmp33019;
  wire tmp33020;
  wire tmp33021;
  wire tmp33022;
  wire tmp33023;
  wire tmp33024;
  wire tmp33025;
  wire tmp33026;
  wire tmp33027;
  wire tmp33028;
  wire tmp33029;
  wire tmp33030;
  wire tmp33031;
  wire tmp33032;
  wire tmp33033;
  wire tmp33034;
  wire tmp33035;
  wire tmp33036;
  wire tmp33037;
  wire tmp33038;
  wire tmp33039;
  wire tmp33040;
  wire tmp33041;
  wire tmp33042;
  wire tmp33043;
  wire tmp33044;
  wire tmp33045;
  wire tmp33046;
  wire tmp33047;
  wire tmp33048;
  wire tmp33049;
  wire tmp33050;
  wire tmp33051;
  wire tmp33052;
  wire tmp33053;
  wire tmp33054;
  wire tmp33055;
  wire tmp33056;
  wire tmp33057;
  wire tmp33058;
  wire tmp33059;
  wire tmp33060;
  wire tmp33061;
  wire tmp33062;
  wire tmp33063;
  wire tmp33064;
  wire tmp33065;
  wire tmp33066;
  wire tmp33067;
  wire tmp33068;
  wire tmp33069;
  wire tmp33070;
  wire tmp33071;
  wire tmp33072;
  wire tmp33073;
  wire tmp33074;
  wire tmp33075;
  wire tmp33076;
  wire tmp33077;
  wire tmp33078;
  wire tmp33079;
  wire tmp33080;
  wire tmp33081;
  wire tmp33082;
  wire tmp33083;
  wire tmp33084;
  wire tmp33085;
  wire tmp33086;
  wire tmp33087;
  wire tmp33088;
  wire tmp33089;
  wire tmp33090;
  wire tmp33091;
  wire tmp33092;
  wire tmp33093;
  wire tmp33094;
  wire tmp33095;
  wire tmp33096;
  wire tmp33097;
  wire tmp33098;
  wire tmp33099;
  wire tmp33100;
  wire tmp33101;
  wire tmp33102;
  wire tmp33103;
  wire tmp33104;
  wire tmp33105;
  wire tmp33106;
  wire tmp33107;
  wire tmp33108;
  wire tmp33109;
  wire tmp33110;
  wire tmp33111;
  wire tmp33112;
  wire tmp33113;
  wire tmp33114;
  wire tmp33115;
  wire tmp33116;
  wire tmp33117;
  wire tmp33118;
  wire tmp33119;
  wire tmp33120;
  wire tmp33121;
  wire tmp33122;
  wire tmp33123;
  wire tmp33124;
  wire tmp33125;
  wire tmp33126;
  wire tmp33127;
  wire tmp33128;
  wire tmp33129;
  wire tmp33130;
  wire tmp33131;
  wire tmp33132;
  wire tmp33133;
  wire tmp33134;
  wire tmp33135;
  wire tmp33136;
  wire tmp33137;
  wire tmp33138;
  wire tmp33139;
  wire tmp33140;
  wire tmp33141;
  wire tmp33142;
  wire tmp33143;
  wire tmp33144;
  wire tmp33145;
  wire tmp33146;
  wire tmp33147;
  wire tmp33148;
  wire tmp33149;
  wire tmp33150;
  wire tmp33151;
  wire tmp33152;
  wire tmp33153;
  wire tmp33154;
  wire tmp33155;
  wire tmp33156;
  wire tmp33157;
  wire tmp33158;
  wire tmp33159;
  wire tmp33160;
  wire tmp33161;
  wire tmp33162;
  wire tmp33163;
  wire tmp33164;
  wire tmp33165;
  wire tmp33166;
  wire tmp33167;
  wire tmp33168;
  wire tmp33169;
  wire tmp33170;
  wire tmp33171;
  wire tmp33172;
  wire tmp33173;
  wire tmp33174;
  wire tmp33175;
  wire tmp33176;
  wire tmp33177;
  wire tmp33178;
  wire tmp33179;
  wire tmp33180;
  wire tmp33181;
  wire tmp33182;
  wire tmp33183;
  wire tmp33184;
  wire tmp33185;
  wire tmp33186;
  wire tmp33187;
  wire tmp33188;
  wire tmp33189;
  wire tmp33190;
  wire tmp33191;
  wire tmp33192;
  wire tmp33193;
  wire tmp33194;
  wire tmp33195;
  wire tmp33196;
  wire tmp33197;
  wire tmp33198;
  wire tmp33199;
  wire tmp33200;
  wire tmp33201;
  wire tmp33202;
  wire tmp33203;
  wire tmp33204;
  wire tmp33205;
  wire tmp33206;
  wire tmp33207;
  wire tmp33208;
  wire tmp33209;
  wire tmp33210;
  wire tmp33211;
  wire tmp33212;
  wire tmp33213;
  wire tmp33214;
  wire tmp33215;
  wire tmp33216;
  wire tmp33217;
  wire tmp33218;
  wire tmp33219;
  wire tmp33220;
  wire tmp33221;
  wire tmp33222;
  wire tmp33223;
  wire tmp33224;
  wire tmp33225;
  wire tmp33226;
  wire tmp33227;
  wire tmp33228;
  wire tmp33229;
  wire tmp33230;
  wire tmp33231;
  wire tmp33232;
  wire tmp33233;
  wire tmp33234;
  wire tmp33235;
  wire tmp33236;
  wire tmp33237;
  wire tmp33238;
  wire tmp33239;
  wire tmp33240;
  wire tmp33241;
  wire tmp33242;
  wire tmp33243;
  wire tmp33244;
  wire tmp33245;
  wire tmp33246;
  wire tmp33247;
  wire tmp33248;
  wire tmp33249;
  wire tmp33250;
  wire tmp33251;
  wire tmp33252;
  wire tmp33253;
  wire tmp33254;
  wire tmp33255;
  wire tmp33256;
  wire tmp33257;
  wire tmp33258;
  wire tmp33259;
  wire tmp33260;
  wire tmp33261;
  wire tmp33262;
  wire tmp33263;
  wire tmp33264;
  wire tmp33265;
  wire tmp33266;
  wire tmp33267;
  wire tmp33268;
  wire tmp33269;
  wire tmp33270;
  wire tmp33271;
  wire tmp33272;
  wire tmp33273;
  wire tmp33274;
  wire tmp33275;
  wire tmp33276;
  wire tmp33277;
  wire tmp33278;
  wire tmp33279;
  wire tmp33280;
  wire tmp33281;
  wire tmp33282;
  wire tmp33283;
  wire tmp33284;
  wire tmp33285;
  wire tmp33286;
  wire tmp33287;
  wire tmp33288;
  wire tmp33289;
  wire tmp33290;
  wire tmp33291;
  wire tmp33292;
  wire tmp33293;
  wire tmp33294;
  wire tmp33295;
  wire tmp33296;
  wire tmp33297;
  wire tmp33298;
  wire tmp33299;
  wire tmp33300;
  wire tmp33301;
  wire tmp33302;
  wire tmp33303;
  wire tmp33304;
  wire tmp33305;
  wire tmp33306;
  wire tmp33307;
  wire tmp33308;
  wire tmp33309;
  wire tmp33310;
  wire tmp33311;
  wire tmp33312;
  wire tmp33313;
  wire tmp33314;
  wire tmp33315;
  wire tmp33316;
  wire tmp33317;
  wire tmp33318;
  wire tmp33319;
  wire tmp33320;
  wire tmp33321;
  wire tmp33322;
  wire tmp33323;
  wire tmp33324;
  wire tmp33325;
  wire tmp33326;
  wire tmp33327;
  wire tmp33328;
  wire tmp33329;
  wire tmp33330;
  wire tmp33331;
  wire tmp33332;
  wire tmp33333;
  wire tmp33334;
  wire tmp33335;
  wire tmp33336;
  wire tmp33337;
  wire tmp33338;
  wire tmp33339;
  wire tmp33340;
  wire tmp33341;
  wire tmp33342;
  wire tmp33343;
  wire tmp33344;
  wire tmp33345;
  wire tmp33346;
  wire tmp33347;
  wire tmp33348;
  wire tmp33349;
  wire tmp33350;
  wire tmp33351;
  wire tmp33352;
  wire tmp33353;
  wire tmp33354;
  wire tmp33355;
  wire tmp33356;
  wire tmp33357;
  wire tmp33358;
  wire tmp33359;
  wire tmp33360;
  wire tmp33361;
  wire tmp33362;
  wire tmp33363;
  wire tmp33364;
  wire tmp33365;
  wire tmp33366;
  wire tmp33367;
  wire tmp33368;
  wire tmp33369;
  wire tmp33370;
  wire tmp33371;
  wire tmp33372;
  wire tmp33373;
  wire tmp33374;
  wire tmp33375;
  wire tmp33376;
  wire tmp33377;
  wire tmp33378;
  wire tmp33379;
  wire tmp33380;
  wire tmp33381;
  wire tmp33382;
  wire tmp33383;
  wire tmp33384;
  wire tmp33385;
  wire tmp33386;
  wire tmp33387;
  wire tmp33388;
  wire tmp33389;
  wire tmp33390;
  wire tmp33391;
  wire tmp33392;
  wire tmp33393;
  wire tmp33394;
  wire tmp33395;
  wire tmp33396;
  wire tmp33397;
  wire tmp33398;
  wire tmp33399;
  wire tmp33400;
  wire tmp33401;
  wire tmp33402;
  wire tmp33403;
  wire tmp33404;
  wire tmp33405;
  wire tmp33406;
  wire tmp33407;
  wire tmp33408;
  wire tmp33409;
  wire tmp33410;
  wire tmp33411;
  wire tmp33412;
  wire tmp33413;
  wire tmp33414;
  wire tmp33415;
  wire tmp33416;
  wire tmp33417;
  wire tmp33418;
  wire tmp33419;
  wire tmp33420;
  wire tmp33421;
  wire tmp33422;
  wire tmp33423;
  wire tmp33424;
  wire tmp33425;
  wire tmp33426;
  wire tmp33427;
  wire tmp33428;
  wire tmp33429;
  wire tmp33430;
  wire tmp33431;
  wire tmp33432;
  wire tmp33433;
  wire tmp33434;
  wire tmp33435;
  wire tmp33436;
  wire tmp33437;
  wire tmp33438;
  wire tmp33439;
  wire tmp33440;
  wire tmp33441;
  wire tmp33442;
  wire tmp33443;
  wire tmp33444;
  wire tmp33445;
  wire tmp33446;
  wire tmp33447;
  wire tmp33448;
  wire tmp33449;
  wire tmp33450;
  wire tmp33451;
  wire tmp33452;
  wire tmp33453;
  wire tmp33454;
  wire tmp33455;
  wire tmp33456;
  wire tmp33457;
  wire tmp33458;
  wire tmp33459;
  wire tmp33460;
  wire tmp33461;
  wire tmp33462;
  wire tmp33463;
  wire tmp33464;
  wire tmp33465;
  wire tmp33466;
  wire tmp33467;
  wire tmp33468;
  wire tmp33469;
  wire tmp33470;
  wire tmp33471;
  wire tmp33472;
  wire tmp33473;
  wire tmp33474;
  wire tmp33475;
  wire tmp33476;
  wire tmp33477;
  wire tmp33478;
  wire tmp33479;
  wire tmp33480;
  wire tmp33481;
  wire tmp33482;
  wire tmp33483;
  wire tmp33484;
  wire tmp33485;
  wire tmp33486;
  wire tmp33487;
  wire tmp33488;
  wire tmp33489;
  wire tmp33490;
  wire tmp33491;
  wire tmp33492;
  wire tmp33493;
  wire tmp33494;
  wire tmp33495;
  wire tmp33496;
  wire tmp33497;
  wire tmp33498;
  wire tmp33499;
  wire tmp33500;
  wire tmp33501;
  wire tmp33502;
  wire tmp33503;
  wire tmp33504;
  wire tmp33505;
  wire tmp33506;
  wire tmp33507;
  wire tmp33508;
  wire tmp33509;
  wire tmp33510;
  wire tmp33511;
  wire tmp33512;
  wire tmp33513;
  wire tmp33514;
  wire tmp33515;
  wire tmp33516;
  wire tmp33517;
  wire tmp33518;
  wire tmp33519;
  wire tmp33520;
  wire tmp33521;
  wire tmp33522;
  wire tmp33523;
  wire tmp33524;
  wire tmp33525;
  wire tmp33526;
  wire tmp33527;
  wire tmp33528;
  wire tmp33529;
  wire tmp33530;
  wire tmp33531;
  wire tmp33532;
  wire tmp33533;
  wire tmp33534;
  wire tmp33535;
  wire tmp33536;
  wire tmp33537;
  wire tmp33538;
  wire tmp33539;
  wire tmp33540;
  wire tmp33541;
  wire tmp33542;
  wire tmp33543;
  wire tmp33544;
  wire tmp33545;
  wire tmp33546;
  wire tmp33547;
  wire tmp33548;
  wire tmp33549;
  wire tmp33550;
  wire tmp33551;
  wire tmp33552;
  wire tmp33553;
  wire tmp33554;
  wire tmp33555;
  wire tmp33556;
  wire tmp33557;
  wire tmp33558;
  wire tmp33559;
  wire tmp33560;
  wire tmp33561;
  wire tmp33562;
  wire tmp33563;
  wire tmp33564;
  wire tmp33565;
  wire tmp33566;
  wire tmp33567;
  wire tmp33568;
  wire tmp33569;
  wire tmp33570;
  wire tmp33571;
  wire tmp33572;
  wire tmp33573;
  wire tmp33574;
  wire tmp33575;
  wire tmp33576;
  wire tmp33577;
  wire tmp33578;
  wire tmp33579;
  wire tmp33580;
  wire tmp33581;
  wire tmp33582;
  wire tmp33583;
  wire tmp33584;
  wire tmp33585;
  wire tmp33586;
  wire tmp33587;
  wire tmp33588;
  wire tmp33589;
  wire tmp33590;
  wire tmp33591;
  wire tmp33592;
  wire tmp33593;
  wire tmp33594;
  wire tmp33595;
  wire tmp33596;
  wire tmp33597;
  wire tmp33598;
  wire tmp33599;
  wire tmp33600;
  wire tmp33601;
  wire tmp33602;
  wire tmp33603;
  wire tmp33604;
  wire tmp33605;
  wire tmp33606;
  wire tmp33607;
  wire tmp33608;
  wire tmp33609;
  wire tmp33610;
  wire tmp33611;
  wire tmp33612;
  wire tmp33613;
  wire tmp33614;
  wire tmp33615;
  wire tmp33616;
  wire tmp33617;
  wire tmp33618;
  wire tmp33619;
  wire tmp33620;
  wire tmp33621;
  wire tmp33622;
  wire tmp33623;
  wire tmp33624;
  wire tmp33625;
  wire tmp33626;
  wire tmp33627;
  wire tmp33628;
  wire tmp33629;
  wire tmp33630;
  wire tmp33631;
  wire tmp33632;
  wire tmp33633;
  wire tmp33634;
  wire tmp33635;
  wire tmp33636;
  wire tmp33637;
  wire tmp33638;
  wire tmp33639;
  wire tmp33640;
  wire tmp33641;
  wire tmp33642;
  wire tmp33643;
  wire tmp33644;
  wire tmp33645;
  wire tmp33646;
  wire tmp33647;
  wire tmp33648;
  wire tmp33649;
  wire tmp33650;
  wire tmp33651;
  wire tmp33652;
  wire tmp33653;
  wire tmp33654;
  wire tmp33655;
  wire tmp33656;
  wire tmp33657;
  wire tmp33658;
  wire tmp33659;
  wire tmp33660;
  wire tmp33661;
  wire tmp33662;
  wire tmp33663;
  wire tmp33664;
  wire tmp33665;
  wire tmp33666;
  wire tmp33667;
  wire tmp33668;
  wire tmp33669;
  wire tmp33670;
  wire tmp33671;
  wire tmp33672;
  wire tmp33673;
  wire tmp33674;
  wire tmp33675;
  wire tmp33676;
  wire tmp33677;
  wire tmp33678;
  wire tmp33679;
  wire tmp33680;
  wire tmp33681;
  wire tmp33682;
  wire tmp33683;
  wire tmp33684;
  wire tmp33685;
  wire tmp33686;
  wire tmp33687;
  wire tmp33688;
  wire tmp33689;
  wire tmp33690;
  wire tmp33691;
  wire tmp33692;
  wire tmp33693;
  wire tmp33694;
  wire tmp33695;
  wire tmp33696;
  wire tmp33697;
  wire tmp33698;
  wire tmp33699;
  wire tmp33700;
  wire tmp33701;
  wire tmp33702;
  wire tmp33703;
  wire tmp33704;
  wire tmp33705;
  wire tmp33706;
  wire tmp33707;
  wire tmp33708;
  wire tmp33709;
  wire tmp33710;
  wire tmp33711;
  wire tmp33712;
  wire tmp33713;
  wire tmp33714;
  wire tmp33715;
  wire tmp33716;
  wire tmp33717;
  wire tmp33718;
  wire tmp33719;
  wire tmp33720;
  wire tmp33721;
  wire tmp33722;
  wire tmp33723;
  wire tmp33724;
  wire tmp33725;
  wire tmp33726;
  wire tmp33727;
  wire tmp33728;
  wire tmp33729;
  wire tmp33730;
  wire tmp33731;
  wire tmp33732;
  wire tmp33733;
  wire tmp33734;
  wire tmp33735;
  wire tmp33736;
  wire tmp33737;
  wire tmp33738;
  wire tmp33739;
  wire tmp33740;
  wire tmp33741;
  wire tmp33742;
  wire tmp33743;
  wire tmp33744;
  wire tmp33745;
  wire tmp33746;
  wire tmp33747;
  wire tmp33748;
  wire tmp33749;
  wire tmp33750;
  wire tmp33751;
  wire tmp33752;
  wire tmp33753;
  wire tmp33754;
  wire tmp33755;
  wire tmp33756;
  wire tmp33757;
  wire tmp33758;
  wire tmp33759;
  wire tmp33760;
  wire tmp33761;
  wire tmp33762;
  wire tmp33763;
  wire tmp33764;
  wire tmp33765;
  wire tmp33766;
  wire tmp33767;
  wire tmp33768;
  wire tmp33769;
  wire tmp33770;
  wire tmp33771;
  wire tmp33772;
  wire tmp33773;
  wire tmp33774;
  wire tmp33775;
  wire tmp33776;
  wire tmp33777;
  wire tmp33778;
  wire tmp33779;
  wire tmp33780;
  wire tmp33781;
  wire tmp33782;
  wire tmp33783;
  wire tmp33784;
  wire tmp33785;
  wire tmp33786;
  wire tmp33787;
  wire tmp33788;
  wire tmp33789;
  wire tmp33790;
  wire tmp33791;
  wire tmp33792;
  wire tmp33793;
  wire tmp33794;
  wire tmp33795;
  wire tmp33796;
  wire tmp33797;
  wire tmp33798;
  wire tmp33799;
  wire tmp33800;
  wire tmp33801;
  wire tmp33802;
  wire tmp33803;
  wire tmp33804;
  wire tmp33805;
  wire tmp33806;
  wire tmp33807;
  wire tmp33808;
  wire tmp33809;
  wire tmp33810;
  wire tmp33811;
  wire tmp33812;
  wire tmp33813;
  wire tmp33814;
  wire tmp33815;
  wire tmp33816;
  wire tmp33817;
  wire tmp33818;
  wire tmp33819;
  wire tmp33820;
  wire tmp33821;
  wire tmp33822;
  wire tmp33823;
  wire tmp33824;
  wire tmp33825;
  wire tmp33826;
  wire tmp33827;
  wire tmp33828;
  wire tmp33829;
  wire tmp33830;
  wire tmp33831;
  wire tmp33832;
  wire tmp33833;
  wire tmp33834;
  wire tmp33835;
  wire tmp33836;
  wire tmp33837;
  wire tmp33838;
  wire tmp33839;
  wire tmp33840;
  wire tmp33841;
  wire tmp33842;
  wire tmp33843;
  wire tmp33844;
  wire tmp33845;
  wire tmp33846;
  wire tmp33847;
  wire tmp33848;
  wire tmp33849;
  wire tmp33850;
  wire tmp33851;
  wire tmp33852;
  wire tmp33853;
  wire tmp33854;
  wire tmp33855;
  wire tmp33856;
  wire tmp33857;
  wire tmp33858;
  wire tmp33859;
  wire tmp33860;
  wire tmp33861;
  wire tmp33862;
  wire tmp33863;
  wire tmp33864;
  wire tmp33865;
  wire tmp33866;
  wire tmp33867;
  wire tmp33868;
  wire tmp33869;
  wire tmp33870;
  wire tmp33871;
  wire tmp33872;
  wire tmp33873;
  wire tmp33874;
  wire tmp33875;
  wire tmp33876;
  wire tmp33877;
  wire tmp33878;
  wire tmp33879;
  wire tmp33880;
  wire tmp33881;
  wire tmp33882;
  wire tmp33883;
  wire tmp33884;
  wire tmp33885;
  wire tmp33886;
  wire tmp33887;
  wire tmp33888;
  wire tmp33889;
  wire tmp33890;
  wire tmp33891;
  wire tmp33892;
  wire tmp33893;
  wire tmp33894;
  wire tmp33895;
  wire tmp33896;
  wire tmp33897;
  wire tmp33898;
  wire tmp33899;
  wire tmp33900;
  wire tmp33901;
  wire tmp33902;
  wire tmp33903;
  wire tmp33904;
  wire tmp33905;
  wire tmp33906;
  wire tmp33907;
  wire tmp33908;
  wire tmp33909;
  wire tmp33910;
  wire tmp33911;
  wire tmp33912;
  wire tmp33913;
  wire tmp33914;
  wire tmp33915;
  wire tmp33916;
  wire tmp33917;
  wire tmp33918;
  wire tmp33919;
  wire tmp33920;
  wire tmp33921;
  wire tmp33922;
  wire tmp33923;
  wire tmp33924;
  wire tmp33925;
  wire tmp33926;
  wire tmp33927;
  wire tmp33928;
  wire tmp33929;
  wire tmp33930;
  wire tmp33931;
  wire tmp33932;
  wire tmp33933;
  wire tmp33934;
  wire tmp33935;
  wire tmp33936;
  wire tmp33937;
  wire tmp33938;
  wire tmp33939;
  wire tmp33940;
  wire tmp33941;
  wire tmp33942;
  wire tmp33943;
  wire tmp33944;
  wire tmp33945;
  wire tmp33946;
  wire tmp33947;
  wire tmp33948;
  wire tmp33949;
  wire tmp33950;
  wire tmp33951;
  wire tmp33952;
  wire tmp33953;
  wire tmp33954;
  wire tmp33955;
  wire tmp33956;
  wire tmp33957;
  wire tmp33958;
  wire tmp33959;
  wire tmp33960;
  wire tmp33961;
  wire tmp33962;
  wire tmp33963;
  wire tmp33964;
  wire tmp33965;
  wire tmp33966;
  wire tmp33967;
  wire tmp33968;
  wire tmp33969;
  wire tmp33970;
  wire tmp33971;
  wire tmp33972;
  wire tmp33973;
  wire tmp33974;
  wire tmp33975;
  wire tmp33976;
  wire tmp33977;
  wire tmp33978;
  wire tmp33979;
  wire tmp33980;
  wire tmp33981;
  wire tmp33982;
  wire tmp33983;
  wire tmp33984;
  wire tmp33985;
  wire tmp33986;
  wire tmp33987;
  wire tmp33988;
  wire tmp33989;
  wire tmp33990;
  wire tmp33991;
  wire tmp33992;
  wire tmp33993;
  wire tmp33994;
  wire tmp33995;
  wire tmp33996;
  wire tmp33997;
  wire tmp33998;
  wire tmp33999;
  wire tmp34000;
  wire tmp34001;
  wire tmp34002;
  wire tmp34003;
  wire tmp34004;
  wire tmp34005;
  wire tmp34006;
  wire tmp34007;
  wire tmp34008;
  wire tmp34009;
  wire tmp34010;
  wire tmp34011;
  wire tmp34012;
  wire tmp34013;
  wire tmp34014;
  wire tmp34015;
  wire tmp34016;
  wire tmp34017;
  wire tmp34018;
  wire tmp34019;
  wire tmp34020;
  wire tmp34021;
  wire tmp34022;
  wire tmp34023;
  wire tmp34024;
  wire tmp34025;
  wire tmp34026;
  wire tmp34027;
  wire tmp34028;
  wire tmp34029;
  wire tmp34030;
  wire tmp34031;
  wire tmp34032;
  wire tmp34033;
  wire tmp34034;
  wire tmp34035;
  wire tmp34036;
  wire tmp34037;
  wire tmp34038;
  wire tmp34039;
  wire tmp34040;
  wire tmp34041;
  wire tmp34042;
  wire tmp34043;
  wire tmp34044;
  wire tmp34045;
  wire tmp34046;
  wire tmp34047;
  wire tmp34048;
  wire tmp34049;
  wire tmp34050;
  wire tmp34051;
  wire tmp34052;
  wire tmp34053;
  wire tmp34054;
  wire tmp34055;
  wire tmp34056;
  wire tmp34057;
  wire tmp34058;
  wire tmp34059;
  wire tmp34060;
  wire tmp34061;
  wire tmp34062;
  wire tmp34063;
  wire tmp34064;
  wire tmp34065;
  wire tmp34066;
  wire tmp34067;
  wire tmp34068;
  wire tmp34069;
  wire tmp34070;
  wire tmp34071;
  wire tmp34072;
  wire tmp34073;
  wire tmp34074;
  wire tmp34075;
  wire tmp34076;
  wire tmp34077;
  wire tmp34078;
  wire tmp34079;
  wire tmp34080;
  wire tmp34081;
  wire tmp34082;
  wire tmp34083;
  wire tmp34084;
  wire tmp34085;
  wire tmp34086;
  wire tmp34087;
  wire tmp34088;
  wire tmp34089;
  wire tmp34090;
  wire tmp34091;
  wire tmp34092;
  wire tmp34093;
  wire tmp34094;
  wire tmp34095;
  wire tmp34096;
  wire tmp34097;
  wire tmp34098;
  wire tmp34099;
  wire tmp34100;
  wire tmp34101;
  wire tmp34102;
  wire tmp34103;
  wire tmp34104;
  wire tmp34105;
  wire tmp34106;
  wire tmp34107;
  wire tmp34108;
  wire tmp34109;
  wire tmp34110;
  wire tmp34111;
  wire tmp34112;
  wire tmp34113;
  wire tmp34114;
  wire tmp34115;
  wire tmp34116;
  wire tmp34117;
  wire tmp34118;
  wire tmp34119;
  wire tmp34120;
  wire tmp34121;
  wire tmp34122;
  wire tmp34123;
  wire tmp34124;
  wire tmp34125;
  wire tmp34126;
  wire tmp34127;
  wire tmp34128;
  wire tmp34129;
  wire tmp34130;
  wire tmp34131;
  wire tmp34132;
  wire tmp34133;
  wire tmp34134;
  wire tmp34135;
  wire tmp34136;
  wire tmp34137;
  wire tmp34138;
  wire tmp34139;
  wire tmp34140;
  wire tmp34141;
  wire tmp34142;
  wire tmp34143;
  wire tmp34144;
  wire tmp34145;
  wire tmp34146;
  wire tmp34147;
  wire tmp34148;
  wire tmp34149;
  wire tmp34150;
  wire tmp34151;
  wire tmp34152;
  wire tmp34153;
  wire tmp34154;
  wire tmp34155;
  wire tmp34156;
  wire tmp34157;
  wire tmp34158;
  wire tmp34159;
  wire tmp34160;
  wire tmp34161;
  wire tmp34162;
  wire tmp34163;
  wire tmp34164;
  wire tmp34165;
  wire tmp34166;
  wire tmp34167;
  wire tmp34168;
  wire tmp34169;
  wire tmp34170;
  wire tmp34171;
  wire tmp34172;
  wire tmp34173;
  wire tmp34174;
  wire tmp34175;
  wire tmp34176;
  wire tmp34177;
  wire tmp34178;
  wire tmp34179;
  wire tmp34180;
  wire tmp34181;
  wire tmp34182;
  wire tmp34183;
  wire tmp34184;
  wire tmp34185;
  wire tmp34186;
  wire tmp34187;
  wire tmp34188;
  wire tmp34189;
  wire tmp34190;
  wire tmp34191;
  wire tmp34192;
  wire tmp34193;
  wire tmp34194;
  wire tmp34195;
  wire tmp34196;
  wire tmp34197;
  wire tmp34198;
  wire tmp34199;
  wire tmp34200;
  wire tmp34201;
  wire tmp34202;
  wire tmp34203;
  wire tmp34204;
  wire tmp34205;
  wire tmp34206;
  wire tmp34207;
  wire tmp34208;
  wire tmp34209;
  wire tmp34210;
  wire tmp34211;
  wire tmp34212;
  wire tmp34213;
  wire tmp34214;
  wire tmp34215;
  wire tmp34216;
  wire tmp34217;
  wire tmp34218;
  wire tmp34219;
  wire tmp34220;
  wire tmp34221;
  wire tmp34222;
  wire tmp34223;
  wire tmp34224;
  wire tmp34225;
  wire tmp34226;
  wire tmp34227;
  wire tmp34228;
  wire tmp34229;
  wire tmp34230;
  wire tmp34231;
  wire tmp34232;
  wire tmp34233;
  wire tmp34234;
  wire tmp34235;
  wire tmp34236;
  wire tmp34237;
  wire tmp34238;
  wire tmp34239;
  wire tmp34240;
  wire tmp34241;
  wire tmp34242;
  wire tmp34243;
  wire tmp34244;
  wire tmp34245;
  wire tmp34246;
  wire tmp34247;
  wire tmp34248;
  wire tmp34249;
  wire tmp34250;
  wire tmp34251;
  wire tmp34252;
  wire tmp34253;
  wire tmp34254;
  wire tmp34255;
  wire tmp34256;
  wire tmp34257;
  wire tmp34258;
  wire tmp34259;
  wire tmp34260;
  wire tmp34261;
  wire tmp34262;
  wire tmp34263;
  wire tmp34264;
  wire tmp34265;
  wire tmp34266;
  wire tmp34267;
  wire tmp34268;
  wire tmp34269;
  wire tmp34270;
  wire tmp34271;
  wire tmp34272;
  wire tmp34273;
  wire tmp34274;
  wire tmp34275;
  wire tmp34276;
  wire tmp34277;
  wire tmp34278;
  wire tmp34279;
  wire tmp34280;
  wire tmp34281;
  wire tmp34282;
  wire tmp34283;
  wire tmp34284;
  wire tmp34285;
  wire tmp34286;
  wire tmp34287;
  wire tmp34288;
  wire tmp34289;
  wire tmp34290;
  wire tmp34291;
  wire tmp34292;
  wire tmp34293;
  wire tmp34294;
  wire tmp34295;
  wire tmp34296;
  wire tmp34297;
  wire tmp34298;
  wire tmp34299;
  wire tmp34300;
  wire tmp34301;
  wire tmp34302;
  wire tmp34303;
  wire tmp34304;
  wire tmp34305;
  wire tmp34306;
  wire tmp34307;
  wire tmp34308;
  wire tmp34309;
  wire tmp34310;
  wire tmp34311;
  wire tmp34312;
  wire tmp34313;
  wire tmp34314;
  wire tmp34315;
  wire tmp34316;
  wire tmp34317;
  wire tmp34318;
  wire tmp34319;
  wire tmp34320;
  wire tmp34321;
  wire tmp34322;
  wire tmp34323;
  wire tmp34324;
  wire tmp34325;
  wire tmp34326;
  wire tmp34327;
  wire tmp34328;
  wire tmp34329;
  wire tmp34330;
  wire tmp34331;
  wire tmp34332;
  wire tmp34333;
  wire tmp34334;
  wire tmp34335;
  wire tmp34336;
  wire tmp34337;
  wire tmp34338;
  wire tmp34339;
  wire tmp34340;
  wire tmp34341;
  wire tmp34342;
  wire tmp34343;
  wire tmp34344;
  wire tmp34345;
  wire tmp34346;
  wire tmp34347;
  wire tmp34348;
  wire tmp34349;
  wire tmp34350;
  wire tmp34351;
  wire tmp34352;
  wire tmp34353;
  wire tmp34354;
  wire tmp34355;
  wire tmp34356;
  wire tmp34357;
  wire tmp34358;
  wire tmp34359;
  wire tmp34360;
  wire tmp34361;
  wire tmp34362;
  wire tmp34363;
  wire tmp34364;
  wire tmp34365;
  wire tmp34366;
  wire tmp34367;
  wire tmp34368;
  wire tmp34369;
  wire tmp34370;
  wire tmp34371;
  wire tmp34372;
  wire tmp34373;
  wire tmp34374;
  wire tmp34375;
  wire tmp34376;
  wire tmp34377;
  wire tmp34378;
  wire tmp34379;
  wire tmp34380;
  wire tmp34381;
  wire tmp34382;
  wire tmp34383;
  wire tmp34384;
  wire tmp34385;
  wire tmp34386;
  wire tmp34387;
  wire tmp34388;
  wire tmp34389;
  wire tmp34390;
  wire tmp34391;
  wire tmp34392;
  wire tmp34393;
  wire tmp34394;
  wire tmp34395;
  wire tmp34396;
  wire tmp34397;
  wire tmp34398;
  wire tmp34399;
  wire tmp34400;
  wire tmp34401;
  wire tmp34402;
  wire tmp34403;
  wire tmp34404;
  wire tmp34405;
  wire tmp34406;
  wire tmp34407;
  wire tmp34408;
  wire tmp34409;
  wire tmp34410;
  wire tmp34411;
  wire tmp34412;
  wire tmp34413;
  wire tmp34414;
  wire tmp34415;
  wire tmp34416;
  wire tmp34417;
  wire tmp34418;
  wire tmp34419;
  wire tmp34420;
  wire tmp34421;
  wire tmp34422;
  wire tmp34423;
  wire tmp34424;
  wire tmp34425;
  wire tmp34426;
  wire tmp34427;
  wire tmp34428;
  wire tmp34429;
  wire tmp34430;
  wire tmp34431;
  wire tmp34432;
  wire tmp34433;
  wire tmp34434;
  wire tmp34435;
  wire tmp34436;
  wire tmp34437;
  wire tmp34438;
  wire tmp34439;
  wire tmp34440;
  wire tmp34441;
  wire tmp34442;
  wire tmp34443;
  wire tmp34444;
  wire tmp34445;
  wire tmp34446;
  wire tmp34447;
  wire tmp34448;
  wire tmp34449;
  wire tmp34450;
  wire tmp34451;
  wire tmp34452;
  wire tmp34453;
  wire tmp34454;
  wire tmp34455;
  wire tmp34456;
  wire tmp34457;
  wire tmp34458;
  wire tmp34459;
  wire tmp34460;
  wire tmp34461;
  wire tmp34462;
  wire tmp34463;
  wire tmp34464;
  wire tmp34465;
  wire tmp34466;
  wire tmp34467;
  wire tmp34468;
  wire tmp34469;
  wire tmp34470;
  wire tmp34471;
  wire tmp34472;
  wire tmp34473;
  wire tmp34474;
  wire tmp34475;
  wire tmp34476;
  wire tmp34477;
  wire tmp34478;
  wire tmp34479;
  wire tmp34480;
  wire tmp34481;
  wire tmp34482;
  wire tmp34483;
  wire tmp34484;
  wire tmp34485;
  wire tmp34486;
  wire tmp34487;
  wire tmp34488;
  wire tmp34489;
  wire tmp34490;
  wire tmp34491;
  wire tmp34492;
  wire tmp34493;
  wire tmp34494;
  wire tmp34495;
  wire tmp34496;
  wire tmp34497;
  wire tmp34498;
  wire tmp34499;
  wire tmp34500;
  wire tmp34501;
  wire tmp34502;
  wire tmp34503;
  wire tmp34504;
  wire tmp34505;
  wire tmp34506;
  wire tmp34507;
  wire tmp34508;
  wire tmp34509;
  wire tmp34510;
  wire tmp34511;
  wire tmp34512;
  wire tmp34513;
  wire tmp34514;
  wire tmp34515;
  wire tmp34516;
  wire tmp34517;
  wire tmp34518;
  wire tmp34519;
  wire tmp34520;
  wire tmp34521;
  wire tmp34522;
  wire tmp34523;
  wire tmp34524;
  wire tmp34525;
  wire tmp34526;
  wire tmp34527;
  wire tmp34528;
  wire tmp34529;
  wire tmp34530;
  wire tmp34531;
  wire tmp34532;
  wire tmp34533;
  wire tmp34534;
  wire tmp34535;
  wire tmp34536;
  wire tmp34537;
  wire tmp34538;
  wire tmp34539;
  wire tmp34540;
  wire tmp34541;
  wire tmp34542;
  wire tmp34543;
  wire tmp34544;
  wire tmp34545;
  wire tmp34546;
  wire tmp34547;
  wire tmp34548;
  wire tmp34549;
  wire tmp34550;
  wire tmp34551;
  wire tmp34552;
  wire tmp34553;
  wire tmp34554;
  wire tmp34555;
  wire tmp34556;
  wire tmp34557;
  wire tmp34558;
  wire tmp34559;
  wire tmp34560;
  wire tmp34561;
  wire tmp34562;
  wire tmp34563;
  wire tmp34564;
  wire tmp34565;
  wire tmp34566;
  wire tmp34567;
  wire tmp34568;
  wire tmp34569;
  wire tmp34570;
  wire tmp34571;
  wire tmp34572;
  wire tmp34573;
  wire tmp34574;
  wire tmp34575;
  wire tmp34576;
  wire tmp34577;
  wire tmp34578;
  wire tmp34579;
  wire tmp34580;
  wire tmp34581;
  wire tmp34582;
  wire tmp34583;
  wire tmp34584;
  wire tmp34585;
  wire tmp34586;
  wire tmp34587;
  wire tmp34588;
  wire tmp34589;
  wire tmp34590;
  wire tmp34591;
  wire tmp34592;
  wire tmp34593;
  wire tmp34594;
  wire tmp34595;
  wire tmp34596;
  wire tmp34597;
  wire tmp34598;
  wire tmp34599;
  wire tmp34600;
  wire tmp34601;
  wire tmp34602;
  wire tmp34603;
  wire tmp34604;
  wire tmp34605;
  wire tmp34606;
  wire tmp34607;
  wire tmp34608;
  wire tmp34609;
  wire tmp34610;
  wire tmp34611;
  wire tmp34612;
  wire tmp34613;
  wire tmp34614;
  wire tmp34615;
  wire tmp34616;
  wire tmp34617;
  wire tmp34618;
  wire tmp34619;
  wire tmp34620;
  wire tmp34621;
  wire tmp34622;
  wire tmp34623;
  wire tmp34624;
  wire tmp34625;
  wire tmp34626;
  wire tmp34627;
  wire tmp34628;
  wire tmp34629;
  wire tmp34630;
  wire tmp34631;
  wire tmp34632;
  wire tmp34633;
  wire tmp34634;
  wire tmp34635;
  wire tmp34636;
  wire tmp34637;
  wire tmp34638;
  wire tmp34639;
  wire tmp34640;
  wire tmp34641;
  wire tmp34642;
  wire tmp34643;
  wire tmp34644;
  wire tmp34645;
  wire tmp34646;
  wire tmp34647;
  wire tmp34648;
  wire tmp34649;
  wire tmp34650;
  wire tmp34651;
  wire tmp34652;
  wire tmp34653;
  wire tmp34654;
  wire tmp34655;
  wire tmp34656;
  wire tmp34657;
  wire tmp34658;
  wire tmp34659;
  wire tmp34660;
  wire tmp34661;
  wire tmp34662;
  wire tmp34663;
  wire tmp34664;
  wire tmp34665;
  wire tmp34666;
  wire tmp34667;
  wire tmp34668;
  wire tmp34669;
  wire tmp34670;
  wire tmp34671;
  wire tmp34672;
  wire tmp34673;
  wire tmp34674;
  wire tmp34675;
  wire tmp34676;
  wire tmp34677;
  wire tmp34678;
  wire tmp34679;
  wire tmp34680;
  wire tmp34681;
  wire tmp34682;
  wire tmp34683;
  wire tmp34684;
  wire tmp34685;
  wire tmp34686;
  wire tmp34687;
  wire tmp34688;
  wire tmp34689;
  wire tmp34690;
  wire tmp34691;
  wire tmp34692;
  wire tmp34693;
  wire tmp34694;
  wire tmp34695;
  wire tmp34696;
  wire tmp34697;
  wire tmp34698;
  wire tmp34699;
  wire tmp34700;
  wire tmp34701;
  wire tmp34702;
  wire tmp34703;
  wire tmp34704;
  wire tmp34705;
  wire tmp34706;
  wire tmp34707;
  wire tmp34708;
  wire tmp34709;
  wire tmp34710;
  wire tmp34711;
  wire tmp34712;
  wire tmp34713;
  wire tmp34714;
  wire tmp34715;
  wire tmp34716;
  wire tmp34717;
  wire tmp34718;
  wire tmp34719;
  wire tmp34720;
  wire tmp34721;
  wire tmp34722;
  wire tmp34723;
  wire tmp34724;
  wire tmp34725;
  wire tmp34726;
  wire tmp34727;
  wire tmp34728;
  wire tmp34729;
  wire tmp34730;
  wire tmp34731;
  wire tmp34732;
  wire tmp34733;
  wire tmp34734;
  wire tmp34735;
  wire tmp34736;
  wire tmp34737;
  wire tmp34738;
  wire tmp34739;
  wire tmp34740;
  wire tmp34741;
  wire tmp34742;
  wire tmp34743;
  wire tmp34744;
  wire tmp34745;
  wire tmp34746;
  wire tmp34747;
  wire tmp34748;
  wire tmp34749;
  wire tmp34750;
  wire tmp34751;
  wire tmp34752;
  wire tmp34753;
  wire tmp34754;
  wire tmp34755;
  wire tmp34756;
  wire tmp34757;
  wire tmp34758;
  wire tmp34759;
  wire tmp34760;
  wire tmp34761;
  wire tmp34762;
  wire tmp34763;
  wire tmp34764;
  wire tmp34765;
  wire tmp34766;
  wire tmp34767;
  wire tmp34768;
  wire tmp34769;
  wire tmp34770;
  wire tmp34771;
  wire tmp34772;
  wire tmp34773;
  wire tmp34774;
  wire tmp34775;
  wire tmp34776;
  wire tmp34777;
  wire tmp34778;
  wire tmp34779;
  wire tmp34780;
  wire tmp34781;
  wire tmp34782;
  wire tmp34783;
  wire tmp34784;
  wire tmp34785;
  wire tmp34786;
  wire tmp34787;
  wire tmp34788;
  wire tmp34789;
  wire tmp34790;
  wire tmp34791;
  wire tmp34792;
  wire tmp34793;
  wire tmp34794;
  wire tmp34795;
  wire tmp34796;
  wire tmp34797;
  wire tmp34798;
  wire tmp34799;
  wire tmp34800;
  wire tmp34801;
  wire tmp34802;
  wire tmp34803;
  wire tmp34804;
  wire tmp34805;
  wire tmp34806;
  wire tmp34807;
  wire tmp34808;
  wire tmp34809;
  wire tmp34810;
  wire tmp34811;
  wire tmp34812;
  wire tmp34813;
  wire tmp34814;
  wire tmp34815;
  wire tmp34816;
  wire tmp34817;
  wire tmp34818;
  wire tmp34819;
  wire tmp34820;
  wire tmp34821;
  wire tmp34822;
  wire tmp34823;
  wire tmp34824;
  wire tmp34825;
  wire tmp34826;
  wire tmp34827;
  wire tmp34828;
  wire tmp34829;
  wire tmp34830;
  wire tmp34831;
  wire tmp34832;
  wire tmp34833;
  wire tmp34834;
  wire tmp34835;
  wire tmp34836;
  wire tmp34837;
  wire tmp34838;
  wire tmp34839;
  wire tmp34840;
  wire tmp34841;
  wire tmp34842;
  wire tmp34843;
  wire tmp34844;
  wire tmp34845;
  wire tmp34846;
  wire tmp34847;
  wire tmp34848;
  wire tmp34849;
  wire tmp34850;
  wire tmp34851;
  wire tmp34852;
  wire tmp34853;
  wire tmp34854;
  wire tmp34855;
  wire tmp34856;
  wire tmp34857;
  wire tmp34858;
  wire tmp34859;
  wire tmp34860;
  wire tmp34861;
  wire tmp34862;
  wire tmp34863;
  wire tmp34864;
  wire tmp34865;
  wire tmp34866;
  wire tmp34867;
  wire tmp34868;
  wire tmp34869;
  wire tmp34870;
  wire tmp34871;
  wire tmp34872;
  wire tmp34873;
  wire tmp34874;
  wire tmp34875;
  wire tmp34876;
  wire tmp34877;
  wire tmp34878;
  wire tmp34879;
  wire tmp34880;
  wire tmp34881;
  wire tmp34882;
  wire tmp34883;
  wire tmp34884;
  wire tmp34885;
  wire tmp34886;
  wire tmp34887;
  wire tmp34888;
  wire tmp34889;
  wire tmp34890;
  wire tmp34891;
  wire tmp34892;
  wire tmp34893;
  wire tmp34894;
  wire tmp34895;
  wire tmp34896;
  wire tmp34897;
  wire tmp34898;
  wire tmp34899;
  wire tmp34900;
  wire tmp34901;
  wire tmp34902;
  wire tmp34903;
  wire tmp34904;
  wire tmp34905;
  wire tmp34906;
  wire tmp34907;
  wire tmp34908;
  wire tmp34909;
  wire tmp34910;
  wire tmp34911;
  wire tmp34912;
  wire tmp34913;
  wire tmp34914;
  wire tmp34915;
  wire tmp34916;
  wire tmp34917;
  wire tmp34918;
  wire tmp34919;
  wire tmp34920;
  wire tmp34921;
  wire tmp34922;
  wire tmp34923;
  wire tmp34924;
  wire tmp34925;
  wire tmp34926;
  wire tmp34927;
  wire tmp34928;
  wire tmp34929;
  wire tmp34930;
  wire tmp34931;
  wire tmp34932;
  wire tmp34933;
  wire tmp34934;
  wire tmp34935;
  wire tmp34936;
  wire tmp34937;
  wire tmp34938;
  wire tmp34939;
  wire tmp34940;
  wire tmp34941;
  wire tmp34942;
  wire tmp34943;
  wire tmp34944;
  wire tmp34945;
  wire tmp34946;
  wire tmp34947;
  wire tmp34948;
  wire tmp34949;
  wire tmp34950;
  wire tmp34951;
  wire tmp34952;
  wire tmp34953;
  wire tmp34954;
  wire tmp34955;
  wire tmp34956;
  wire tmp34957;
  wire tmp34958;
  wire tmp34959;
  wire tmp34960;
  wire tmp34961;
  wire tmp34962;
  wire tmp34963;
  wire tmp34964;
  wire tmp34965;
  wire tmp34966;
  wire tmp34967;
  wire tmp34968;
  wire tmp34969;
  wire tmp34970;
  wire tmp34971;
  wire tmp34972;
  wire tmp34973;
  wire tmp34974;
  wire tmp34975;
  wire tmp34976;
  wire tmp34977;
  wire tmp34978;
  wire tmp34979;
  wire tmp34980;
  wire tmp34981;
  wire tmp34982;
  wire tmp34983;
  wire tmp34984;
  wire tmp34985;
  wire tmp34986;
  wire tmp34987;
  wire tmp34988;
  wire tmp34989;
  wire tmp34990;
  wire tmp34991;
  wire tmp34992;
  wire tmp34993;
  wire tmp34994;
  wire tmp34995;
  wire tmp34996;
  wire tmp34997;
  wire tmp34998;
  wire tmp34999;
  wire tmp35000;
  wire tmp35001;
  wire tmp35002;
  wire tmp35003;
  wire tmp35004;
  wire tmp35005;
  wire tmp35006;
  wire tmp35007;
  wire tmp35008;
  wire tmp35009;
  wire tmp35010;
  wire tmp35011;
  wire tmp35012;
  wire tmp35013;
  wire tmp35014;
  wire tmp35015;
  wire tmp35016;
  wire tmp35017;
  wire tmp35018;
  wire tmp35019;
  wire tmp35020;
  wire tmp35021;
  wire tmp35022;
  wire tmp35023;
  wire tmp35024;
  wire tmp35025;
  wire tmp35026;
  wire tmp35027;
  wire tmp35028;
  wire tmp35029;
  wire tmp35030;
  wire tmp35031;
  wire tmp35032;
  wire tmp35033;
  wire tmp35034;
  wire tmp35035;
  wire tmp35036;
  wire tmp35037;
  wire tmp35038;
  wire tmp35039;
  wire tmp35040;
  wire tmp35041;
  wire tmp35042;
  wire tmp35043;
  wire tmp35044;
  wire tmp35045;
  wire tmp35046;
  wire tmp35047;
  wire tmp35048;
  wire tmp35049;
  wire tmp35050;
  wire tmp35051;
  wire tmp35052;
  wire tmp35053;
  wire tmp35054;
  wire tmp35055;
  wire tmp35056;
  wire tmp35057;
  wire tmp35058;
  wire tmp35059;
  wire tmp35060;
  wire tmp35061;
  wire tmp35062;
  wire tmp35063;
  wire tmp35064;
  wire tmp35065;
  wire tmp35066;
  wire tmp35067;
  wire tmp35068;
  wire tmp35069;
  wire tmp35070;
  wire tmp35071;
  wire tmp35072;
  wire tmp35073;
  wire tmp35074;
  wire tmp35075;
  wire tmp35076;
  wire tmp35077;
  wire tmp35078;
  wire tmp35079;
  wire tmp35080;
  wire tmp35081;
  wire tmp35082;
  wire tmp35083;
  wire tmp35084;
  wire tmp35085;
  wire tmp35086;
  wire tmp35087;
  wire tmp35088;
  wire tmp35089;
  wire tmp35090;
  wire tmp35091;
  wire tmp35092;
  wire tmp35093;
  wire tmp35094;
  wire tmp35095;
  wire tmp35096;
  wire tmp35097;
  wire tmp35098;
  wire tmp35099;
  wire tmp35100;
  wire tmp35101;
  wire tmp35102;
  wire tmp35103;
  wire tmp35104;
  wire tmp35105;
  wire tmp35106;
  wire tmp35107;
  wire tmp35108;
  wire tmp35109;
  wire tmp35110;
  wire tmp35111;
  wire tmp35112;
  wire tmp35113;
  wire tmp35114;
  wire tmp35115;
  wire tmp35116;
  wire tmp35117;
  wire tmp35118;
  wire tmp35119;
  wire tmp35120;
  wire tmp35121;
  wire tmp35122;
  wire tmp35123;
  wire tmp35124;
  wire tmp35125;
  wire tmp35126;
  wire tmp35127;
  wire tmp35128;
  wire tmp35129;
  wire tmp35130;
  wire tmp35131;
  wire tmp35132;
  wire tmp35133;
  wire tmp35134;
  wire tmp35135;
  wire tmp35136;
  wire tmp35137;
  wire tmp35138;
  wire tmp35139;
  wire tmp35140;
  wire tmp35141;
  wire tmp35142;
  wire tmp35143;
  wire tmp35144;
  wire tmp35145;
  wire tmp35146;
  wire tmp35147;
  wire tmp35148;
  wire tmp35149;
  wire tmp35150;
  wire tmp35151;
  wire tmp35152;
  wire tmp35153;
  wire tmp35154;
  wire tmp35155;
  wire tmp35156;
  wire tmp35157;
  wire tmp35158;
  wire tmp35159;
  wire tmp35160;
  wire tmp35161;
  wire tmp35162;
  wire tmp35163;
  wire tmp35164;
  wire tmp35165;
  wire tmp35166;
  wire tmp35167;
  wire tmp35168;
  wire tmp35169;
  wire tmp35170;
  wire tmp35171;
  wire tmp35172;
  wire tmp35173;
  wire tmp35174;
  wire tmp35175;
  wire tmp35176;
  wire tmp35177;
  wire tmp35178;
  wire tmp35179;
  wire tmp35180;
  wire tmp35181;
  wire tmp35182;
  wire tmp35183;
  wire tmp35184;
  wire tmp35185;
  wire tmp35186;
  wire tmp35187;
  wire tmp35188;
  wire tmp35189;
  wire tmp35190;
  wire tmp35191;
  wire tmp35192;
  wire tmp35193;
  wire tmp35194;
  wire tmp35195;
  wire tmp35196;
  wire tmp35197;
  wire tmp35198;
  wire tmp35199;
  wire tmp35200;
  wire tmp35201;
  wire tmp35202;
  wire tmp35203;
  wire tmp35204;
  wire tmp35205;
  wire tmp35206;
  wire tmp35207;
  wire tmp35208;
  wire tmp35209;
  wire tmp35210;
  wire tmp35211;
  wire tmp35212;
  wire tmp35213;
  wire tmp35214;
  wire tmp35215;
  wire tmp35216;
  wire tmp35217;
  wire tmp35218;
  wire tmp35219;
  wire tmp35220;
  wire tmp35221;
  wire tmp35222;
  wire tmp35223;
  wire tmp35224;
  wire tmp35225;
  wire tmp35226;
  wire tmp35227;
  wire tmp35228;
  wire tmp35229;
  wire tmp35230;
  wire tmp35231;
  wire tmp35232;
  wire tmp35233;
  wire tmp35234;
  wire tmp35235;
  wire tmp35236;
  wire tmp35237;
  wire tmp35238;
  wire tmp35239;
  wire tmp35240;
  wire tmp35241;
  wire tmp35242;
  wire tmp35243;
  wire tmp35244;
  wire tmp35245;
  wire tmp35246;
  wire tmp35247;
  wire tmp35248;
  wire tmp35249;
  wire tmp35250;
  wire tmp35251;
  wire tmp35252;
  wire tmp35253;
  wire tmp35254;
  wire tmp35255;
  wire tmp35256;
  wire tmp35257;
  wire tmp35258;
  wire tmp35259;
  wire tmp35260;
  wire tmp35261;
  wire tmp35262;
  wire tmp35263;
  wire tmp35264;
  wire tmp35265;
  wire tmp35266;
  wire tmp35267;
  wire tmp35268;
  wire tmp35269;
  wire tmp35270;
  wire tmp35271;
  wire tmp35272;
  wire tmp35273;
  wire tmp35274;
  wire tmp35275;
  wire tmp35276;
  wire tmp35277;
  wire tmp35278;
  wire tmp35279;
  wire tmp35280;
  wire tmp35281;
  wire tmp35282;
  wire tmp35283;
  wire tmp35284;
  wire tmp35285;
  wire tmp35286;
  wire tmp35287;
  wire tmp35288;
  wire tmp35289;
  wire tmp35290;
  wire tmp35291;
  wire tmp35292;
  wire tmp35293;
  wire tmp35294;
  wire tmp35295;
  wire tmp35296;
  wire tmp35297;
  wire tmp35298;
  wire tmp35299;
  wire tmp35300;
  wire tmp35301;
  wire tmp35302;
  wire tmp35303;
  wire tmp35304;
  wire tmp35305;
  wire tmp35306;
  wire tmp35307;
  wire tmp35308;
  wire tmp35309;
  wire tmp35310;
  wire tmp35311;
  wire tmp35312;
  wire tmp35313;
  wire tmp35314;
  wire tmp35315;
  wire tmp35316;
  wire tmp35317;
  wire tmp35318;
  wire tmp35319;
  wire tmp35320;
  wire tmp35321;
  wire tmp35322;
  wire tmp35323;
  wire tmp35324;
  wire tmp35325;
  wire tmp35326;
  wire tmp35327;
  wire tmp35328;
  wire tmp35329;
  wire tmp35330;
  wire tmp35331;
  wire tmp35332;
  wire tmp35333;
  wire tmp35334;
  wire tmp35335;
  wire tmp35336;
  wire tmp35337;
  wire tmp35338;
  wire tmp35339;
  wire tmp35340;
  wire tmp35341;
  wire tmp35342;
  wire tmp35343;
  wire tmp35344;
  wire tmp35345;
  wire tmp35346;
  wire tmp35347;
  wire tmp35348;
  wire tmp35349;
  wire tmp35350;
  wire tmp35351;
  wire tmp35352;
  wire tmp35353;
  wire tmp35354;
  wire tmp35355;
  wire tmp35356;
  wire tmp35357;
  wire tmp35358;
  wire tmp35359;
  wire tmp35360;
  wire tmp35361;
  wire tmp35362;
  wire tmp35363;
  wire tmp35364;
  wire tmp35365;
  wire tmp35366;
  wire tmp35367;
  wire tmp35368;
  wire tmp35369;
  wire tmp35370;
  wire tmp35371;
  wire tmp35372;
  wire tmp35373;
  wire tmp35374;
  wire tmp35375;
  wire tmp35376;
  wire tmp35377;
  wire tmp35378;
  wire tmp35379;
  wire tmp35380;
  wire tmp35381;
  wire tmp35382;
  wire tmp35383;
  wire tmp35384;
  wire tmp35385;
  wire tmp35386;
  wire tmp35387;
  wire tmp35388;
  wire tmp35389;
  wire tmp35390;
  wire tmp35391;
  wire tmp35392;
  wire tmp35393;
  wire tmp35394;
  wire tmp35395;
  wire tmp35396;
  wire tmp35397;
  wire tmp35398;
  wire tmp35399;
  wire tmp35400;
  wire tmp35401;
  wire tmp35402;
  wire tmp35403;
  wire tmp35404;
  wire tmp35405;
  wire tmp35406;
  wire tmp35407;
  wire tmp35408;
  wire tmp35409;
  wire tmp35410;
  wire tmp35411;
  wire tmp35412;
  wire tmp35413;
  wire tmp35414;
  wire tmp35415;
  wire tmp35416;
  wire tmp35417;
  wire tmp35418;
  wire tmp35419;
  wire tmp35420;
  wire tmp35421;
  wire tmp35422;
  wire tmp35423;
  wire tmp35424;
  wire tmp35425;
  wire tmp35426;
  wire tmp35427;
  wire tmp35428;
  wire tmp35429;
  wire tmp35430;
  wire tmp35431;
  wire tmp35432;
  wire tmp35433;
  wire tmp35434;
  wire tmp35435;
  wire tmp35436;
  wire tmp35437;
  wire tmp35438;
  wire tmp35439;
  wire tmp35440;
  wire tmp35441;
  wire tmp35442;
  wire tmp35443;
  wire tmp35444;
  wire tmp35445;
  wire tmp35446;
  wire tmp35447;
  wire tmp35448;
  wire tmp35449;
  wire tmp35450;
  wire tmp35451;
  wire tmp35452;
  wire tmp35453;
  wire tmp35454;
  wire tmp35455;
  wire tmp35456;
  wire tmp35457;
  wire tmp35458;
  wire tmp35459;
  wire tmp35460;
  wire tmp35461;
  wire tmp35462;
  wire tmp35463;
  wire tmp35464;
  wire tmp35465;
  wire tmp35466;
  wire tmp35467;
  wire tmp35468;
  wire tmp35469;
  wire tmp35470;
  wire tmp35471;
  wire tmp35472;
  wire tmp35473;
  wire tmp35474;
  wire tmp35475;
  wire tmp35476;
  wire tmp35477;
  wire tmp35478;
  wire tmp35479;
  wire tmp35480;
  wire tmp35481;
  wire tmp35482;
  wire tmp35483;
  wire tmp35484;
  wire tmp35485;
  wire tmp35486;
  wire tmp35487;
  wire tmp35488;
  wire tmp35489;
  wire tmp35490;
  wire tmp35491;
  wire tmp35492;
  wire tmp35493;
  wire tmp35494;
  wire tmp35495;
  wire tmp35496;
  wire tmp35497;
  wire tmp35498;
  wire tmp35499;
  wire tmp35500;
  wire tmp35501;
  wire tmp35502;
  wire tmp35503;
  wire tmp35504;
  wire tmp35505;
  wire tmp35506;
  wire tmp35507;
  wire tmp35508;
  wire tmp35509;
  wire tmp35510;
  wire tmp35511;
  wire tmp35512;
  wire tmp35513;
  wire tmp35514;
  wire tmp35515;
  wire tmp35516;
  wire tmp35517;
  wire tmp35518;
  wire tmp35519;
  wire tmp35520;
  wire tmp35521;
  wire tmp35522;
  wire tmp35523;
  wire tmp35524;
  wire tmp35525;
  wire tmp35526;
  wire tmp35527;
  wire tmp35528;
  wire tmp35529;
  wire tmp35530;
  wire tmp35531;
  wire tmp35532;
  wire tmp35533;
  wire tmp35534;
  wire tmp35535;
  wire tmp35536;
  wire tmp35537;
  wire tmp35538;
  wire tmp35539;
  wire tmp35540;
  wire tmp35541;
  wire tmp35542;
  wire tmp35543;
  wire tmp35544;
  wire tmp35545;
  wire tmp35546;
  wire tmp35547;
  wire tmp35548;
  wire tmp35549;
  wire tmp35550;
  wire tmp35551;
  wire tmp35552;
  wire tmp35553;
  wire tmp35554;
  wire tmp35555;
  wire tmp35556;
  wire tmp35557;
  wire tmp35558;
  wire tmp35559;
  wire tmp35560;
  wire tmp35561;
  wire tmp35562;
  wire tmp35563;
  wire tmp35564;
  wire tmp35565;
  wire tmp35566;
  wire tmp35567;
  wire tmp35568;
  wire tmp35569;
  wire tmp35570;
  wire tmp35571;
  wire tmp35572;
  wire tmp35573;
  wire tmp35574;
  wire tmp35575;
  wire tmp35576;
  wire tmp35577;
  wire tmp35578;
  wire tmp35579;
  wire tmp35580;
  wire tmp35581;
  wire tmp35582;
  wire tmp35583;
  wire tmp35584;
  wire tmp35585;
  wire tmp35586;
  wire tmp35587;
  wire tmp35588;
  wire tmp35589;
  wire tmp35590;
  wire tmp35591;
  wire tmp35592;
  wire tmp35593;
  wire tmp35594;
  wire tmp35595;
  wire tmp35596;
  wire tmp35597;
  wire tmp35598;
  wire tmp35599;
  wire tmp35600;
  wire tmp35601;
  wire tmp35602;
  wire tmp35603;
  wire tmp35604;
  wire tmp35605;
  wire tmp35606;
  wire tmp35607;
  wire tmp35608;
  wire tmp35609;
  wire tmp35610;
  wire tmp35611;
  wire tmp35612;
  wire tmp35613;
  wire tmp35614;
  wire tmp35615;
  wire tmp35616;
  wire tmp35617;
  wire tmp35618;
  wire tmp35619;
  wire tmp35620;
  wire tmp35621;
  wire tmp35622;
  wire tmp35623;
  wire tmp35624;
  wire tmp35625;
  wire tmp35626;
  wire tmp35627;
  wire tmp35628;
  wire tmp35629;
  wire tmp35630;
  wire tmp35631;
  wire tmp35632;
  wire tmp35633;
  wire tmp35634;
  wire tmp35635;
  wire tmp35636;
  wire tmp35637;
  wire tmp35638;
  wire tmp35639;
  wire tmp35640;
  wire tmp35641;
  wire tmp35642;
  wire tmp35643;
  wire tmp35644;
  wire tmp35645;
  wire tmp35646;
  wire tmp35647;
  wire tmp35648;
  wire tmp35649;
  wire tmp35650;
  wire tmp35651;
  wire tmp35652;
  wire tmp35653;
  wire tmp35654;
  wire tmp35655;
  wire tmp35656;
  wire tmp35657;
  wire tmp35658;
  wire tmp35659;
  wire tmp35660;
  wire tmp35661;
  wire tmp35662;
  wire tmp35663;
  wire tmp35664;
  wire tmp35665;
  wire tmp35666;
  wire tmp35667;
  wire tmp35668;
  wire tmp35669;
  wire tmp35670;
  wire tmp35671;
  wire tmp35672;
  wire tmp35673;
  wire tmp35674;
  wire tmp35675;
  wire tmp35676;
  wire tmp35677;
  wire tmp35678;
  wire tmp35679;
  wire tmp35680;
  wire tmp35681;
  wire tmp35682;
  wire tmp35683;
  wire tmp35684;
  wire tmp35685;
  wire tmp35686;
  wire tmp35687;
  wire tmp35688;
  wire tmp35689;
  wire tmp35690;
  wire tmp35691;
  wire tmp35692;
  wire tmp35693;
  wire tmp35694;
  wire tmp35695;
  wire tmp35696;
  wire tmp35697;
  wire tmp35698;
  wire tmp35699;
  wire tmp35700;
  wire tmp35701;
  wire tmp35702;
  wire tmp35703;
  wire tmp35704;
  wire tmp35705;
  wire tmp35706;
  wire tmp35707;
  wire tmp35708;
  wire tmp35709;
  wire tmp35710;
  wire tmp35711;
  wire tmp35712;
  wire tmp35713;
  wire tmp35714;
  wire tmp35715;
  wire tmp35716;
  wire tmp35717;
  wire tmp35718;
  wire tmp35719;
  wire tmp35720;
  wire tmp35721;
  wire tmp35722;
  wire tmp35723;
  wire tmp35724;
  wire tmp35725;
  wire tmp35726;
  wire tmp35727;
  wire tmp35728;
  wire tmp35729;
  wire tmp35730;
  wire tmp35731;
  wire tmp35732;
  wire tmp35733;
  wire tmp35734;
  wire tmp35735;
  wire tmp35736;
  wire tmp35737;
  wire tmp35738;
  wire tmp35739;
  wire tmp35740;
  wire tmp35741;
  wire tmp35742;
  wire tmp35743;
  wire tmp35744;
  wire tmp35745;
  wire tmp35746;
  wire tmp35747;
  wire tmp35748;
  wire tmp35749;
  wire tmp35750;
  wire tmp35751;
  wire tmp35752;
  wire tmp35753;
  wire tmp35754;
  wire tmp35755;
  wire tmp35756;
  wire tmp35757;
  wire tmp35758;
  wire tmp35759;
  wire tmp35760;
  wire tmp35761;
  wire tmp35762;
  wire tmp35763;
  wire tmp35764;
  wire tmp35765;
  wire tmp35766;
  wire tmp35767;
  wire tmp35768;
  wire tmp35769;
  wire tmp35770;
  wire tmp35771;
  wire tmp35772;
  wire tmp35773;
  wire tmp35774;
  wire tmp35775;
  wire tmp35776;
  wire tmp35777;
  wire tmp35778;
  wire tmp35779;
  wire tmp35780;
  wire tmp35781;
  wire tmp35782;
  wire tmp35783;
  wire tmp35784;
  wire tmp35785;
  wire tmp35786;
  wire tmp35787;
  wire tmp35788;
  wire tmp35789;
  wire tmp35790;
  wire tmp35791;
  wire tmp35792;
  wire tmp35793;
  wire tmp35794;
  wire tmp35795;
  wire tmp35796;
  wire tmp35797;
  wire tmp35798;
  wire tmp35799;
  wire tmp35800;
  wire tmp35801;
  wire tmp35802;
  wire tmp35803;
  wire tmp35804;
  wire tmp35805;
  wire tmp35806;
  wire tmp35807;
  wire tmp35808;
  wire tmp35809;
  wire tmp35810;
  wire tmp35811;
  wire tmp35812;
  wire tmp35813;
  wire tmp35814;
  wire tmp35815;
  wire tmp35816;
  wire tmp35817;
  wire tmp35818;
  wire tmp35819;
  wire tmp35820;
  wire tmp35821;
  wire tmp35822;
  wire tmp35823;
  wire tmp35824;
  wire tmp35825;
  wire tmp35826;
  wire tmp35827;
  wire tmp35828;
  wire tmp35829;
  wire tmp35830;
  wire tmp35831;
  wire tmp35832;
  wire tmp35833;
  wire tmp35834;
  wire tmp35835;
  wire tmp35836;
  wire tmp35837;
  wire tmp35838;
  wire tmp35839;
  wire tmp35840;
  wire tmp35841;
  wire tmp35842;
  wire tmp35843;
  wire tmp35844;
  wire tmp35845;
  wire tmp35846;
  wire tmp35847;
  wire tmp35848;
  wire tmp35849;
  wire tmp35850;
  wire tmp35851;
  wire tmp35852;
  wire tmp35853;
  wire tmp35854;
  wire tmp35855;
  wire tmp35856;
  wire tmp35857;
  wire tmp35858;
  wire tmp35859;
  wire tmp35860;
  wire tmp35861;
  wire tmp35862;
  wire tmp35863;
  wire tmp35864;
  wire tmp35865;
  wire tmp35866;
  wire tmp35867;
  wire tmp35868;
  wire tmp35869;
  wire tmp35870;
  wire tmp35871;
  wire tmp35872;
  wire tmp35873;
  wire tmp35874;
  wire tmp35875;
  wire tmp35876;
  wire tmp35877;
  wire tmp35878;
  wire tmp35879;
  wire tmp35880;
  wire tmp35881;
  wire tmp35882;
  wire tmp35883;
  wire tmp35884;
  wire tmp35885;
  wire tmp35886;
  wire tmp35887;
  wire tmp35888;
  wire tmp35889;
  wire tmp35890;
  wire tmp35891;
  wire tmp35892;
  wire tmp35893;
  wire tmp35894;
  wire tmp35895;
  wire tmp35896;
  wire tmp35897;
  wire tmp35898;
  wire tmp35899;
  wire tmp35900;
  wire tmp35901;
  wire tmp35902;
  wire tmp35903;
  wire tmp35904;
  wire tmp35905;
  wire tmp35906;
  wire tmp35907;
  wire tmp35908;
  wire tmp35909;
  wire tmp35910;
  wire tmp35911;
  wire tmp35912;
  wire tmp35913;
  wire tmp35914;
  wire tmp35915;
  wire tmp35916;
  wire tmp35917;
  wire tmp35918;
  wire tmp35919;
  wire tmp35920;
  wire tmp35921;
  wire tmp35922;
  wire tmp35923;
  wire tmp35924;
  wire tmp35925;
  wire tmp35926;
  wire tmp35927;
  wire tmp35928;
  wire tmp35929;
  wire tmp35930;
  wire tmp35931;
  wire tmp35932;
  wire tmp35933;
  wire tmp35934;
  wire tmp35935;
  wire tmp35936;
  wire tmp35937;
  wire tmp35938;
  wire tmp35939;
  wire tmp35940;
  wire tmp35941;
  wire tmp35942;
  wire tmp35943;
  wire tmp35944;
  wire tmp35945;
  wire tmp35946;
  wire tmp35947;
  wire tmp35948;
  wire tmp35949;
  wire tmp35950;
  wire tmp35951;
  wire tmp35952;
  wire tmp35953;
  wire tmp35954;
  wire tmp35955;
  wire tmp35956;
  wire tmp35957;
  wire tmp35958;
  wire tmp35959;
  wire tmp35960;
  wire tmp35961;
  wire tmp35962;
  wire tmp35963;
  wire tmp35964;
  wire tmp35965;
  wire tmp35966;
  wire tmp35967;
  wire tmp35968;
  wire tmp35969;
  wire tmp35970;
  wire tmp35971;
  wire tmp35972;
  wire tmp35973;
  wire tmp35974;
  wire tmp35975;
  wire tmp35976;
  wire tmp35977;
  wire tmp35978;
  wire tmp35979;
  wire tmp35980;
  wire tmp35981;
  wire tmp35982;
  wire tmp35983;
  wire tmp35984;
  wire tmp35985;
  wire tmp35986;
  wire tmp35987;
  wire tmp35988;
  wire tmp35989;
  wire tmp35990;
  wire tmp35991;
  wire tmp35992;
  wire tmp35993;
  wire tmp35994;
  wire tmp35995;
  wire tmp35996;
  wire tmp35997;
  wire tmp35998;
  wire tmp35999;
  wire tmp36000;
  wire tmp36001;
  wire tmp36002;
  wire tmp36003;
  wire tmp36004;
  wire tmp36005;
  wire tmp36006;
  wire tmp36007;
  wire tmp36008;
  wire tmp36009;
  wire tmp36010;
  wire tmp36011;
  wire tmp36012;
  wire tmp36013;
  wire tmp36014;
  wire tmp36015;
  wire tmp36016;
  wire tmp36017;
  wire tmp36018;
  wire tmp36019;
  wire tmp36020;
  wire tmp36021;
  wire tmp36022;
  wire tmp36023;
  wire tmp36024;
  wire tmp36025;
  wire tmp36026;
  wire tmp36027;
  wire tmp36028;
  wire tmp36029;
  wire tmp36030;
  wire tmp36031;
  wire tmp36032;
  wire tmp36033;
  wire tmp36034;
  wire tmp36035;
  wire tmp36036;
  wire tmp36037;
  wire tmp36038;
  wire tmp36039;
  wire tmp36040;
  wire tmp36041;
  wire tmp36042;
  wire tmp36043;
  wire tmp36044;
  wire tmp36045;
  wire tmp36046;
  wire tmp36047;
  wire tmp36048;
  wire tmp36049;
  wire tmp36050;
  wire tmp36051;
  wire tmp36052;
  wire tmp36053;
  wire tmp36054;
  wire tmp36055;
  wire tmp36056;
  wire tmp36057;
  wire tmp36058;
  wire tmp36059;
  wire tmp36060;
  wire tmp36061;
  wire tmp36062;
  wire tmp36063;
  wire tmp36064;
  wire tmp36065;
  wire tmp36066;
  wire tmp36067;
  wire tmp36068;
  wire tmp36069;
  wire tmp36070;
  wire tmp36071;
  wire tmp36072;
  wire tmp36073;
  wire tmp36074;
  wire tmp36075;
  wire tmp36076;
  wire tmp36077;
  wire tmp36078;
  wire tmp36079;
  wire tmp36080;
  wire tmp36081;
  wire tmp36082;
  wire tmp36083;
  wire tmp36084;
  wire tmp36085;
  wire tmp36086;
  wire tmp36087;
  wire tmp36088;
  wire tmp36089;
  wire tmp36090;
  wire tmp36091;
  wire tmp36092;
  wire tmp36093;
  wire tmp36094;
  wire tmp36095;
  wire tmp36096;
  wire tmp36097;
  wire tmp36098;
  wire tmp36099;
  wire tmp36100;
  wire tmp36101;
  wire tmp36102;
  wire tmp36103;
  wire tmp36104;
  wire tmp36105;
  wire tmp36106;
  wire tmp36107;
  wire tmp36108;
  wire tmp36109;
  wire tmp36110;
  wire tmp36111;
  wire tmp36112;
  wire tmp36113;
  wire tmp36114;
  wire tmp36115;
  wire tmp36116;
  wire tmp36117;
  wire tmp36118;
  wire tmp36119;
  wire tmp36120;
  wire tmp36121;
  wire tmp36122;
  wire tmp36123;
  wire tmp36124;
  wire tmp36125;
  wire tmp36126;
  wire tmp36127;
  wire tmp36128;
  wire tmp36129;
  wire tmp36130;
  wire tmp36131;
  wire tmp36132;
  wire tmp36133;
  wire tmp36134;
  wire tmp36135;
  wire tmp36136;
  wire tmp36137;
  wire tmp36138;
  wire tmp36139;
  wire tmp36140;
  wire tmp36141;
  wire tmp36142;
  wire tmp36143;
  wire tmp36144;
  wire tmp36145;
  wire tmp36146;
  wire tmp36147;
  wire tmp36148;
  wire tmp36149;
  wire tmp36150;
  wire tmp36151;
  wire tmp36152;
  wire tmp36153;
  wire tmp36154;
  wire tmp36155;
  wire tmp36156;
  wire tmp36157;
  wire tmp36158;
  wire tmp36159;
  wire tmp36160;
  wire tmp36161;
  wire tmp36162;
  wire tmp36163;
  wire tmp36164;
  wire tmp36165;
  wire tmp36166;
  wire tmp36167;
  wire tmp36168;
  wire tmp36169;
  wire tmp36170;
  wire tmp36171;
  wire tmp36172;
  wire tmp36173;
  wire tmp36174;
  wire tmp36175;
  wire tmp36176;
  wire tmp36177;
  wire tmp36178;
  wire tmp36179;
  wire tmp36180;
  wire tmp36181;
  wire tmp36182;
  wire tmp36183;
  wire tmp36184;
  wire tmp36185;
  wire tmp36186;
  wire tmp36187;
  wire tmp36188;
  wire tmp36189;
  wire tmp36190;
  wire tmp36191;
  wire tmp36192;
  wire tmp36193;
  wire tmp36194;
  wire tmp36195;
  wire tmp36196;
  wire tmp36197;
  wire tmp36198;
  wire tmp36199;
  wire tmp36200;
  wire tmp36201;
  wire tmp36202;
  wire tmp36203;
  wire tmp36204;
  wire tmp36205;
  wire tmp36206;
  wire tmp36207;
  wire tmp36208;
  wire tmp36209;
  wire tmp36210;
  wire tmp36211;
  wire tmp36212;
  wire tmp36213;
  wire tmp36214;
  wire tmp36215;
  wire tmp36216;
  wire tmp36217;
  wire tmp36218;
  wire tmp36219;
  wire tmp36220;
  wire tmp36221;
  wire tmp36222;
  wire tmp36223;
  wire tmp36224;
  wire tmp36225;
  wire tmp36226;
  wire tmp36227;
  wire tmp36228;
  wire tmp36229;
  wire tmp36230;
  wire tmp36231;
  wire tmp36232;
  wire tmp36233;
  wire tmp36234;
  wire tmp36235;
  wire tmp36236;
  wire tmp36237;
  wire tmp36238;
  wire tmp36239;
  wire tmp36240;
  wire tmp36241;
  wire tmp36242;
  wire tmp36243;
  wire tmp36244;
  wire tmp36245;
  wire tmp36246;
  wire tmp36247;
  wire tmp36248;
  wire tmp36249;
  wire tmp36250;
  wire tmp36251;
  wire tmp36252;
  wire tmp36253;
  wire tmp36254;
  wire tmp36255;
  wire tmp36256;
  wire tmp36257;
  wire tmp36258;
  wire tmp36259;
  wire tmp36260;
  wire tmp36261;
  wire tmp36262;
  wire tmp36263;
  wire tmp36264;
  wire tmp36265;
  wire tmp36266;
  wire tmp36267;
  wire tmp36268;
  wire tmp36269;
  wire tmp36270;
  wire tmp36271;
  wire tmp36272;
  wire tmp36273;
  wire tmp36274;
  wire tmp36275;
  wire tmp36276;
  wire tmp36277;
  wire tmp36278;
  wire tmp36279;
  wire tmp36280;
  wire tmp36281;
  wire tmp36282;
  wire tmp36283;
  wire tmp36284;
  wire tmp36285;
  wire tmp36286;
  wire tmp36287;
  wire tmp36288;
  wire tmp36289;
  wire tmp36290;
  wire tmp36291;
  wire tmp36292;
  wire tmp36293;
  wire tmp36294;
  wire tmp36295;
  wire tmp36296;
  wire tmp36297;
  wire tmp36298;
  wire tmp36299;
  wire tmp36300;
  wire tmp36301;
  wire tmp36302;
  wire tmp36303;
  wire tmp36304;
  wire tmp36305;
  wire tmp36306;
  wire tmp36307;
  wire tmp36308;
  wire tmp36309;
  wire tmp36310;
  wire tmp36311;
  wire tmp36312;
  wire tmp36313;
  wire tmp36314;
  wire tmp36315;
  wire tmp36316;
  wire tmp36317;
  wire tmp36318;
  wire tmp36319;
  wire tmp36320;
  wire tmp36321;
  wire tmp36322;
  wire tmp36323;
  wire tmp36324;
  wire tmp36325;
  wire tmp36326;
  wire tmp36327;
  wire tmp36328;
  wire tmp36329;
  wire tmp36330;
  wire tmp36331;
  wire tmp36332;
  wire tmp36333;
  wire tmp36334;
  wire tmp36335;
  wire tmp36336;
  wire tmp36337;
  wire tmp36338;
  wire tmp36339;
  wire tmp36340;
  wire tmp36341;
  wire tmp36342;
  wire tmp36343;
  wire tmp36344;
  wire tmp36345;
  wire tmp36346;
  wire tmp36347;
  wire tmp36348;
  wire tmp36349;
  wire tmp36350;
  wire tmp36351;
  wire tmp36352;
  wire tmp36353;
  wire tmp36354;
  wire tmp36355;
  wire tmp36356;
  wire tmp36357;
  wire tmp36358;
  wire tmp36359;
  wire tmp36360;
  wire tmp36361;
  wire tmp36362;
  wire tmp36363;
  wire tmp36364;
  wire tmp36365;
  wire tmp36366;
  wire tmp36367;
  wire tmp36368;
  wire tmp36369;
  wire tmp36370;
  wire tmp36371;
  wire tmp36372;
  wire tmp36373;
  wire tmp36374;
  wire tmp36375;
  wire tmp36376;
  wire tmp36377;
  wire tmp36378;
  wire tmp36379;
  wire tmp36380;
  wire tmp36381;
  wire tmp36382;
  wire tmp36383;
  wire tmp36384;
  wire tmp36385;
  wire tmp36386;
  wire tmp36387;
  wire tmp36388;
  wire tmp36389;
  wire tmp36390;
  wire tmp36391;
  wire tmp36392;
  wire tmp36393;
  wire tmp36394;
  wire tmp36395;
  wire tmp36396;
  wire tmp36397;
  wire tmp36398;
  wire tmp36399;
  wire tmp36400;
  wire tmp36401;
  wire tmp36402;
  wire tmp36403;
  wire tmp36404;
  wire tmp36405;
  wire tmp36406;
  wire tmp36407;
  wire tmp36408;
  wire tmp36409;
  wire tmp36410;
  wire tmp36411;
  wire tmp36412;
  wire tmp36413;
  wire tmp36414;
  wire tmp36415;
  wire tmp36416;
  wire tmp36417;
  wire tmp36418;
  wire tmp36419;
  wire tmp36420;
  wire tmp36421;
  wire tmp36422;
  wire tmp36423;
  wire tmp36424;
  wire tmp36425;
  wire tmp36426;
  wire tmp36427;
  wire tmp36428;
  wire tmp36429;
  wire tmp36430;
  wire tmp36431;
  wire tmp36432;
  wire tmp36433;
  wire tmp36434;
  wire tmp36435;
  wire tmp36436;
  wire tmp36437;
  wire tmp36438;
  wire tmp36439;
  wire tmp36440;
  wire tmp36441;
  wire tmp36442;
  wire tmp36443;
  wire tmp36444;
  wire tmp36445;
  wire tmp36446;
  wire tmp36447;
  wire tmp36448;
  wire tmp36449;
  wire tmp36450;
  wire tmp36451;
  wire tmp36452;
  wire tmp36453;
  wire tmp36454;
  wire tmp36455;
  wire tmp36456;
  wire tmp36457;
  wire tmp36458;
  wire tmp36459;
  wire tmp36460;
  wire tmp36461;
  wire tmp36462;
  wire tmp36463;
  wire tmp36464;
  wire tmp36465;
  wire tmp36466;
  wire tmp36467;
  wire tmp36468;
  wire tmp36469;
  wire tmp36470;
  wire tmp36471;
  wire tmp36472;
  wire tmp36473;
  wire tmp36474;
  wire tmp36475;
  wire tmp36476;
  wire tmp36477;
  wire tmp36478;
  wire tmp36479;
  wire tmp36480;
  wire tmp36481;
  wire tmp36482;
  wire tmp36483;
  wire tmp36484;
  wire tmp36485;
  wire tmp36486;
  wire tmp36487;
  wire tmp36488;
  wire tmp36489;
  wire tmp36490;
  wire tmp36491;
  wire tmp36492;
  wire tmp36493;
  wire tmp36494;
  wire tmp36495;
  wire tmp36496;
  wire tmp36497;
  wire tmp36498;
  wire tmp36499;
  wire tmp36500;
  wire tmp36501;
  wire tmp36502;
  wire tmp36503;
  wire tmp36504;
  wire tmp36505;
  wire tmp36506;
  wire tmp36507;
  wire tmp36508;
  wire tmp36509;
  wire tmp36510;
  wire tmp36511;
  wire tmp36512;
  wire tmp36513;
  wire tmp36514;
  wire tmp36515;
  wire tmp36516;
  wire tmp36517;
  wire tmp36518;
  wire tmp36519;
  wire tmp36520;
  wire tmp36521;
  wire tmp36522;
  wire tmp36523;
  wire tmp36524;
  wire tmp36525;
  wire tmp36526;
  wire tmp36527;
  wire tmp36528;
  wire tmp36529;
  wire tmp36530;
  wire tmp36531;
  wire tmp36532;
  wire tmp36533;
  wire tmp36534;
  wire tmp36535;
  wire tmp36536;
  wire tmp36537;
  wire tmp36538;
  wire tmp36539;
  wire tmp36540;
  wire tmp36541;
  wire tmp36542;
  wire tmp36543;
  wire tmp36544;
  wire tmp36545;
  wire tmp36546;
  wire tmp36547;
  wire tmp36548;
  wire tmp36549;
  wire tmp36550;
  wire tmp36551;
  wire tmp36552;
  wire tmp36553;
  wire tmp36554;
  wire tmp36555;
  wire tmp36556;
  wire tmp36557;
  wire tmp36558;
  wire tmp36559;
  wire tmp36560;
  wire tmp36561;
  wire tmp36562;
  wire tmp36563;
  wire tmp36564;
  wire tmp36565;
  wire tmp36566;
  wire tmp36567;
  wire tmp36568;
  wire tmp36569;
  wire tmp36570;
  wire tmp36571;
  wire tmp36572;
  wire tmp36573;
  wire tmp36574;
  wire tmp36575;
  wire tmp36576;
  wire tmp36577;
  wire tmp36578;
  wire tmp36579;
  wire tmp36580;
  wire tmp36581;
  wire tmp36582;
  wire tmp36583;
  wire tmp36584;
  wire tmp36585;
  wire tmp36586;
  wire tmp36587;
  wire tmp36588;
  wire tmp36589;
  wire tmp36590;
  wire tmp36591;
  wire tmp36592;
  wire tmp36593;
  wire tmp36594;
  wire tmp36595;
  wire tmp36596;
  wire tmp36597;
  wire tmp36598;
  wire tmp36599;
  wire tmp36600;
  wire tmp36601;
  wire tmp36602;
  wire tmp36603;
  wire tmp36604;
  wire tmp36605;
  wire tmp36606;
  wire tmp36607;
  wire tmp36608;
  wire tmp36609;
  wire tmp36610;
  wire tmp36611;
  wire tmp36612;
  wire tmp36613;
  wire tmp36614;
  wire tmp36615;
  wire tmp36616;
  wire tmp36617;
  wire tmp36618;
  wire tmp36619;
  wire tmp36620;
  wire tmp36621;
  wire tmp36622;
  wire tmp36623;
  wire tmp36624;
  wire tmp36625;
  wire tmp36626;
  wire tmp36627;
  wire tmp36628;
  wire tmp36629;
  wire tmp36630;
  wire tmp36631;
  wire tmp36632;
  wire tmp36633;
  wire tmp36634;
  wire tmp36635;
  wire tmp36636;
  wire tmp36637;
  wire tmp36638;
  wire tmp36639;
  wire tmp36640;
  wire tmp36641;
  wire tmp36642;
  wire tmp36643;
  wire tmp36644;
  wire tmp36645;
  wire tmp36646;
  wire tmp36647;
  wire tmp36648;
  wire tmp36649;
  wire tmp36650;
  wire tmp36651;
  wire tmp36652;
  wire tmp36653;
  wire tmp36654;
  wire tmp36655;
  wire tmp36656;
  wire tmp36657;
  wire tmp36658;
  wire tmp36659;
  wire tmp36660;
  wire tmp36661;
  wire tmp36662;
  wire tmp36663;
  wire tmp36664;
  wire tmp36665;
  wire tmp36666;
  wire tmp36667;
  wire tmp36668;
  wire tmp36669;
  wire tmp36670;
  wire tmp36671;
  wire tmp36672;
  wire tmp36673;
  wire tmp36674;
  wire tmp36675;
  wire tmp36676;
  wire tmp36677;
  wire tmp36678;
  wire tmp36679;
  wire tmp36680;
  wire tmp36681;
  wire tmp36682;
  wire tmp36683;
  wire tmp36684;
  wire tmp36685;
  wire tmp36686;
  wire tmp36687;
  wire tmp36688;
  wire tmp36689;
  wire tmp36690;
  wire tmp36691;
  wire tmp36692;
  wire tmp36693;
  wire tmp36694;
  wire tmp36695;
  wire tmp36696;
  wire tmp36697;
  wire tmp36698;
  wire tmp36699;
  wire tmp36700;
  wire tmp36701;
  wire tmp36702;
  wire tmp36703;
  wire tmp36704;
  wire tmp36705;
  wire tmp36706;
  wire tmp36707;
  wire tmp36708;
  wire tmp36709;
  wire tmp36710;
  wire tmp36711;
  wire tmp36712;
  wire tmp36713;
  wire tmp36714;
  wire tmp36715;
  wire tmp36716;
  wire tmp36717;
  wire tmp36718;
  wire tmp36719;
  wire tmp36720;
  wire tmp36721;
  wire tmp36722;
  wire tmp36723;
  wire tmp36724;
  wire tmp36725;
  wire tmp36726;
  wire tmp36727;
  wire tmp36728;
  wire tmp36729;
  wire tmp36730;
  wire tmp36731;
  wire tmp36732;
  wire tmp36733;
  wire tmp36734;
  wire tmp36735;
  wire tmp36736;
  wire tmp36737;
  wire tmp36738;
  wire tmp36739;
  wire tmp36740;
  wire tmp36741;
  wire tmp36742;
  wire tmp36743;
  wire tmp36744;
  wire tmp36745;
  wire tmp36746;
  wire tmp36747;
  wire tmp36748;
  wire tmp36749;
  wire tmp36750;
  wire tmp36751;
  wire tmp36752;
  wire tmp36753;
  wire tmp36754;
  wire tmp36755;
  wire tmp36756;
  wire tmp36757;
  wire tmp36758;
  wire tmp36759;
  wire tmp36760;
  wire tmp36761;
  wire tmp36762;
  wire tmp36763;
  wire tmp36764;
  wire tmp36765;
  wire tmp36766;
  wire tmp36767;
  wire tmp36768;
  wire tmp36769;
  wire tmp36770;
  wire tmp36771;
  wire tmp36772;
  wire tmp36773;
  wire tmp36774;
  wire tmp36775;
  wire tmp36776;
  wire tmp36777;
  wire tmp36778;
  wire tmp36779;
  wire tmp36780;
  wire tmp36781;
  wire tmp36782;
  wire tmp36783;
  wire tmp36784;
  wire tmp36785;
  wire tmp36786;
  wire tmp36787;
  wire tmp36788;
  wire tmp36789;
  wire tmp36790;
  wire tmp36791;
  wire tmp36792;
  wire tmp36793;
  wire tmp36794;
  wire tmp36795;
  wire tmp36796;
  wire tmp36797;
  wire tmp36798;
  wire tmp36799;
  wire tmp36800;
  wire tmp36801;
  wire tmp36802;
  wire tmp36803;
  wire tmp36804;
  wire tmp36805;
  wire tmp36806;
  wire tmp36807;
  wire tmp36808;
  wire tmp36809;
  wire tmp36810;
  wire tmp36811;
  wire tmp36812;
  wire tmp36813;
  wire tmp36814;
  wire tmp36815;
  wire tmp36816;
  wire tmp36817;
  wire tmp36818;
  wire tmp36819;
  wire tmp36820;
  wire tmp36821;
  wire tmp36822;
  wire tmp36823;
  wire tmp36824;
  wire tmp36825;
  wire tmp36826;
  wire tmp36827;
  wire tmp36828;
  wire tmp36829;
  wire tmp36830;
  wire tmp36831;
  wire tmp36832;
  wire tmp36833;
  wire tmp36834;
  wire tmp36835;
  wire tmp36836;
  wire tmp36837;
  wire tmp36838;
  wire tmp36839;
  wire tmp36840;
  wire tmp36841;
  wire tmp36842;
  wire tmp36843;
  wire tmp36844;
  wire tmp36845;
  wire tmp36846;
  wire tmp36847;
  wire tmp36848;
  wire tmp36849;
  wire tmp36850;
  wire tmp36851;
  wire tmp36852;
  wire tmp36853;
  wire tmp36854;
  wire tmp36855;
  wire tmp36856;
  wire tmp36857;
  wire tmp36858;
  wire tmp36859;
  wire tmp36860;
  wire tmp36861;
  wire tmp36862;
  wire tmp36863;
  wire tmp36864;
  wire tmp36865;
  wire tmp36866;
  wire tmp36867;
  wire tmp36868;
  wire tmp36869;
  wire tmp36870;
  wire tmp36871;
  wire tmp36872;
  wire tmp36873;
  wire tmp36874;
  wire tmp36875;
  wire tmp36876;
  wire tmp36877;
  wire tmp36878;
  wire tmp36879;
  wire tmp36880;
  wire tmp36881;
  wire tmp36882;
  wire tmp36883;
  wire tmp36884;
  wire tmp36885;
  wire tmp36886;
  wire tmp36887;
  wire tmp36888;
  wire tmp36889;
  wire tmp36890;
  wire tmp36891;
  wire tmp36892;
  wire tmp36893;
  wire tmp36894;
  wire tmp36895;
  wire tmp36896;
  wire tmp36897;
  wire tmp36898;
  wire tmp36899;
  wire tmp36900;
  wire tmp36901;
  wire tmp36902;
  wire tmp36903;
  wire tmp36904;
  wire tmp36905;
  wire tmp36906;
  wire tmp36907;
  wire tmp36908;
  wire tmp36909;
  wire tmp36910;
  wire tmp36911;
  wire tmp36912;
  wire tmp36913;
  wire tmp36914;
  wire tmp36915;
  wire tmp36916;
  wire tmp36917;
  wire tmp36918;
  wire tmp36919;
  wire tmp36920;
  wire tmp36921;
  wire tmp36922;
  wire tmp36923;
  wire tmp36924;
  wire tmp36925;
  wire tmp36926;
  wire tmp36927;
  wire tmp36928;
  wire tmp36929;
  wire tmp36930;
  wire tmp36931;
  wire tmp36932;
  wire tmp36933;
  wire tmp36934;
  wire tmp36935;
  wire tmp36936;
  wire tmp36937;
  wire tmp36938;
  wire tmp36939;
  wire tmp36940;
  wire tmp36941;
  wire tmp36942;
  wire tmp36943;
  wire tmp36944;
  wire tmp36945;
  wire tmp36946;
  wire tmp36947;
  wire tmp36948;
  wire tmp36949;
  wire tmp36950;
  wire tmp36951;
  wire tmp36952;
  wire tmp36953;
  wire tmp36954;
  wire tmp36955;
  wire tmp36956;
  wire tmp36957;
  wire tmp36958;
  wire tmp36959;
  wire tmp36960;
  wire tmp36961;
  wire tmp36962;
  wire tmp36963;
  wire tmp36964;
  wire tmp36965;
  wire tmp36966;
  wire tmp36967;
  wire tmp36968;
  wire tmp36969;
  wire tmp36970;
  wire tmp36971;
  wire tmp36972;
  wire tmp36973;
  wire tmp36974;
  wire tmp36975;
  wire tmp36976;
  wire tmp36977;
  wire tmp36978;
  wire tmp36979;
  wire tmp36980;
  wire tmp36981;
  wire tmp36982;
  wire tmp36983;
  wire tmp36984;
  wire tmp36985;
  wire tmp36986;
  wire tmp36987;
  wire tmp36988;
  wire tmp36989;
  wire tmp36990;
  wire tmp36991;
  wire tmp36992;
  wire tmp36993;
  wire tmp36994;
  wire tmp36995;
  wire tmp36996;
  wire tmp36997;
  wire tmp36998;
  wire tmp36999;
  wire tmp37000;
  wire tmp37001;
  wire tmp37002;
  wire tmp37003;
  wire tmp37004;
  wire tmp37005;
  wire tmp37006;
  wire tmp37007;
  wire tmp37008;
  wire tmp37009;
  wire tmp37010;
  wire tmp37011;
  wire tmp37012;
  wire tmp37013;
  wire tmp37014;
  wire tmp37015;
  wire tmp37016;
  wire tmp37017;
  wire tmp37018;
  wire tmp37019;
  wire tmp37020;
  wire tmp37021;
  wire tmp37022;
  wire tmp37023;
  wire tmp37024;
  wire tmp37025;
  wire tmp37026;
  wire tmp37027;
  wire tmp37028;
  wire tmp37029;
  wire tmp37030;
  wire tmp37031;
  wire tmp37032;
  wire tmp37033;
  wire tmp37034;
  wire tmp37035;
  wire tmp37036;
  wire tmp37037;
  wire tmp37038;
  wire tmp37039;
  wire tmp37040;
  wire tmp37041;
  wire tmp37042;
  wire tmp37043;
  wire tmp37044;
  wire tmp37045;
  wire tmp37046;
  wire tmp37047;
  wire tmp37048;
  wire tmp37049;
  wire tmp37050;
  wire tmp37051;
  wire tmp37052;
  wire tmp37053;
  wire tmp37054;
  wire tmp37055;
  wire tmp37056;
  wire tmp37057;
  wire tmp37058;
  wire tmp37059;
  wire tmp37060;
  wire tmp37061;
  wire tmp37062;
  wire tmp37063;
  wire tmp37064;
  wire tmp37065;
  wire tmp37066;
  wire tmp37067;
  wire tmp37068;
  wire tmp37069;
  wire tmp37070;
  wire tmp37071;
  wire tmp37072;
  wire tmp37073;
  wire tmp37074;
  wire tmp37075;
  wire tmp37076;
  wire tmp37077;
  wire tmp37078;
  wire tmp37079;
  wire tmp37080;
  wire tmp37081;
  wire tmp37082;
  wire tmp37083;
  wire tmp37084;
  wire tmp37085;
  wire tmp37086;
  wire tmp37087;
  wire tmp37088;
  wire tmp37089;
  wire tmp37090;
  wire tmp37091;
  wire tmp37092;
  wire tmp37093;
  wire tmp37094;
  wire tmp37095;
  wire tmp37096;
  wire tmp37097;
  wire tmp37098;
  wire tmp37099;
  wire tmp37100;
  wire tmp37101;
  wire tmp37102;
  wire tmp37103;
  wire tmp37104;
  wire tmp37105;
  wire tmp37106;
  wire tmp37107;
  wire tmp37108;
  wire tmp37109;
  wire tmp37110;
  wire tmp37111;
  wire tmp37112;
  wire tmp37113;
  wire tmp37114;
  wire tmp37115;
  wire tmp37116;
  wire tmp37117;
  wire tmp37118;
  wire tmp37119;
  wire tmp37120;
  wire tmp37121;
  wire tmp37122;
  wire tmp37123;
  wire tmp37124;
  wire tmp37125;
  wire tmp37126;
  wire tmp37127;
  wire tmp37128;
  wire tmp37129;
  wire tmp37130;
  wire tmp37131;
  wire tmp37132;
  wire tmp37133;
  wire tmp37134;
  wire tmp37135;
  wire tmp37136;
  wire tmp37137;
  wire tmp37138;
  wire tmp37139;
  wire tmp37140;
  wire tmp37141;
  wire tmp37142;
  wire tmp37143;
  wire tmp37144;
  wire tmp37145;
  wire tmp37146;
  wire tmp37147;
  wire tmp37148;
  wire tmp37149;
  wire tmp37150;
  wire tmp37151;
  wire tmp37152;
  wire tmp37153;
  wire tmp37154;
  wire tmp37155;
  wire tmp37156;
  wire tmp37157;
  wire tmp37158;
  wire tmp37159;
  wire tmp37160;
  wire tmp37161;
  wire tmp37162;
  wire tmp37163;
  wire tmp37164;
  wire tmp37165;
  wire tmp37166;
  wire tmp37167;
  wire tmp37168;
  wire tmp37169;
  wire tmp37170;
  wire tmp37171;
  wire tmp37172;
  wire tmp37173;
  wire tmp37174;
  wire tmp37175;
  wire tmp37176;
  wire tmp37177;
  wire tmp37178;
  wire tmp37179;
  wire tmp37180;
  wire tmp37181;
  wire tmp37182;
  wire tmp37183;
  wire tmp37184;
  wire tmp37185;
  wire tmp37186;
  wire tmp37187;
  wire tmp37188;
  wire tmp37189;
  wire tmp37190;
  wire tmp37191;
  wire tmp37192;
  wire tmp37193;
  wire tmp37194;
  wire tmp37195;
  wire tmp37196;
  wire tmp37197;
  wire tmp37198;
  wire tmp37199;
  wire tmp37200;
  wire tmp37201;
  wire tmp37202;
  wire tmp37203;
  wire tmp37204;
  wire tmp37205;
  wire tmp37206;
  wire tmp37207;
  wire tmp37208;
  wire tmp37209;
  wire tmp37210;
  wire tmp37211;
  wire tmp37212;
  wire tmp37213;
  wire tmp37214;
  wire tmp37215;
  wire tmp37216;
  wire tmp37217;
  wire tmp37218;
  wire tmp37219;
  wire tmp37220;
  wire tmp37221;
  wire tmp37222;
  wire tmp37223;
  wire tmp37224;
  wire tmp37225;
  wire tmp37226;
  wire tmp37227;
  wire tmp37228;
  wire tmp37229;
  wire tmp37230;
  wire tmp37231;
  wire tmp37232;
  wire tmp37233;
  wire tmp37234;
  wire tmp37235;
  wire tmp37236;
  wire tmp37237;
  wire tmp37238;
  wire tmp37239;
  wire tmp37240;
  wire tmp37241;
  wire tmp37242;
  wire tmp37243;
  wire tmp37244;
  wire tmp37245;
  wire tmp37246;
  wire tmp37247;
  wire tmp37248;
  wire tmp37249;
  wire tmp37250;
  wire tmp37251;
  wire tmp37252;
  wire tmp37253;
  wire tmp37254;
  wire tmp37255;
  wire tmp37256;
  wire tmp37257;
  wire tmp37258;
  wire tmp37259;
  wire tmp37260;
  wire tmp37261;
  wire tmp37262;
  wire tmp37263;
  wire tmp37264;
  wire tmp37265;
  wire tmp37266;
  wire tmp37267;
  wire tmp37268;
  wire tmp37269;
  wire tmp37270;
  wire tmp37271;
  wire tmp37272;
  wire tmp37273;
  wire tmp37274;
  wire tmp37275;
  wire tmp37276;
  wire tmp37277;
  wire tmp37278;
  wire tmp37279;
  wire tmp37280;
  wire tmp37281;
  wire tmp37282;
  wire tmp37283;
  wire tmp37284;
  wire tmp37285;
  wire tmp37286;
  wire tmp37287;
  wire tmp37288;
  wire tmp37289;
  wire tmp37290;
  wire tmp37291;
  wire tmp37292;
  wire tmp37293;
  wire tmp37294;
  wire tmp37295;
  wire tmp37296;
  wire tmp37297;
  wire tmp37298;
  wire tmp37299;
  wire tmp37300;
  wire tmp37301;
  wire tmp37302;
  wire tmp37303;
  wire tmp37304;
  wire tmp37305;
  wire tmp37306;
  wire tmp37307;
  wire tmp37308;
  wire tmp37309;
  wire tmp37310;
  wire tmp37311;
  wire tmp37312;
  wire tmp37313;
  wire tmp37314;
  wire tmp37315;
  wire tmp37316;
  wire tmp37317;
  wire tmp37318;
  wire tmp37319;
  wire tmp37320;
  wire tmp37321;
  wire tmp37322;
  wire tmp37323;
  wire tmp37324;
  wire tmp37325;
  wire tmp37326;
  wire tmp37327;
  wire tmp37328;
  wire tmp37329;
  wire tmp37330;
  wire tmp37331;
  wire tmp37332;
  wire tmp37333;
  wire tmp37334;
  wire tmp37335;
  wire tmp37336;
  wire tmp37337;
  wire tmp37338;
  wire tmp37339;
  wire tmp37340;
  wire tmp37341;
  wire tmp37342;
  wire tmp37343;
  wire tmp37344;
  wire tmp37345;
  wire tmp37346;
  wire tmp37347;
  wire tmp37348;
  wire tmp37349;
  wire tmp37350;
  wire tmp37351;
  wire tmp37352;
  wire tmp37353;
  wire tmp37354;
  wire tmp37355;
  wire tmp37356;
  wire tmp37357;
  wire tmp37358;
  wire tmp37359;
  wire tmp37360;
  wire tmp37361;
  wire tmp37362;
  wire tmp37363;
  wire tmp37364;
  wire tmp37365;
  wire tmp37366;
  wire tmp37367;
  wire tmp37368;
  wire tmp37369;
  wire tmp37370;
  wire tmp37371;
  wire tmp37372;
  wire tmp37373;
  wire tmp37374;
  wire tmp37375;
  wire tmp37376;
  wire tmp37377;
  wire tmp37378;
  wire tmp37379;
  wire tmp37380;
  wire tmp37381;
  wire tmp37382;
  wire tmp37383;
  wire tmp37384;
  wire tmp37385;
  wire tmp37386;
  wire tmp37387;
  wire tmp37388;
  wire tmp37389;
  wire tmp37390;
  wire tmp37391;
  wire tmp37392;
  wire tmp37393;
  wire tmp37394;
  wire tmp37395;
  wire tmp37396;
  wire tmp37397;
  wire tmp37398;
  wire tmp37399;
  wire tmp37400;
  wire tmp37401;
  wire tmp37402;
  wire tmp37403;
  wire tmp37404;
  wire tmp37405;
  wire tmp37406;
  wire tmp37407;
  wire tmp37408;
  wire tmp37409;
  wire tmp37410;
  wire tmp37411;
  wire tmp37412;
  wire tmp37413;
  wire tmp37414;
  wire tmp37415;
  wire tmp37416;
  wire tmp37417;
  wire tmp37418;
  wire tmp37419;
  wire tmp37420;
  wire tmp37421;
  wire tmp37422;
  wire tmp37423;
  wire tmp37424;
  wire tmp37425;
  wire tmp37426;
  wire tmp37427;
  wire tmp37428;
  wire tmp37429;
  wire tmp37430;
  wire tmp37431;
  wire tmp37432;
  wire tmp37433;
  wire tmp37434;
  wire tmp37435;
  wire tmp37436;
  wire tmp37437;
  wire tmp37438;
  wire tmp37439;
  wire tmp37440;
  wire tmp37441;
  wire tmp37442;
  wire tmp37443;
  wire tmp37444;
  wire tmp37445;
  wire tmp37446;
  wire tmp37447;
  wire tmp37448;
  wire tmp37449;
  wire tmp37450;
  wire tmp37451;
  wire tmp37452;
  wire tmp37453;
  wire tmp37454;
  wire tmp37455;
  wire tmp37456;
  wire tmp37457;
  wire tmp37458;
  wire tmp37459;
  wire tmp37460;
  wire tmp37461;
  wire tmp37462;
  wire tmp37463;
  wire tmp37464;
  wire tmp37465;
  wire tmp37466;
  wire tmp37467;
  wire tmp37468;
  wire tmp37469;
  wire tmp37470;
  wire tmp37471;
  wire tmp37472;
  wire tmp37473;
  wire tmp37474;
  wire tmp37475;
  wire tmp37476;
  wire tmp37477;
  wire tmp37478;
  wire tmp37479;
  wire tmp37480;
  wire tmp37481;
  wire tmp37482;
  wire tmp37483;
  wire tmp37484;
  wire tmp37485;
  wire tmp37486;
  wire tmp37487;
  wire tmp37488;
  wire tmp37489;
  wire tmp37490;
  wire tmp37491;
  wire tmp37492;
  wire tmp37493;
  wire tmp37494;
  wire tmp37495;
  wire tmp37496;
  wire tmp37497;
  wire tmp37498;
  wire tmp37499;
  wire tmp37500;
  wire tmp37501;
  wire tmp37502;
  wire tmp37503;
  wire tmp37504;
  wire tmp37505;
  wire tmp37506;
  wire tmp37507;
  wire tmp37508;
  wire tmp37509;
  wire tmp37510;
  wire tmp37511;
  wire tmp37512;
  wire tmp37513;
  wire tmp37514;
  wire tmp37515;
  wire tmp37516;
  wire tmp37517;
  wire tmp37518;
  wire tmp37519;
  wire tmp37520;
  wire tmp37521;
  wire tmp37522;
  wire tmp37523;
  wire tmp37524;
  wire tmp37525;
  wire tmp37526;
  wire tmp37527;
  wire tmp37528;
  wire tmp37529;
  wire tmp37530;
  wire tmp37531;
  wire tmp37532;
  wire tmp37533;
  wire tmp37534;
  wire tmp37535;
  wire tmp37536;
  wire tmp37537;
  wire tmp37538;
  wire tmp37539;
  wire tmp37540;
  wire tmp37541;
  wire tmp37542;
  wire tmp37543;
  wire tmp37544;
  wire tmp37545;
  wire tmp37546;
  wire tmp37547;
  wire tmp37548;
  wire tmp37549;
  wire tmp37550;
  wire tmp37551;
  wire tmp37552;
  wire tmp37553;
  wire tmp37554;
  wire tmp37555;
  wire tmp37556;
  wire tmp37557;
  wire tmp37558;
  wire tmp37559;
  wire tmp37560;
  wire tmp37561;
  wire tmp37562;
  wire tmp37563;
  wire tmp37564;
  wire tmp37565;
  wire tmp37566;
  wire tmp37567;
  wire tmp37568;
  wire tmp37569;
  wire tmp37570;
  wire tmp37571;
  wire tmp37572;
  wire tmp37573;
  wire tmp37574;
  wire tmp37575;
  wire tmp37576;
  wire tmp37577;
  wire tmp37578;
  wire tmp37579;
  wire tmp37580;
  wire tmp37581;
  wire tmp37582;
  wire tmp37583;
  wire tmp37584;
  wire tmp37585;
  wire tmp37586;
  wire tmp37587;
  wire tmp37588;
  wire tmp37589;
  wire tmp37590;
  wire tmp37591;
  wire tmp37592;
  wire tmp37593;
  wire tmp37594;
  wire tmp37595;
  wire tmp37596;
  wire tmp37597;
  wire tmp37598;
  wire tmp37599;
  wire tmp37600;
  wire tmp37601;
  wire tmp37602;
  wire tmp37603;
  wire tmp37604;
  wire tmp37605;
  wire tmp37606;
  wire tmp37607;
  wire tmp37608;
  wire tmp37609;
  wire tmp37610;
  wire tmp37611;
  wire tmp37612;
  wire tmp37613;
  wire tmp37614;
  wire tmp37615;
  wire tmp37616;
  wire tmp37617;
  wire tmp37618;
  wire tmp37619;
  wire tmp37620;
  wire tmp37621;
  wire tmp37622;
  wire tmp37623;
  wire tmp37624;
  wire tmp37625;
  wire tmp37626;
  wire tmp37627;
  wire tmp37628;
  wire tmp37629;
  wire tmp37630;
  wire tmp37631;
  wire tmp37632;
  wire tmp37633;
  wire tmp37634;
  wire tmp37635;
  wire tmp37636;
  wire tmp37637;
  wire tmp37638;
  wire tmp37639;
  wire tmp37640;
  wire tmp37641;
  wire tmp37642;
  wire tmp37643;
  wire tmp37644;
  wire tmp37645;
  wire tmp37646;
  wire tmp37647;
  wire tmp37648;
  wire tmp37649;
  wire tmp37650;
  wire tmp37651;
  wire tmp37652;
  wire tmp37653;
  wire tmp37654;
  wire tmp37655;
  wire tmp37656;
  wire tmp37657;
  wire tmp37658;
  wire tmp37659;
  wire tmp37660;
  wire tmp37661;
  wire tmp37662;
  wire tmp37663;
  wire tmp37664;
  wire tmp37665;
  wire tmp37666;
  wire tmp37667;
  wire tmp37668;
  wire tmp37669;
  wire tmp37670;
  wire tmp37671;
  wire tmp37672;
  wire tmp37673;
  wire tmp37674;
  wire tmp37675;
  wire tmp37676;
  wire tmp37677;
  wire tmp37678;
  wire tmp37679;
  wire tmp37680;
  wire tmp37681;
  wire tmp37682;
  wire tmp37683;
  wire tmp37684;
  wire tmp37685;
  wire tmp37686;
  wire tmp37687;
  wire tmp37688;
  wire tmp37689;
  wire tmp37690;
  wire tmp37691;
  wire tmp37692;
  wire tmp37693;
  wire tmp37694;
  wire tmp37695;
  wire tmp37696;
  wire tmp37697;
  wire tmp37698;
  wire tmp37699;
  wire tmp37700;
  wire tmp37701;
  wire tmp37702;
  wire tmp37703;
  wire tmp37704;
  wire tmp37705;
  wire tmp37706;
  wire tmp37707;
  wire tmp37708;
  wire tmp37709;
  wire tmp37710;
  wire tmp37711;
  wire tmp37712;
  wire tmp37713;
  wire tmp37714;
  wire tmp37715;
  wire tmp37716;
  wire tmp37717;
  wire tmp37718;
  wire tmp37719;
  wire tmp37720;
  wire tmp37721;
  wire tmp37722;
  wire tmp37723;
  wire tmp37724;
  wire tmp37725;
  wire tmp37726;
  wire tmp37727;
  wire tmp37728;
  wire tmp37729;
  wire tmp37730;
  wire tmp37731;
  wire tmp37732;
  wire tmp37733;
  wire tmp37734;
  wire tmp37735;
  wire tmp37736;
  wire tmp37737;
  wire tmp37738;
  wire tmp37739;
  wire tmp37740;
  wire tmp37741;
  wire tmp37742;
  wire tmp37743;
  wire tmp37744;
  wire tmp37745;
  wire tmp37746;
  wire tmp37747;
  wire tmp37748;
  wire tmp37749;
  wire tmp37750;
  wire tmp37751;
  wire tmp37752;
  wire tmp37753;
  wire tmp37754;
  wire tmp37755;
  wire tmp37756;
  wire tmp37757;
  wire tmp37758;
  wire tmp37759;
  wire tmp37760;
  wire tmp37761;
  wire tmp37762;
  wire tmp37763;
  wire tmp37764;
  wire tmp37765;
  wire tmp37766;
  wire tmp37767;
  wire tmp37768;
  wire tmp37769;
  wire tmp37770;
  wire tmp37771;
  wire tmp37772;
  wire tmp37773;
  wire tmp37774;
  wire tmp37775;
  wire tmp37776;
  wire tmp37777;
  wire tmp37778;
  wire tmp37779;
  wire tmp37780;
  wire tmp37781;
  wire tmp37782;
  wire tmp37783;
  wire tmp37784;
  wire tmp37785;
  wire tmp37786;
  wire tmp37787;
  wire tmp37788;
  wire tmp37789;
  wire tmp37790;
  wire tmp37791;
  wire tmp37792;
  wire tmp37793;
  wire tmp37794;
  wire tmp37795;
  wire tmp37796;
  wire tmp37797;
  wire tmp37798;
  wire tmp37799;
  wire tmp37800;
  wire tmp37801;
  wire tmp37802;
  wire tmp37803;
  wire tmp37804;
  wire tmp37805;
  wire tmp37806;
  wire tmp37807;
  wire tmp37808;
  wire tmp37809;
  wire tmp37810;
  wire tmp37811;
  wire tmp37812;
  wire tmp37813;
  wire tmp37814;
  wire tmp37815;
  wire tmp37816;
  wire tmp37817;
  wire tmp37818;
  wire tmp37819;
  wire tmp37820;
  wire tmp37821;
  wire tmp37822;
  wire tmp37823;
  wire tmp37824;
  wire tmp37825;
  wire tmp37826;
  wire tmp37827;
  wire tmp37828;
  wire tmp37829;
  wire tmp37830;
  wire tmp37831;
  wire tmp37832;
  wire tmp37833;
  wire tmp37834;
  wire tmp37835;
  wire tmp37836;
  wire tmp37837;
  wire tmp37838;
  wire tmp37839;
  wire tmp37840;
  wire tmp37841;
  wire tmp37842;
  wire tmp37843;
  wire tmp37844;
  wire tmp37845;
  wire tmp37846;
  wire tmp37847;
  wire tmp37848;
  wire tmp37849;
  wire tmp37850;
  wire tmp37851;
  wire tmp37852;
  wire tmp37853;
  wire tmp37854;
  wire tmp37855;
  wire tmp37856;
  wire tmp37857;
  wire tmp37858;
  wire tmp37859;
  wire tmp37860;
  wire tmp37861;
  wire tmp37862;
  wire tmp37863;
  wire tmp37864;
  wire tmp37865;
  wire tmp37866;
  wire tmp37867;
  wire tmp37868;
  wire tmp37869;
  wire tmp37870;
  wire tmp37871;
  wire tmp37872;
  wire tmp37873;
  wire tmp37874;
  wire tmp37875;
  wire tmp37876;
  wire tmp37877;
  wire tmp37878;
  wire tmp37879;
  wire tmp37880;
  wire tmp37881;
  wire tmp37882;
  wire tmp37883;
  wire tmp37884;
  wire tmp37885;
  wire tmp37886;
  wire tmp37887;
  wire tmp37888;
  wire tmp37889;
  wire tmp37890;
  wire tmp37891;
  wire tmp37892;
  wire tmp37893;
  wire tmp37894;
  wire tmp37895;
  wire tmp37896;
  wire tmp37897;
  wire tmp37898;
  wire tmp37899;
  wire tmp37900;
  wire tmp37901;
  wire tmp37902;
  wire tmp37903;
  wire tmp37904;
  wire tmp37905;
  wire tmp37906;
  wire tmp37907;
  wire tmp37908;
  wire tmp37909;
  wire tmp37910;
  wire tmp37911;
  wire tmp37912;
  wire tmp37913;
  wire tmp37914;
  wire tmp37915;
  wire tmp37916;
  wire tmp37917;
  wire tmp37918;
  wire tmp37919;
  wire tmp37920;
  wire tmp37921;
  wire tmp37922;
  wire tmp37923;
  wire tmp37924;
  wire tmp37925;
  wire tmp37926;
  wire tmp37927;
  wire tmp37928;
  wire tmp37929;
  wire tmp37930;
  wire tmp37931;
  wire tmp37932;
  wire tmp37933;
  wire tmp37934;
  wire tmp37935;
  wire tmp37936;
  wire tmp37937;
  wire tmp37938;
  wire tmp37939;
  wire tmp37940;
  wire tmp37941;
  wire tmp37942;
  wire tmp37943;
  wire tmp37944;
  wire tmp37945;
  wire tmp37946;
  wire tmp37947;
  wire tmp37948;
  wire tmp37949;
  wire tmp37950;
  wire tmp37951;
  wire tmp37952;
  wire tmp37953;
  wire tmp37954;
  wire tmp37955;
  wire tmp37956;
  wire tmp37957;
  wire tmp37958;
  wire tmp37959;
  wire tmp37960;
  wire tmp37961;
  wire tmp37962;
  wire tmp37963;
  wire tmp37964;
  wire tmp37965;
  wire tmp37966;
  wire tmp37967;
  wire tmp37968;
  wire tmp37969;
  wire tmp37970;
  wire tmp37971;
  wire tmp37972;
  wire tmp37973;
  wire tmp37974;
  wire tmp37975;
  wire tmp37976;
  wire tmp37977;
  wire tmp37978;
  wire tmp37979;
  wire tmp37980;
  wire tmp37981;
  wire tmp37982;
  wire tmp37983;
  wire tmp37984;
  wire tmp37985;
  wire tmp37986;
  wire tmp37987;
  wire tmp37988;
  wire tmp37989;
  wire tmp37990;
  wire tmp37991;
  wire tmp37992;
  wire tmp37993;
  wire tmp37994;
  wire tmp37995;
  wire tmp37996;
  wire tmp37997;
  wire tmp37998;
  wire tmp37999;
  wire tmp38000;
  wire tmp38001;
  wire tmp38002;
  wire tmp38003;
  wire tmp38004;
  wire tmp38005;
  wire tmp38006;
  wire tmp38007;
  wire tmp38008;
  wire tmp38009;
  wire tmp38010;
  wire tmp38011;
  wire tmp38012;
  wire tmp38013;
  wire tmp38014;
  wire tmp38015;
  wire tmp38016;
  wire tmp38017;
  wire tmp38018;
  wire tmp38019;
  wire tmp38020;
  wire tmp38021;
  wire tmp38022;
  wire tmp38023;
  wire tmp38024;
  wire tmp38025;
  wire tmp38026;
  wire tmp38027;
  wire tmp38028;
  wire tmp38029;
  wire tmp38030;
  wire tmp38031;
  wire tmp38032;
  wire tmp38033;
  wire tmp38034;
  wire tmp38035;
  wire tmp38036;
  wire tmp38037;
  wire tmp38038;
  wire tmp38039;
  wire tmp38040;
  wire tmp38041;
  wire tmp38042;
  wire tmp38043;
  wire tmp38044;
  wire tmp38045;
  wire tmp38046;
  wire tmp38047;
  wire tmp38048;
  wire tmp38049;
  wire tmp38050;
  wire tmp38051;
  wire tmp38052;
  wire tmp38053;
  wire tmp38054;
  wire tmp38055;
  wire tmp38056;
  wire tmp38057;
  wire tmp38058;
  wire tmp38059;
  wire tmp38060;
  wire tmp38061;
  wire tmp38062;
  wire tmp38063;
  wire tmp38064;
  wire tmp38065;
  wire tmp38066;
  wire tmp38067;
  wire tmp38068;
  wire tmp38069;
  wire tmp38070;
  wire tmp38071;
  wire tmp38072;
  wire tmp38073;
  wire tmp38074;
  wire tmp38075;
  wire tmp38076;
  wire tmp38077;
  wire tmp38078;
  wire tmp38079;
  wire tmp38080;
  wire tmp38081;
  wire tmp38082;
  wire tmp38083;
  wire tmp38084;
  wire tmp38085;
  wire tmp38086;
  wire tmp38087;
  wire tmp38088;
  wire tmp38089;
  wire tmp38090;
  wire tmp38091;
  wire tmp38092;
  wire tmp38093;
  wire tmp38094;
  wire tmp38095;
  wire tmp38096;
  wire tmp38097;
  wire tmp38098;
  wire tmp38099;
  wire tmp38100;
  wire tmp38101;
  wire tmp38102;
  wire tmp38103;
  wire tmp38104;
  wire tmp38105;
  wire tmp38106;
  wire tmp38107;
  wire tmp38108;
  wire tmp38109;
  wire tmp38110;
  wire tmp38111;
  wire tmp38112;
  wire tmp38113;
  wire tmp38114;
  wire tmp38115;
  wire tmp38116;
  wire tmp38117;
  wire tmp38118;
  wire tmp38119;
  wire tmp38120;
  wire tmp38121;
  wire tmp38122;
  wire tmp38123;
  wire tmp38124;
  wire tmp38125;
  wire tmp38126;
  wire tmp38127;
  wire tmp38128;
  wire tmp38129;
  wire tmp38130;
  wire tmp38131;
  wire tmp38132;
  wire tmp38133;
  wire tmp38134;
  wire tmp38135;
  wire tmp38136;
  wire tmp38137;
  wire tmp38138;
  wire tmp38139;
  wire tmp38140;
  wire tmp38141;
  wire tmp38142;
  wire tmp38143;
  wire tmp38144;
  wire tmp38145;
  wire tmp38146;
  wire tmp38147;
  wire tmp38148;
  wire tmp38149;
  wire tmp38150;
  wire tmp38151;
  wire tmp38152;
  wire tmp38153;
  wire tmp38154;
  wire tmp38155;
  wire tmp38156;
  wire tmp38157;
  wire tmp38158;
  wire tmp38159;
  wire tmp38160;
  wire tmp38161;
  wire tmp38162;
  wire tmp38163;
  wire tmp38164;
  wire tmp38165;
  wire tmp38166;
  wire tmp38167;
  wire tmp38168;
  wire tmp38169;
  wire tmp38170;
  wire tmp38171;
  wire tmp38172;
  wire tmp38173;
  wire tmp38174;
  wire tmp38175;
  wire tmp38176;
  wire tmp38177;
  wire tmp38178;
  wire tmp38179;
  wire tmp38180;
  wire tmp38181;
  wire tmp38182;
  wire tmp38183;
  wire tmp38184;
  wire tmp38185;
  wire tmp38186;
  wire tmp38187;
  wire tmp38188;
  wire tmp38189;
  wire tmp38190;
  wire tmp38191;
  wire tmp38192;
  wire tmp38193;
  wire tmp38194;
  wire tmp38195;
  wire tmp38196;
  wire tmp38197;
  wire tmp38198;
  wire tmp38199;
  wire tmp38200;
  wire tmp38201;
  wire tmp38202;
  wire tmp38203;
  wire tmp38204;
  wire tmp38205;
  wire tmp38206;
  wire tmp38207;
  wire tmp38208;
  wire tmp38209;
  wire tmp38210;
  wire tmp38211;
  wire tmp38212;
  wire tmp38213;
  wire tmp38214;
  wire tmp38215;
  wire tmp38216;
  wire tmp38217;
  wire tmp38218;
  wire tmp38219;
  wire tmp38220;
  wire tmp38221;
  wire tmp38222;
  wire tmp38223;
  wire tmp38224;
  wire tmp38225;
  wire tmp38226;
  wire tmp38227;
  wire tmp38228;
  wire tmp38229;
  wire tmp38230;
  wire tmp38231;
  wire tmp38232;
  wire tmp38233;
  wire tmp38234;
  wire tmp38235;
  wire tmp38236;
  wire tmp38237;
  wire tmp38238;
  wire tmp38239;
  wire tmp38240;
  wire tmp38241;
  wire tmp38242;
  wire tmp38243;
  wire tmp38244;
  wire tmp38245;
  wire tmp38246;
  wire tmp38247;
  wire tmp38248;
  wire tmp38249;
  wire tmp38250;
  wire tmp38251;
  wire tmp38252;
  wire tmp38253;
  wire tmp38254;
  wire tmp38255;
  wire tmp38256;
  wire tmp38257;
  wire tmp38258;
  wire tmp38259;
  wire tmp38260;
  wire tmp38261;
  wire tmp38262;
  wire tmp38263;
  wire tmp38264;
  wire tmp38265;
  wire tmp38266;
  wire tmp38267;
  wire tmp38268;
  wire tmp38269;
  wire tmp38270;
  wire tmp38271;
  wire tmp38272;
  wire tmp38273;
  wire tmp38274;
  wire tmp38275;
  wire tmp38276;
  wire tmp38277;
  wire tmp38278;
  wire tmp38279;
  wire tmp38280;
  wire tmp38281;
  wire tmp38282;
  wire tmp38283;
  wire tmp38284;
  wire tmp38285;
  wire tmp38286;
  wire tmp38287;
  wire tmp38288;
  wire tmp38289;
  wire tmp38290;
  wire tmp38291;
  wire tmp38292;
  wire tmp38293;
  wire tmp38294;
  wire tmp38295;
  wire tmp38296;
  wire tmp38297;
  wire tmp38298;
  wire tmp38299;
  wire tmp38300;
  wire tmp38301;
  wire tmp38302;
  wire tmp38303;
  wire tmp38304;
  wire tmp38305;
  wire tmp38306;
  wire tmp38307;
  wire tmp38308;
  wire tmp38309;
  wire tmp38310;
  wire tmp38311;
  wire tmp38312;
  wire tmp38313;
  wire tmp38314;
  wire tmp38315;
  wire tmp38316;
  wire tmp38317;
  wire tmp38318;
  wire tmp38319;
  wire tmp38320;
  wire tmp38321;
  wire tmp38322;
  wire tmp38323;
  wire tmp38324;
  wire tmp38325;
  wire tmp38326;
  wire tmp38327;
  wire tmp38328;
  wire tmp38329;
  wire tmp38330;
  wire tmp38331;
  wire tmp38332;
  wire tmp38333;
  wire tmp38334;
  wire tmp38335;
  wire tmp38336;
  wire tmp38337;
  wire tmp38338;
  wire tmp38339;
  wire tmp38340;
  wire tmp38341;
  wire tmp38342;
  wire tmp38343;
  wire tmp38344;
  wire tmp38345;
  wire tmp38346;
  wire tmp38347;
  wire tmp38348;
  wire tmp38349;
  wire tmp38350;
  wire tmp38351;
  wire tmp38352;
  wire tmp38353;
  wire tmp38354;
  wire tmp38355;
  wire tmp38356;
  wire tmp38357;
  wire tmp38358;
  wire tmp38359;
  wire tmp38360;
  wire tmp38361;
  wire tmp38362;
  wire tmp38363;
  wire tmp38364;
  wire tmp38365;
  wire tmp38366;
  wire tmp38367;
  wire tmp38368;
  wire tmp38369;
  wire tmp38370;
  wire tmp38371;
  wire tmp38372;
  wire tmp38373;
  wire tmp38374;
  wire tmp38375;
  wire tmp38376;
  wire tmp38377;
  wire tmp38378;
  wire tmp38379;
  wire tmp38380;
  wire tmp38381;
  wire tmp38382;
  wire tmp38383;
  wire tmp38384;
  wire tmp38385;
  wire tmp38386;
  wire tmp38387;
  wire tmp38388;
  wire tmp38389;
  wire tmp38390;
  wire tmp38391;
  wire tmp38392;
  wire tmp38393;
  wire tmp38394;
  wire tmp38395;
  wire tmp38396;
  wire tmp38397;
  wire tmp38398;
  wire tmp38399;
  wire tmp38400;
  wire tmp38401;
  wire tmp38402;
  wire tmp38403;
  wire tmp38404;
  wire tmp38405;
  wire tmp38406;
  wire tmp38407;
  wire tmp38408;
  wire tmp38409;
  wire tmp38410;
  wire tmp38411;
  wire tmp38412;
  wire tmp38413;
  wire tmp38414;
  wire tmp38415;
  wire tmp38416;
  wire tmp38417;
  wire tmp38418;
  wire tmp38419;
  wire tmp38420;
  wire tmp38421;
  wire tmp38422;
  wire tmp38423;
  wire tmp38424;
  wire tmp38425;
  wire tmp38426;
  wire tmp38427;
  wire tmp38428;
  wire tmp38429;
  wire tmp38430;
  wire tmp38431;
  wire tmp38432;
  wire tmp38433;
  wire tmp38434;
  wire tmp38435;
  wire tmp38436;
  wire tmp38437;
  wire tmp38438;
  wire tmp38439;
  wire tmp38440;
  wire tmp38441;
  wire tmp38442;
  wire tmp38443;
  wire tmp38444;
  wire tmp38445;
  wire tmp38446;
  wire tmp38447;
  wire tmp38448;
  wire tmp38449;
  wire tmp38450;
  wire tmp38451;
  wire tmp38452;
  wire tmp38453;
  wire tmp38454;
  wire tmp38455;
  wire tmp38456;
  wire tmp38457;
  wire tmp38458;
  wire tmp38459;
  wire tmp38460;
  wire tmp38461;
  wire tmp38462;
  wire tmp38463;
  wire tmp38464;
  wire tmp38465;
  wire tmp38466;
  wire tmp38467;
  wire tmp38468;
  wire tmp38469;
  wire tmp38470;
  wire tmp38471;
  wire tmp38472;
  wire tmp38473;
  wire tmp38474;
  wire tmp38475;
  wire tmp38476;
  wire tmp38477;
  wire tmp38478;
  wire tmp38479;
  wire tmp38480;
  wire tmp38481;
  wire tmp38482;
  wire tmp38483;
  wire tmp38484;
  wire tmp38485;
  wire tmp38486;
  wire tmp38487;
  wire tmp38488;
  wire tmp38489;
  wire tmp38490;
  wire tmp38491;
  wire tmp38492;
  wire tmp38493;
  wire tmp38494;
  wire tmp38495;
  wire tmp38496;
  wire tmp38497;
  wire tmp38498;
  wire tmp38499;
  wire tmp38500;
  wire tmp38501;
  wire tmp38502;
  wire tmp38503;
  wire tmp38504;
  wire tmp38505;
  wire tmp38506;
  wire tmp38507;
  wire tmp38508;
  wire tmp38509;
  wire tmp38510;
  wire tmp38511;
  wire tmp38512;
  wire tmp38513;
  wire tmp38514;
  wire tmp38515;
  wire tmp38516;
  wire tmp38517;
  wire tmp38518;
  wire tmp38519;
  wire tmp38520;
  wire tmp38521;
  wire tmp38522;
  wire tmp38523;
  wire tmp38524;
  wire tmp38525;
  wire tmp38526;
  wire tmp38527;
  wire tmp38528;
  wire tmp38529;
  wire tmp38530;
  wire tmp38531;
  wire tmp38532;
  wire tmp38533;
  wire tmp38534;
  wire tmp38535;
  wire tmp38536;
  wire tmp38537;
  wire tmp38538;
  wire tmp38539;
  wire tmp38540;
  wire tmp38541;
  wire tmp38542;
  wire tmp38543;
  wire tmp38544;
  wire tmp38545;
  wire tmp38546;
  wire tmp38547;
  wire tmp38548;
  wire tmp38549;
  wire tmp38550;
  wire tmp38551;
  wire tmp38552;
  wire tmp38553;
  wire tmp38554;
  wire tmp38555;
  wire tmp38556;
  wire tmp38557;
  wire tmp38558;
  wire tmp38559;
  wire tmp38560;
  wire tmp38561;
  wire tmp38562;
  wire tmp38563;
  wire tmp38564;
  wire tmp38565;
  wire tmp38566;
  wire tmp38567;
  wire tmp38568;
  wire tmp38569;
  wire tmp38570;
  wire tmp38571;
  wire tmp38572;
  wire tmp38573;
  wire tmp38574;
  wire tmp38575;
  wire tmp38576;
  wire tmp38577;
  wire tmp38578;
  wire tmp38579;
  wire tmp38580;
  wire tmp38581;
  wire tmp38582;
  wire tmp38583;
  wire tmp38584;
  wire tmp38585;
  wire tmp38586;
  wire tmp38587;
  wire tmp38588;
  wire tmp38589;
  wire tmp38590;
  wire tmp38591;
  wire tmp38592;
  wire tmp38593;
  wire tmp38594;
  wire tmp38595;
  wire tmp38596;
  wire tmp38597;
  wire tmp38598;
  wire tmp38599;
  wire tmp38600;
  wire tmp38601;
  wire tmp38602;
  wire tmp38603;
  wire tmp38604;
  wire tmp38605;
  wire tmp38606;
  wire tmp38607;
  wire tmp38608;
  wire tmp38609;
  wire tmp38610;
  wire tmp38611;
  wire tmp38612;
  wire tmp38613;
  wire tmp38614;
  wire tmp38615;
  wire tmp38616;
  wire tmp38617;
  wire tmp38618;
  wire tmp38619;
  wire tmp38620;
  wire tmp38621;
  wire tmp38622;
  wire tmp38623;
  wire tmp38624;
  wire tmp38625;
  wire tmp38626;
  wire tmp38627;
  wire tmp38628;
  wire tmp38629;
  wire tmp38630;
  wire tmp38631;
  wire tmp38632;
  wire tmp38633;
  wire tmp38634;
  wire tmp38635;
  wire tmp38636;
  wire tmp38637;
  wire tmp38638;
  wire tmp38639;
  wire tmp38640;
  wire tmp38641;
  wire tmp38642;
  wire tmp38643;
  wire tmp38644;
  wire tmp38645;
  wire tmp38646;
  wire tmp38647;
  wire tmp38648;
  wire tmp38649;
  wire tmp38650;
  wire tmp38651;
  wire tmp38652;
  wire tmp38653;
  wire tmp38654;
  wire tmp38655;
  wire tmp38656;
  wire tmp38657;
  wire tmp38658;
  wire tmp38659;
  wire tmp38660;
  wire tmp38661;
  wire tmp38662;
  wire tmp38663;
  wire tmp38664;
  wire tmp38665;
  wire tmp38666;
  wire tmp38667;
  wire tmp38668;
  wire tmp38669;
  wire tmp38670;
  wire tmp38671;
  wire tmp38672;
  wire tmp38673;
  wire tmp38674;
  wire tmp38675;
  wire tmp38676;
  wire tmp38677;
  wire tmp38678;
  wire tmp38679;
  wire tmp38680;
  wire tmp38681;
  wire tmp38682;
  wire tmp38683;
  wire tmp38684;
  wire tmp38685;
  wire tmp38686;
  wire tmp38687;
  wire tmp38688;
  wire tmp38689;
  wire tmp38690;
  wire tmp38691;
  wire tmp38692;
  wire tmp38693;
  wire tmp38694;
  wire tmp38695;
  wire tmp38696;
  wire tmp38697;
  wire tmp38698;
  wire tmp38699;
  wire tmp38700;
  wire tmp38701;
  wire tmp38702;
  wire tmp38703;
  wire tmp38704;
  wire tmp38705;
  wire tmp38706;
  wire tmp38707;
  wire tmp38708;
  wire tmp38709;
  wire tmp38710;
  wire tmp38711;
  wire tmp38712;
  wire tmp38713;
  wire tmp38714;
  wire tmp38715;
  wire tmp38716;
  wire tmp38717;
  wire tmp38718;
  wire tmp38719;
  wire tmp38720;
  wire tmp38721;
  wire tmp38722;
  wire tmp38723;
  wire tmp38724;
  wire tmp38725;
  wire tmp38726;
  wire tmp38727;
  wire tmp38728;
  wire tmp38729;
  wire tmp38730;
  wire tmp38731;
  wire tmp38732;
  wire tmp38733;
  wire tmp38734;
  wire tmp38735;
  wire tmp38736;
  wire tmp38737;
  wire tmp38738;
  wire tmp38739;
  wire tmp38740;
  wire tmp38741;
  wire tmp38742;
  wire tmp38743;
  wire tmp38744;
  wire tmp38745;
  wire tmp38746;
  wire tmp38747;
  wire tmp38748;
  wire tmp38749;
  wire tmp38750;
  wire tmp38751;
  wire tmp38752;
  wire tmp38753;
  wire tmp38754;
  wire tmp38755;
  wire tmp38756;
  wire tmp38757;
  wire tmp38758;
  wire tmp38759;
  wire tmp38760;
  wire tmp38761;
  wire tmp38762;
  wire tmp38763;
  wire tmp38764;
  wire tmp38765;
  wire tmp38766;
  wire tmp38767;
  wire tmp38768;
  wire tmp38769;
  wire tmp38770;
  wire tmp38771;
  wire tmp38772;
  wire tmp38773;
  wire tmp38774;
  wire tmp38775;
  wire tmp38776;
  wire tmp38777;
  wire tmp38778;
  wire tmp38779;
  wire tmp38780;
  wire tmp38781;
  wire tmp38782;
  wire tmp38783;
  wire tmp38784;
  wire tmp38785;
  wire tmp38786;
  wire tmp38787;
  wire tmp38788;
  wire tmp38789;
  wire tmp38790;
  wire tmp38791;
  wire tmp38792;
  wire tmp38793;
  wire tmp38794;
  wire tmp38795;
  wire tmp38796;
  wire tmp38797;
  wire tmp38798;
  wire tmp38799;
  wire tmp38800;
  wire tmp38801;
  wire tmp38802;
  wire tmp38803;
  wire tmp38804;
  wire tmp38805;
  wire tmp38806;
  wire tmp38807;
  wire tmp38808;
  wire tmp38809;
  wire tmp38810;
  wire tmp38811;
  wire tmp38812;
  wire tmp38813;
  wire tmp38814;
  wire tmp38815;
  wire tmp38816;
  wire tmp38817;
  wire tmp38818;
  wire tmp38819;
  wire tmp38820;
  wire tmp38821;
  wire tmp38822;
  wire tmp38823;
  wire tmp38824;
  wire tmp38825;
  wire tmp38826;
  wire tmp38827;
  wire tmp38828;
  wire tmp38829;
  wire tmp38830;
  wire tmp38831;
  wire tmp38832;
  wire tmp38833;
  wire tmp38834;
  wire tmp38835;
  wire tmp38836;
  wire tmp38837;
  wire tmp38838;
  wire tmp38839;
  wire tmp38840;
  wire tmp38841;
  wire tmp38842;
  wire tmp38843;
  wire tmp38844;
  wire tmp38845;
  wire tmp38846;
  wire tmp38847;
  wire tmp38848;
  wire tmp38849;
  wire tmp38850;
  wire tmp38851;
  wire tmp38852;
  wire tmp38853;
  wire tmp38854;
  wire tmp38855;
  wire tmp38856;
  wire tmp38857;
  wire tmp38858;
  wire tmp38859;
  wire tmp38860;
  wire tmp38861;
  wire tmp38862;
  wire tmp38863;
  wire tmp38864;
  wire tmp38865;
  wire tmp38866;
  wire tmp38867;
  wire tmp38868;
  wire tmp38869;
  wire tmp38870;
  wire tmp38871;
  wire tmp38872;
  wire tmp38873;
  wire tmp38874;
  wire tmp38875;
  wire tmp38876;
  wire tmp38877;
  wire tmp38878;
  wire tmp38879;
  wire tmp38880;
  wire tmp38881;
  wire tmp38882;
  wire tmp38883;
  wire tmp38884;
  wire tmp38885;
  wire tmp38886;
  wire tmp38887;
  wire tmp38888;
  wire tmp38889;
  wire tmp38890;
  wire tmp38891;
  wire tmp38892;
  wire tmp38893;
  wire tmp38894;
  wire tmp38895;
  wire tmp38896;
  wire tmp38897;
  wire tmp38898;
  wire tmp38899;
  wire tmp38900;
  wire tmp38901;
  wire tmp38902;
  wire tmp38903;
  wire tmp38904;
  wire tmp38905;
  wire tmp38906;
  wire tmp38907;
  wire tmp38908;
  wire tmp38909;
  wire tmp38910;
  wire tmp38911;
  wire tmp38912;
  wire tmp38913;
  wire tmp38914;
  wire tmp38915;
  wire tmp38916;
  wire tmp38917;
  wire tmp38918;
  wire tmp38919;
  wire tmp38920;
  wire tmp38921;
  wire tmp38922;
  wire tmp38923;
  wire tmp38924;
  wire tmp38925;
  wire tmp38926;
  wire tmp38927;
  wire tmp38928;
  wire tmp38929;
  wire tmp38930;
  wire tmp38931;
  wire tmp38932;
  wire tmp38933;
  wire tmp38934;
  wire tmp38935;
  wire tmp38936;
  wire tmp38937;
  wire tmp38938;
  wire tmp38939;
  wire tmp38940;
  wire tmp38941;
  wire tmp38942;
  wire tmp38943;
  wire tmp38944;
  wire tmp38945;
  wire tmp38946;
  wire tmp38947;
  wire tmp38948;
  wire tmp38949;
  wire tmp38950;
  wire tmp38951;
  wire tmp38952;
  wire tmp38953;
  wire tmp38954;
  wire tmp38955;
  wire tmp38956;
  wire tmp38957;
  wire tmp38958;
  wire tmp38959;
  wire tmp38960;
  wire tmp38961;
  wire tmp38962;
  wire tmp38963;
  wire tmp38964;
  wire tmp38965;
  wire tmp38966;
  wire tmp38967;
  wire tmp38968;
  wire tmp38969;
  wire tmp38970;
  wire tmp38971;
  wire tmp38972;
  wire tmp38973;
  wire tmp38974;
  wire tmp38975;
  wire tmp38976;
  wire tmp38977;
  wire tmp38978;
  wire tmp38979;
  wire tmp38980;
  wire tmp38981;
  wire tmp38982;
  wire tmp38983;
  wire tmp38984;
  wire tmp38985;
  wire tmp38986;
  wire tmp38987;
  wire tmp38988;
  wire tmp38989;
  wire tmp38990;
  wire tmp38991;
  wire tmp38992;
  wire tmp38993;
  wire tmp38994;
  wire tmp38995;
  wire tmp38996;
  wire tmp38997;
  wire tmp38998;
  wire tmp38999;
  wire tmp39000;
  wire tmp39001;
  wire tmp39002;
  wire tmp39003;
  wire tmp39004;
  wire tmp39005;
  wire tmp39006;
  wire tmp39007;
  wire tmp39008;
  wire tmp39009;
  wire tmp39010;
  wire tmp39011;
  wire tmp39012;
  wire tmp39013;
  wire tmp39014;
  wire tmp39015;
  wire tmp39016;
  wire tmp39017;
  wire tmp39018;
  wire tmp39019;
  wire tmp39020;
  wire tmp39021;
  wire tmp39022;
  wire tmp39023;
  wire tmp39024;
  wire tmp39025;
  wire tmp39026;
  wire tmp39027;
  wire tmp39028;
  wire tmp39029;
  wire tmp39030;
  wire tmp39031;
  wire tmp39032;
  wire tmp39033;
  wire tmp39034;
  wire tmp39035;
  wire tmp39036;
  wire tmp39037;
  wire tmp39038;
  wire tmp39039;
  wire tmp39040;
  wire tmp39041;
  wire tmp39042;
  wire tmp39043;
  wire tmp39044;
  wire tmp39045;
  wire tmp39046;
  wire tmp39047;
  wire tmp39048;
  wire tmp39049;
  wire tmp39050;
  wire tmp39051;
  wire tmp39052;
  wire tmp39053;
  wire tmp39054;
  wire tmp39055;
  wire tmp39056;
  wire tmp39057;
  wire tmp39058;
  wire tmp39059;
  wire tmp39060;
  wire tmp39061;
  wire tmp39062;
  wire tmp39063;
  wire tmp39064;
  wire tmp39065;
  wire tmp39066;
  wire tmp39067;
  wire tmp39068;
  wire tmp39069;
  wire tmp39070;
  wire tmp39071;
  wire tmp39072;
  wire tmp39073;
  wire tmp39074;
  wire tmp39075;
  wire tmp39076;
  wire tmp39077;
  wire tmp39078;
  wire tmp39079;
  wire tmp39080;
  wire tmp39081;
  wire tmp39082;
  wire tmp39083;
  wire tmp39084;
  wire tmp39085;
  wire tmp39086;
  wire tmp39087;
  wire tmp39088;
  wire tmp39089;
  wire tmp39090;
  wire tmp39091;
  wire tmp39092;
  wire tmp39093;
  wire tmp39094;
  wire tmp39095;
  wire tmp39096;
  wire tmp39097;
  wire tmp39098;
  wire tmp39099;
  wire tmp39100;
  wire tmp39101;
  wire tmp39102;
  wire tmp39103;
  wire tmp39104;
  wire tmp39105;
  wire tmp39106;
  wire tmp39107;
  wire tmp39108;
  wire tmp39109;
  wire tmp39110;
  wire tmp39111;
  wire tmp39112;
  wire tmp39113;
  wire tmp39114;
  wire tmp39115;
  wire tmp39116;
  wire tmp39117;
  wire tmp39118;
  wire tmp39119;
  wire tmp39120;
  wire tmp39121;
  wire tmp39122;
  wire tmp39123;
  wire tmp39124;
  wire tmp39125;
  wire tmp39126;
  wire tmp39127;
  wire tmp39128;
  wire tmp39129;
  wire tmp39130;
  wire tmp39131;
  wire tmp39132;
  wire tmp39133;
  wire tmp39134;
  wire tmp39135;
  wire tmp39136;
  wire tmp39137;
  wire tmp39138;
  wire tmp39139;
  wire tmp39140;
  wire tmp39141;
  wire tmp39142;
  wire tmp39143;
  wire tmp39144;
  wire tmp39145;
  wire tmp39146;
  wire tmp39147;
  wire tmp39148;
  wire tmp39149;
  wire tmp39150;
  wire tmp39151;
  wire tmp39152;
  wire tmp39153;
  wire tmp39154;
  wire tmp39155;
  wire tmp39156;
  wire tmp39157;
  wire tmp39158;
  wire tmp39159;
  wire tmp39160;
  wire tmp39161;
  wire tmp39162;
  wire tmp39163;
  wire tmp39164;
  wire tmp39165;
  wire tmp39166;
  wire tmp39167;
  wire tmp39168;
  wire tmp39169;
  wire tmp39170;
  wire tmp39171;
  wire tmp39172;
  wire tmp39173;
  wire tmp39174;
  wire tmp39175;
  wire tmp39176;
  wire tmp39177;
  wire tmp39178;
  wire tmp39179;
  wire tmp39180;
  wire tmp39181;
  wire tmp39182;
  wire tmp39183;
  wire tmp39184;
  wire tmp39185;
  wire tmp39186;
  wire tmp39187;
  wire tmp39188;
  wire tmp39189;
  wire tmp39190;
  wire tmp39191;
  wire tmp39192;
  wire tmp39193;
  wire tmp39194;
  wire tmp39195;
  wire tmp39196;
  wire tmp39197;
  wire tmp39198;
  wire tmp39199;
  wire tmp39200;
  wire tmp39201;
  wire tmp39202;
  wire tmp39203;
  wire tmp39204;
  wire tmp39205;
  wire tmp39206;
  wire tmp39207;
  wire tmp39208;
  wire tmp39209;
  wire tmp39210;
  wire tmp39211;
  wire tmp39212;
  wire tmp39213;
  wire tmp39214;
  wire tmp39215;
  wire tmp39216;
  wire tmp39217;
  wire tmp39218;
  wire tmp39219;
  wire tmp39220;
  wire tmp39221;
  wire tmp39222;
  wire tmp39223;
  wire tmp39224;
  wire tmp39225;
  wire tmp39226;
  wire tmp39227;
  wire tmp39228;
  wire tmp39229;
  wire tmp39230;
  wire tmp39231;
  wire tmp39232;
  wire tmp39233;
  wire tmp39234;
  wire tmp39235;
  wire tmp39236;
  wire tmp39237;
  wire tmp39238;
  wire tmp39239;
  wire tmp39240;
  wire tmp39241;
  wire tmp39242;
  wire tmp39243;
  wire tmp39244;
  wire tmp39245;
  wire tmp39246;
  wire tmp39247;
  wire tmp39248;
  wire tmp39249;
  wire tmp39250;
  wire tmp39251;
  wire tmp39252;
  wire tmp39253;
  wire tmp39254;
  wire tmp39255;
  wire tmp39256;
  wire tmp39257;
  wire tmp39258;
  wire tmp39259;
  wire tmp39260;
  wire tmp39261;
  wire tmp39262;
  wire tmp39263;
  wire tmp39264;
  wire tmp39265;
  wire tmp39266;
  wire tmp39267;
  wire tmp39268;
  wire tmp39269;
  wire tmp39270;
  wire tmp39271;
  wire tmp39272;
  wire tmp39273;
  wire tmp39274;
  wire tmp39275;
  wire tmp39276;
  wire tmp39277;
  wire tmp39278;
  wire tmp39279;
  wire tmp39280;
  wire tmp39281;
  wire tmp39282;
  wire tmp39283;
  wire tmp39284;
  wire tmp39285;
  wire tmp39286;
  wire tmp39287;
  wire tmp39288;
  wire tmp39289;
  wire tmp39290;
  wire tmp39291;
  wire tmp39292;
  wire tmp39293;
  wire tmp39294;
  wire tmp39295;
  wire tmp39296;
  wire tmp39297;
  wire tmp39298;
  wire tmp39299;
  wire tmp39300;
  wire tmp39301;
  wire tmp39302;
  wire tmp39303;
  wire tmp39304;
  wire tmp39305;
  wire tmp39306;
  wire tmp39307;
  wire tmp39308;
  wire tmp39309;
  wire tmp39310;
  wire tmp39311;
  wire tmp39312;
  wire tmp39313;
  wire tmp39314;
  wire tmp39315;
  wire tmp39316;
  wire tmp39317;
  wire tmp39318;
  wire tmp39319;
  wire tmp39320;
  wire tmp39321;
  wire tmp39322;
  wire tmp39323;
  wire tmp39324;
  wire tmp39325;
  wire tmp39326;
  wire tmp39327;
  wire tmp39328;
  wire tmp39329;
  wire tmp39330;
  wire tmp39331;
  wire tmp39332;
  wire tmp39333;
  wire tmp39334;
  wire tmp39335;
  wire tmp39336;
  wire tmp39337;
  wire tmp39338;
  wire tmp39339;
  wire tmp39340;
  wire tmp39341;
  wire tmp39342;
  wire tmp39343;
  wire tmp39344;
  wire tmp39345;
  wire tmp39346;
  wire tmp39347;
  wire tmp39348;
  wire tmp39349;
  wire tmp39350;
  wire tmp39351;
  wire tmp39352;
  wire tmp39353;
  wire tmp39354;
  wire tmp39355;
  wire tmp39356;
  wire tmp39357;
  wire tmp39358;
  wire tmp39359;
  wire tmp39360;
  wire tmp39361;
  wire tmp39362;
  wire tmp39363;
  wire tmp39364;
  wire tmp39365;
  wire tmp39366;
  wire tmp39367;
  wire tmp39368;
  wire tmp39369;
  wire tmp39370;
  wire tmp39371;
  wire tmp39372;
  wire tmp39373;
  wire tmp39374;
  wire tmp39375;
  wire tmp39376;
  wire tmp39377;
  wire tmp39378;
  wire tmp39379;
  wire tmp39380;
  wire tmp39381;
  wire tmp39382;
  wire tmp39383;
  wire tmp39384;
  wire tmp39385;
  wire tmp39386;
  wire tmp39387;
  wire tmp39388;
  wire tmp39389;
  wire tmp39390;
  wire tmp39391;
  wire tmp39392;
  wire tmp39393;
  wire tmp39394;
  wire tmp39395;
  wire tmp39396;
  wire tmp39397;
  wire tmp39398;
  wire tmp39399;
  wire tmp39400;
  wire tmp39401;
  wire tmp39402;
  wire tmp39403;
  wire tmp39404;
  wire tmp39405;
  wire tmp39406;
  wire tmp39407;
  wire tmp39408;
  wire tmp39409;
  wire tmp39410;
  wire tmp39411;
  wire tmp39412;
  wire tmp39413;
  wire tmp39414;
  wire tmp39415;
  wire tmp39416;
  wire tmp39417;
  wire tmp39418;
  wire tmp39419;
  wire tmp39420;
  wire tmp39421;
  wire tmp39422;
  wire tmp39423;
  wire tmp39424;
  wire tmp39425;
  wire tmp39426;
  wire tmp39427;
  wire tmp39428;
  wire tmp39429;
  wire tmp39430;
  wire tmp39431;
  wire tmp39432;
  wire tmp39433;
  wire tmp39434;
  wire tmp39435;
  wire tmp39436;
  wire tmp39437;
  wire tmp39438;
  wire tmp39439;
  wire tmp39440;
  wire tmp39441;
  wire tmp39442;
  wire tmp39443;
  wire tmp39444;
  wire tmp39445;
  wire tmp39446;
  wire tmp39447;
  wire tmp39448;
  wire tmp39449;
  wire tmp39450;
  wire tmp39451;
  wire tmp39452;
  wire tmp39453;
  wire tmp39454;
  wire tmp39455;
  wire tmp39456;
  wire tmp39457;
  wire tmp39458;
  wire tmp39459;
  wire tmp39460;
  wire tmp39461;
  wire tmp39462;
  wire tmp39463;
  wire tmp39464;
  wire tmp39465;
  wire tmp39466;
  wire tmp39467;
  wire tmp39468;
  wire tmp39469;
  wire tmp39470;
  wire tmp39471;
  wire tmp39472;
  wire tmp39473;
  wire tmp39474;
  wire tmp39475;
  wire tmp39476;
  wire tmp39477;
  wire tmp39478;
  wire tmp39479;
  wire tmp39480;
  wire tmp39481;
  wire tmp39482;
  wire tmp39483;
  wire tmp39484;
  wire tmp39485;
  wire tmp39486;
  wire tmp39487;
  wire tmp39488;
  wire tmp39489;
  wire tmp39490;
  wire tmp39491;
  wire tmp39492;
  wire tmp39493;
  wire tmp39494;
  wire tmp39495;
  wire tmp39496;
  wire tmp39497;
  wire tmp39498;
  wire tmp39499;
  wire tmp39500;
  wire tmp39501;
  wire tmp39502;
  wire tmp39503;
  wire tmp39504;
  wire tmp39505;
  wire tmp39506;
  wire tmp39507;
  wire tmp39508;
  wire tmp39509;
  wire tmp39510;
  wire tmp39511;
  wire tmp39512;
  wire tmp39513;
  wire tmp39514;
  wire tmp39515;
  wire tmp39516;
  wire tmp39517;
  wire tmp39518;
  wire tmp39519;
  wire tmp39520;
  wire tmp39521;
  wire tmp39522;
  wire tmp39523;
  wire tmp39524;
  wire tmp39525;
  wire tmp39526;
  wire tmp39527;
  wire tmp39528;
  wire tmp39529;
  wire tmp39530;
  wire tmp39531;
  wire tmp39532;
  wire tmp39533;
  wire tmp39534;
  wire tmp39535;
  wire tmp39536;
  wire tmp39537;
  wire tmp39538;
  wire tmp39539;
  wire tmp39540;
  wire tmp39541;
  wire tmp39542;
  wire tmp39543;
  wire tmp39544;
  wire tmp39545;
  wire tmp39546;
  wire tmp39547;
  wire tmp39548;
  wire tmp39549;
  wire tmp39550;
  wire tmp39551;
  wire tmp39552;
  wire tmp39553;
  wire tmp39554;
  wire tmp39555;
  wire tmp39556;
  wire tmp39557;
  wire tmp39558;
  wire tmp39559;
  wire tmp39560;
  wire tmp39561;
  wire tmp39562;
  wire tmp39563;
  wire tmp39564;
  wire tmp39565;
  wire tmp39566;
  wire tmp39567;
  wire tmp39568;
  wire tmp39569;
  wire tmp39570;
  wire tmp39571;
  wire tmp39572;
  wire tmp39573;
  wire tmp39574;
  wire tmp39575;
  wire tmp39576;
  wire tmp39577;
  wire tmp39578;
  wire tmp39579;
  wire tmp39580;
  wire tmp39581;
  wire tmp39582;
  wire tmp39583;
  wire tmp39584;
  wire tmp39585;
  wire tmp39586;
  wire tmp39587;
  wire tmp39588;
  wire tmp39589;
  wire tmp39590;
  wire tmp39591;
  wire tmp39592;
  wire tmp39593;
  wire tmp39594;
  wire tmp39595;
  wire tmp39596;
  wire tmp39597;
  wire tmp39598;
  wire tmp39599;
  wire tmp39600;
  wire tmp39601;
  wire tmp39602;
  wire tmp39603;
  wire tmp39604;
  wire tmp39605;
  wire tmp39606;
  wire tmp39607;
  wire tmp39608;
  wire tmp39609;
  wire tmp39610;
  wire tmp39611;
  wire tmp39612;
  wire tmp39613;
  wire tmp39614;
  wire tmp39615;
  wire tmp39616;
  wire tmp39617;
  wire tmp39618;
  wire tmp39619;
  wire tmp39620;
  wire tmp39621;
  wire tmp39622;
  wire tmp39623;
  wire tmp39624;
  wire tmp39625;
  wire tmp39626;
  wire tmp39627;
  wire tmp39628;
  wire tmp39629;
  wire tmp39630;
  wire tmp39631;
  wire tmp39632;
  wire tmp39633;
  wire tmp39634;
  wire tmp39635;
  wire tmp39636;
  wire tmp39637;
  wire tmp39638;
  wire tmp39639;
  wire tmp39640;
  wire tmp39641;
  wire tmp39642;
  wire tmp39643;
  wire tmp39644;
  wire tmp39645;
  wire tmp39646;
  wire tmp39647;
  wire tmp39648;
  wire tmp39649;
  wire tmp39650;
  wire tmp39651;
  wire tmp39652;
  wire tmp39653;
  wire tmp39654;
  wire tmp39655;
  wire tmp39656;
  wire tmp39657;
  wire tmp39658;
  wire tmp39659;
  wire tmp39660;
  wire tmp39661;
  wire tmp39662;
  wire tmp39663;
  wire tmp39664;
  wire tmp39665;
  wire tmp39666;
  wire tmp39667;
  wire tmp39668;
  wire tmp39669;
  wire tmp39670;
  wire tmp39671;
  wire tmp39672;
  wire tmp39673;
  wire tmp39674;
  wire tmp39675;
  wire tmp39676;
  wire tmp39677;
  wire tmp39678;
  wire tmp39679;
  wire tmp39680;
  wire tmp39681;
  wire tmp39682;
  wire tmp39683;
  wire tmp39684;
  wire tmp39685;
  wire tmp39686;
  wire tmp39687;
  wire tmp39688;
  wire tmp39689;
  wire tmp39690;
  wire tmp39691;
  wire tmp39692;
  wire tmp39693;
  wire tmp39694;
  wire tmp39695;
  wire tmp39696;
  wire tmp39697;
  wire tmp39698;
  wire tmp39699;
  wire tmp39700;
  wire tmp39701;
  wire tmp39702;
  wire tmp39703;
  wire tmp39704;
  wire tmp39705;
  wire tmp39706;
  wire tmp39707;
  wire tmp39708;
  wire tmp39709;
  wire tmp39710;
  wire tmp39711;
  wire tmp39712;
  wire tmp39713;
  wire tmp39714;
  wire tmp39715;
  wire tmp39716;
  wire tmp39717;
  wire tmp39718;
  wire tmp39719;
  wire tmp39720;
  wire tmp39721;
  wire tmp39722;
  wire tmp39723;
  wire tmp39724;
  wire tmp39725;
  wire tmp39726;
  wire tmp39727;
  wire tmp39728;
  wire tmp39729;
  wire tmp39730;
  wire tmp39731;
  wire tmp39732;
  wire tmp39733;
  wire tmp39734;
  wire tmp39735;
  wire tmp39736;
  wire tmp39737;
  wire tmp39738;
  wire tmp39739;
  wire tmp39740;
  wire tmp39741;
  wire tmp39742;
  wire tmp39743;
  wire tmp39744;
  wire tmp39745;
  wire tmp39746;
  wire tmp39747;
  wire tmp39748;
  wire tmp39749;
  wire tmp39750;
  wire tmp39751;
  wire tmp39752;
  wire tmp39753;
  wire tmp39754;
  wire tmp39755;
  wire tmp39756;
  wire tmp39757;
  wire tmp39758;
  wire tmp39759;
  wire tmp39760;
  wire tmp39761;
  wire tmp39762;
  wire tmp39763;
  wire tmp39764;
  wire tmp39765;
  wire tmp39766;
  wire tmp39767;
  wire tmp39768;
  wire tmp39769;
  wire tmp39770;
  wire tmp39771;
  wire tmp39772;
  wire tmp39773;
  wire tmp39774;
  wire tmp39775;
  wire tmp39776;
  wire tmp39777;
  wire tmp39778;
  wire tmp39779;
  wire tmp39780;
  wire tmp39781;
  wire tmp39782;
  wire tmp39783;
  wire tmp39784;
  wire tmp39785;
  wire tmp39786;
  wire tmp39787;
  wire tmp39788;
  wire tmp39789;
  wire tmp39790;
  wire tmp39791;
  wire tmp39792;
  wire tmp39793;
  wire tmp39794;
  wire tmp39795;
  wire tmp39796;
  wire tmp39797;
  wire tmp39798;
  wire tmp39799;
  wire tmp39800;
  wire tmp39801;
  wire tmp39802;
  wire tmp39803;
  wire tmp39804;
  wire tmp39805;
  wire tmp39806;
  wire tmp39807;
  wire tmp39808;
  wire tmp39809;
  wire tmp39810;
  wire tmp39811;
  wire tmp39812;
  wire tmp39813;
  wire tmp39814;
  wire tmp39815;
  wire tmp39816;
  wire tmp39817;
  wire tmp39818;
  wire tmp39819;
  wire tmp39820;
  wire tmp39821;
  wire tmp39822;
  wire tmp39823;
  wire tmp39824;
  wire tmp39825;
  wire tmp39826;
  wire tmp39827;
  wire tmp39828;
  wire tmp39829;
  wire tmp39830;
  wire tmp39831;
  wire tmp39832;
  wire tmp39833;
  wire tmp39834;
  wire tmp39835;
  wire tmp39836;
  wire tmp39837;
  wire tmp39838;
  wire tmp39839;
  wire tmp39840;
  wire tmp39841;
  wire tmp39842;
  wire tmp39843;
  wire tmp39844;
  wire tmp39845;
  wire tmp39846;
  wire tmp39847;
  wire tmp39848;
  wire tmp39849;
  wire tmp39850;
  wire tmp39851;
  wire tmp39852;
  wire tmp39853;
  wire tmp39854;
  wire tmp39855;
  wire tmp39856;
  wire tmp39857;
  wire tmp39858;
  wire tmp39859;
  wire tmp39860;
  wire tmp39861;
  wire tmp39862;
  wire tmp39863;
  wire tmp39864;
  wire tmp39865;
  wire tmp39866;
  wire tmp39867;
  wire tmp39868;
  wire tmp39869;
  wire tmp39870;
  wire tmp39871;
  wire tmp39872;
  wire tmp39873;
  wire tmp39874;
  wire tmp39875;
  wire tmp39876;
  wire tmp39877;
  wire tmp39878;
  wire tmp39879;
  wire tmp39880;
  wire tmp39881;
  wire tmp39882;
  wire tmp39883;
  wire tmp39884;
  wire tmp39885;
  wire tmp39886;
  wire tmp39887;
  wire tmp39888;
  wire tmp39889;
  wire tmp39890;
  wire tmp39891;
  wire tmp39892;
  wire tmp39893;
  wire tmp39894;
  wire tmp39895;
  wire tmp39896;
  wire tmp39897;
  wire tmp39898;
  wire tmp39899;
  wire tmp39900;
  wire tmp39901;
  wire tmp39902;
  wire tmp39903;
  wire tmp39904;
  wire tmp39905;
  wire tmp39906;
  wire tmp39907;
  wire tmp39908;
  wire tmp39909;
  wire tmp39910;
  wire tmp39911;
  wire tmp39912;
  wire tmp39913;
  wire tmp39914;
  wire tmp39915;
  wire tmp39916;
  wire tmp39917;
  wire tmp39918;
  wire tmp39919;
  wire tmp39920;
  wire tmp39921;
  wire tmp39922;
  wire tmp39923;
  wire tmp39924;
  wire tmp39925;
  wire tmp39926;
  wire tmp39927;
  wire tmp39928;
  wire tmp39929;
  wire tmp39930;
  wire tmp39931;
  wire tmp39932;
  wire tmp39933;
  wire tmp39934;
  wire tmp39935;
  wire tmp39936;
  wire tmp39937;
  wire tmp39938;
  wire tmp39939;
  wire tmp39940;
  wire tmp39941;
  wire tmp39942;
  wire tmp39943;
  wire tmp39944;
  wire tmp39945;
  wire tmp39946;
  wire tmp39947;
  wire tmp39948;
  wire tmp39949;
  wire tmp39950;
  wire tmp39951;
  wire tmp39952;
  wire tmp39953;
  wire tmp39954;
  wire tmp39955;
  wire tmp39956;
  wire tmp39957;
  wire tmp39958;
  wire tmp39959;
  wire tmp39960;
  wire tmp39961;
  wire tmp39962;
  wire tmp39963;
  wire tmp39964;
  wire tmp39965;
  wire tmp39966;
  wire tmp39967;
  wire tmp39968;
  wire tmp39969;
  wire tmp39970;
  wire tmp39971;
  wire tmp39972;
  wire tmp39973;
  wire tmp39974;
  wire tmp39975;
  wire tmp39976;
  wire tmp39977;
  wire tmp39978;
  wire tmp39979;
  wire tmp39980;
  wire tmp39981;
  wire tmp39982;
  wire tmp39983;
  wire tmp39984;
  wire tmp39985;
  wire tmp39986;
  wire tmp39987;
  wire tmp39988;
  wire tmp39989;
  wire tmp39990;
  wire tmp39991;
  wire tmp39992;
  wire tmp39993;
  wire tmp39994;
  wire tmp39995;
  wire tmp39996;
  wire tmp39997;
  wire tmp39998;
  wire tmp39999;
  wire tmp40000;
  wire tmp40001;
  wire tmp40002;
  wire tmp40003;
  wire tmp40004;
  wire tmp40005;
  wire tmp40006;
  wire tmp40007;
  wire tmp40008;
  wire tmp40009;
  wire tmp40010;
  wire tmp40011;
  wire tmp40012;
  wire tmp40013;
  wire tmp40014;
  wire tmp40015;
  wire tmp40016;
  wire tmp40017;
  wire tmp40018;
  wire tmp40019;
  wire tmp40020;
  wire tmp40021;
  wire tmp40022;
  wire tmp40023;
  wire tmp40024;
  wire tmp40025;
  wire tmp40026;
  wire tmp40027;
  wire tmp40028;
  wire tmp40029;
  wire tmp40030;
  wire tmp40031;
  wire tmp40032;
  wire tmp40033;
  wire tmp40034;
  wire tmp40035;
  wire tmp40036;
  wire tmp40037;
  wire tmp40038;
  wire tmp40039;
  wire tmp40040;
  wire tmp40041;
  wire tmp40042;
  wire tmp40043;
  wire tmp40044;
  wire tmp40045;
  wire tmp40046;
  wire tmp40047;
  wire tmp40048;
  wire tmp40049;
  wire tmp40050;
  wire tmp40051;
  wire tmp40052;
  wire tmp40053;
  wire tmp40054;
  wire tmp40055;
  wire tmp40056;
  wire tmp40057;
  wire tmp40058;
  wire tmp40059;
  wire tmp40060;
  wire tmp40061;
  wire tmp40062;
  wire tmp40063;
  wire tmp40064;
  wire tmp40065;
  wire tmp40066;
  wire tmp40067;
  wire tmp40068;
  wire tmp40069;
  wire tmp40070;
  wire tmp40071;
  wire tmp40072;
  wire tmp40073;
  wire tmp40074;
  wire tmp40075;
  wire tmp40076;
  wire tmp40077;
  wire tmp40078;
  wire tmp40079;
  wire tmp40080;
  wire tmp40081;
  wire tmp40082;
  wire tmp40083;
  wire tmp40084;
  wire tmp40085;
  wire tmp40086;
  wire tmp40087;
  wire tmp40088;
  wire tmp40089;
  wire tmp40090;
  wire tmp40091;
  wire tmp40092;
  wire tmp40093;
  wire tmp40094;
  wire tmp40095;
  wire tmp40096;
  wire tmp40097;
  wire tmp40098;
  wire tmp40099;
  wire tmp40100;
  wire tmp40101;
  wire tmp40102;
  wire tmp40103;
  wire tmp40104;
  wire tmp40105;
  wire tmp40106;
  wire tmp40107;
  wire tmp40108;
  wire tmp40109;
  wire tmp40110;
  wire tmp40111;
  wire tmp40112;
  wire tmp40113;
  wire tmp40114;
  wire tmp40115;
  wire tmp40116;
  wire tmp40117;
  wire tmp40118;
  wire tmp40119;
  wire tmp40120;
  wire tmp40121;
  wire tmp40122;
  wire tmp40123;
  wire tmp40124;
  wire tmp40125;
  wire tmp40126;
  wire tmp40127;
  wire tmp40128;
  wire tmp40129;
  wire tmp40130;
  wire tmp40131;
  wire tmp40132;
  wire tmp40133;
  wire tmp40134;
  wire tmp40135;
  wire tmp40136;
  wire tmp40137;
  wire tmp40138;
  wire tmp40139;
  wire tmp40140;
  wire tmp40141;
  wire tmp40142;
  wire tmp40143;
  wire tmp40144;
  wire tmp40145;
  wire tmp40146;
  wire tmp40147;
  wire tmp40148;
  wire tmp40149;
  wire tmp40150;
  wire tmp40151;
  wire tmp40152;
  wire tmp40153;
  wire tmp40154;
  wire tmp40155;
  wire tmp40156;
  wire tmp40157;
  wire tmp40158;
  wire tmp40159;
  wire tmp40160;
  wire tmp40161;
  wire tmp40162;
  wire tmp40163;
  wire tmp40164;
  wire tmp40165;
  wire tmp40166;
  wire tmp40167;
  wire tmp40168;
  wire tmp40169;
  wire tmp40170;
  wire tmp40171;
  wire tmp40172;
  wire tmp40173;
  wire tmp40174;
  wire tmp40175;
  wire tmp40176;
  wire tmp40177;
  wire tmp40178;
  wire tmp40179;
  wire tmp40180;
  wire tmp40181;
  wire tmp40182;
  wire tmp40183;
  wire tmp40184;
  wire tmp40185;
  wire tmp40186;
  wire tmp40187;
  wire tmp40188;
  wire tmp40189;
  wire tmp40190;
  wire tmp40191;
  wire tmp40192;
  wire tmp40193;
  wire tmp40194;
  wire tmp40195;
  wire tmp40196;
  wire tmp40197;
  wire tmp40198;
  wire tmp40199;
  wire tmp40200;
  wire tmp40201;
  wire tmp40202;
  wire tmp40203;
  wire tmp40204;
  wire tmp40205;
  wire tmp40206;
  wire tmp40207;
  wire tmp40208;
  wire tmp40209;
  wire tmp40210;
  wire tmp40211;
  wire tmp40212;
  wire tmp40213;
  wire tmp40214;
  wire tmp40215;
  wire tmp40216;
  wire tmp40217;
  wire tmp40218;
  wire tmp40219;
  wire tmp40220;
  wire tmp40221;
  wire tmp40222;
  wire tmp40223;
  wire tmp40224;
  wire tmp40225;
  wire tmp40226;
  wire tmp40227;
  wire tmp40228;
  wire tmp40229;
  wire tmp40230;
  wire tmp40231;
  wire tmp40232;
  wire tmp40233;
  wire tmp40234;
  wire tmp40235;
  wire tmp40236;
  wire tmp40237;
  wire tmp40238;
  wire tmp40239;
  wire tmp40240;
  wire tmp40241;
  wire tmp40242;
  wire tmp40243;
  wire tmp40244;
  wire tmp40245;
  wire tmp40246;
  wire tmp40247;
  wire tmp40248;
  wire tmp40249;
  wire tmp40250;
  wire tmp40251;
  wire tmp40252;
  wire tmp40253;
  wire tmp40254;
  wire tmp40255;
  wire tmp40256;
  wire tmp40257;
  wire tmp40258;
  wire tmp40259;
  wire tmp40260;
  wire tmp40261;
  wire tmp40262;
  wire tmp40263;
  wire tmp40264;
  wire tmp40265;
  wire tmp40266;
  wire tmp40267;
  wire tmp40268;
  wire tmp40269;
  wire tmp40270;
  wire tmp40271;
  wire tmp40272;
  wire tmp40273;
  wire tmp40274;
  wire tmp40275;
  wire tmp40276;
  wire tmp40277;
  wire tmp40278;
  wire tmp40279;
  wire tmp40280;
  wire tmp40281;
  wire tmp40282;
  wire tmp40283;
  wire tmp40284;
  wire tmp40285;
  wire tmp40286;
  wire tmp40287;
  wire tmp40288;
  wire tmp40289;
  wire tmp40290;
  wire tmp40291;
  wire tmp40292;
  wire tmp40293;
  wire tmp40294;
  wire tmp40295;
  wire tmp40296;
  wire tmp40297;
  wire tmp40298;
  wire tmp40299;
  wire tmp40300;
  wire tmp40301;
  wire tmp40302;
  wire tmp40303;
  wire tmp40304;
  wire tmp40305;
  wire tmp40306;
  wire tmp40307;
  wire tmp40308;
  wire tmp40309;
  wire tmp40310;
  wire tmp40311;
  wire tmp40312;
  wire tmp40313;
  wire tmp40314;
  wire tmp40315;
  wire tmp40316;
  wire tmp40317;
  wire tmp40318;
  wire tmp40319;
  wire tmp40320;
  wire tmp40321;
  wire tmp40322;
  wire tmp40323;
  wire tmp40324;
  wire tmp40325;
  wire tmp40326;
  wire tmp40327;
  wire tmp40328;
  wire tmp40329;
  wire tmp40330;
  wire tmp40331;
  wire tmp40332;
  wire tmp40333;
  wire tmp40334;
  wire tmp40335;
  wire tmp40336;
  wire tmp40337;
  wire tmp40338;
  wire tmp40339;
  wire tmp40340;
  wire tmp40341;
  wire tmp40342;
  wire tmp40343;
  wire tmp40344;
  wire tmp40345;
  wire tmp40346;
  wire tmp40347;
  wire tmp40348;
  wire tmp40349;
  wire tmp40350;
  wire tmp40351;
  wire tmp40352;
  wire tmp40353;
  wire tmp40354;
  wire tmp40355;
  wire tmp40356;
  wire tmp40357;
  wire tmp40358;
  wire tmp40359;
  wire tmp40360;
  wire tmp40361;
  wire tmp40362;
  wire tmp40363;
  wire tmp40364;
  wire tmp40365;
  wire tmp40366;
  wire tmp40367;
  wire tmp40368;
  wire tmp40369;
  wire tmp40370;
  wire tmp40371;
  wire tmp40372;
  wire tmp40373;
  wire tmp40374;
  wire tmp40375;
  wire tmp40376;
  wire tmp40377;
  wire tmp40378;
  wire tmp40379;
  wire tmp40380;
  wire tmp40381;
  wire tmp40382;
  wire tmp40383;
  wire tmp40384;
  wire tmp40385;
  wire tmp40386;
  wire tmp40387;
  wire tmp40388;
  wire tmp40389;
  wire tmp40390;
  wire tmp40391;
  wire tmp40392;
  wire tmp40393;
  wire tmp40394;
  wire tmp40395;
  wire tmp40396;
  wire tmp40397;
  wire tmp40398;
  wire tmp40399;
  wire tmp40400;
  wire tmp40401;
  wire tmp40402;
  wire tmp40403;
  wire tmp40404;
  wire tmp40405;
  wire tmp40406;
  wire tmp40407;
  wire tmp40408;
  wire tmp40409;
  wire tmp40410;
  wire tmp40411;
  wire tmp40412;
  wire tmp40413;
  wire tmp40414;
  wire tmp40415;
  wire tmp40416;
  wire tmp40417;
  wire tmp40418;
  wire tmp40419;
  wire tmp40420;
  wire tmp40421;
  wire tmp40422;
  wire tmp40423;
  wire tmp40424;
  wire tmp40425;
  wire tmp40426;
  wire tmp40427;
  wire tmp40428;
  wire tmp40429;
  wire tmp40430;
  wire tmp40431;
  wire tmp40432;
  wire tmp40433;
  wire tmp40434;
  wire tmp40435;
  wire tmp40436;
  wire tmp40437;
  wire tmp40438;
  wire tmp40439;
  wire tmp40440;
  wire tmp40441;
  wire tmp40442;
  wire tmp40443;
  wire tmp40444;
  wire tmp40445;
  wire tmp40446;
  wire tmp40447;
  wire tmp40448;
  wire tmp40449;
  wire tmp40450;
  wire tmp40451;
  wire tmp40452;
  wire tmp40453;
  wire tmp40454;
  wire tmp40455;
  wire tmp40456;
  wire tmp40457;
  wire tmp40458;
  wire tmp40459;
  wire tmp40460;
  wire tmp40461;
  wire tmp40462;
  wire tmp40463;
  wire tmp40464;
  wire tmp40465;
  wire tmp40466;
  wire tmp40467;
  wire tmp40468;
  wire tmp40469;
  wire tmp40470;
  wire tmp40471;
  wire tmp40472;
  wire tmp40473;
  wire tmp40474;
  wire tmp40475;
  wire tmp40476;
  wire tmp40477;
  wire tmp40478;
  wire tmp40479;
  wire tmp40480;
  wire tmp40481;
  wire tmp40482;
  wire tmp40483;
  wire tmp40484;
  wire tmp40485;
  wire tmp40486;
  wire tmp40487;
  wire tmp40488;
  wire tmp40489;
  wire tmp40490;
  wire tmp40491;
  wire tmp40492;
  wire tmp40493;
  wire tmp40494;
  wire tmp40495;
  wire tmp40496;
  wire tmp40497;
  wire tmp40498;
  wire tmp40499;
  wire tmp40500;
  wire tmp40501;
  wire tmp40502;
  wire tmp40503;
  wire tmp40504;
  wire tmp40505;
  wire tmp40506;
  wire tmp40507;
  wire tmp40508;
  wire tmp40509;
  wire tmp40510;
  wire tmp40511;
  wire tmp40512;
  wire tmp40513;
  wire tmp40514;
  wire tmp40515;
  wire tmp40516;
  wire tmp40517;
  wire tmp40518;
  wire tmp40519;
  wire tmp40520;
  wire tmp40521;
  wire tmp40522;
  wire tmp40523;
  wire tmp40524;
  wire tmp40525;
  wire tmp40526;
  wire tmp40527;
  wire tmp40528;
  wire tmp40529;
  wire tmp40530;
  wire tmp40531;
  wire tmp40532;
  wire tmp40533;
  wire tmp40534;
  wire tmp40535;
  wire tmp40536;
  wire tmp40537;
  wire tmp40538;
  wire tmp40539;
  wire tmp40540;
  wire tmp40541;
  wire tmp40542;
  wire tmp40543;
  wire tmp40544;
  wire tmp40545;
  wire tmp40546;
  wire tmp40547;
  wire tmp40548;
  wire tmp40549;
  wire tmp40550;
  wire tmp40551;
  wire tmp40552;
  wire tmp40553;
  wire tmp40554;
  wire tmp40555;
  wire tmp40556;
  wire tmp40557;
  wire tmp40558;
  wire tmp40559;
  wire tmp40560;
  wire tmp40561;
  wire tmp40562;
  wire tmp40563;
  wire tmp40564;
  wire tmp40565;
  wire tmp40566;
  wire tmp40567;
  wire tmp40568;
  wire tmp40569;
  wire tmp40570;
  wire tmp40571;
  wire tmp40572;
  wire tmp40573;
  wire tmp40574;
  wire tmp40575;
  wire tmp40576;
  wire tmp40577;
  wire tmp40578;
  wire tmp40579;
  wire tmp40580;
  wire tmp40581;
  wire tmp40582;
  wire tmp40583;
  wire tmp40584;
  wire tmp40585;
  wire tmp40586;
  wire tmp40587;
  wire tmp40588;
  wire tmp40589;
  wire tmp40590;
  wire tmp40591;
  wire tmp40592;
  wire tmp40593;
  wire tmp40594;
  wire tmp40595;
  wire tmp40596;
  wire tmp40597;
  wire tmp40598;
  wire tmp40599;
  wire tmp40600;
  wire tmp40601;
  wire tmp40602;
  wire tmp40603;
  wire tmp40604;
  wire tmp40605;
  wire tmp40606;
  wire tmp40607;
  wire tmp40608;
  wire tmp40609;
  wire tmp40610;
  wire tmp40611;
  wire tmp40612;
  wire tmp40613;
  wire tmp40614;
  wire tmp40615;
  wire tmp40616;
  wire tmp40617;
  wire tmp40618;
  wire tmp40619;
  wire tmp40620;
  wire tmp40621;
  wire tmp40622;
  wire tmp40623;
  wire tmp40624;
  wire tmp40625;
  wire tmp40626;
  wire tmp40627;
  wire tmp40628;
  wire tmp40629;
  wire tmp40630;
  wire tmp40631;
  wire tmp40632;
  wire tmp40633;
  wire tmp40634;
  wire tmp40635;
  wire tmp40636;
  wire tmp40637;
  wire tmp40638;
  wire tmp40639;
  wire tmp40640;
  wire tmp40641;
  wire tmp40642;
  wire tmp40643;
  wire tmp40644;
  wire tmp40645;
  wire tmp40646;
  wire tmp40647;
  wire tmp40648;
  wire tmp40649;
  wire tmp40650;
  wire tmp40651;
  wire tmp40652;
  wire tmp40653;
  wire tmp40654;
  wire tmp40655;
  wire tmp40656;
  wire tmp40657;
  wire tmp40658;
  wire tmp40659;
  wire tmp40660;
  wire tmp40661;
  wire tmp40662;
  wire tmp40663;
  wire tmp40664;
  wire tmp40665;
  wire tmp40666;
  wire tmp40667;
  wire tmp40668;
  wire tmp40669;
  wire tmp40670;
  wire tmp40671;
  wire tmp40672;
  wire tmp40673;
  wire tmp40674;
  wire tmp40675;
  wire tmp40676;
  wire tmp40677;
  wire tmp40678;
  wire tmp40679;
  wire tmp40680;
  wire tmp40681;
  wire tmp40682;
  wire tmp40683;
  wire tmp40684;
  wire tmp40685;
  wire tmp40686;
  wire tmp40687;
  wire tmp40688;
  wire tmp40689;
  wire tmp40690;
  wire tmp40691;
  wire tmp40692;
  wire tmp40693;
  wire tmp40694;
  wire tmp40695;
  wire tmp40696;
  wire tmp40697;
  wire tmp40698;
  wire tmp40699;
  wire tmp40700;
  wire tmp40701;
  wire tmp40702;
  wire tmp40703;
  wire tmp40704;
  wire tmp40705;
  wire tmp40706;
  wire tmp40707;
  wire tmp40708;
  wire tmp40709;
  wire tmp40710;
  wire tmp40711;
  wire tmp40712;
  wire tmp40713;
  wire tmp40714;
  wire tmp40715;
  wire tmp40716;
  wire tmp40717;
  wire tmp40718;
  wire tmp40719;
  wire tmp40720;
  wire tmp40721;
  wire tmp40722;
  wire tmp40723;
  wire tmp40724;
  wire tmp40725;
  wire tmp40726;
  wire tmp40727;
  wire tmp40728;
  wire tmp40729;
  wire tmp40730;
  wire tmp40731;
  wire tmp40732;
  wire tmp40733;
  wire tmp40734;
  wire tmp40735;
  wire tmp40736;
  wire tmp40737;
  wire tmp40738;
  wire tmp40739;
  wire tmp40740;
  wire tmp40741;
  wire tmp40742;
  wire tmp40743;
  wire tmp40744;
  wire tmp40745;
  wire tmp40746;
  wire tmp40747;
  wire tmp40748;
  wire tmp40749;
  wire tmp40750;
  wire tmp40751;
  wire tmp40752;
  wire tmp40753;
  wire tmp40754;
  wire tmp40755;
  wire tmp40756;
  wire tmp40757;
  wire tmp40758;
  wire tmp40759;
  wire tmp40760;
  wire tmp40761;
  wire tmp40762;
  wire tmp40763;
  wire tmp40764;
  wire tmp40765;
  wire tmp40766;
  wire tmp40767;
  wire tmp40768;
  wire tmp40769;
  wire tmp40770;
  wire tmp40771;
  wire tmp40772;
  wire tmp40773;
  wire tmp40774;
  wire tmp40775;
  wire tmp40776;
  wire tmp40777;
  wire tmp40778;
  wire tmp40779;
  wire tmp40780;
  wire tmp40781;
  wire tmp40782;
  wire tmp40783;
  wire tmp40784;
  wire tmp40785;
  wire tmp40786;
  wire tmp40787;
  wire tmp40788;
  wire tmp40789;
  wire tmp40790;
  wire tmp40791;
  wire tmp40792;
  wire tmp40793;
  wire tmp40794;
  wire tmp40795;
  wire tmp40796;
  wire tmp40797;
  wire tmp40798;
  wire tmp40799;
  wire tmp40800;
  wire tmp40801;
  wire tmp40802;
  wire tmp40803;
  wire tmp40804;
  wire tmp40805;
  wire tmp40806;
  wire tmp40807;
  wire tmp40808;
  wire tmp40809;
  wire tmp40810;
  wire tmp40811;
  wire tmp40812;
  wire tmp40813;
  wire tmp40814;
  wire tmp40815;
  wire tmp40816;
  wire tmp40817;
  wire tmp40818;
  wire tmp40819;
  wire tmp40820;
  wire tmp40821;
  wire tmp40822;
  wire tmp40823;
  wire tmp40824;
  wire tmp40825;
  wire tmp40826;
  wire tmp40827;
  wire tmp40828;
  wire tmp40829;
  wire tmp40830;
  wire tmp40831;
  wire tmp40832;
  wire tmp40833;
  wire tmp40834;
  wire tmp40835;
  wire tmp40836;
  wire tmp40837;
  wire tmp40838;
  wire tmp40839;
  wire tmp40840;
  wire tmp40841;
  wire tmp40842;
  wire tmp40843;
  wire tmp40844;
  wire tmp40845;
  wire tmp40846;
  wire tmp40847;
  wire tmp40848;
  wire tmp40849;
  wire tmp40850;
  wire tmp40851;
  wire tmp40852;
  wire tmp40853;
  wire tmp40854;
  wire tmp40855;
  wire tmp40856;
  wire tmp40857;
  wire tmp40858;
  wire tmp40859;
  wire tmp40860;
  wire tmp40861;
  wire tmp40862;
  wire tmp40863;
  wire tmp40864;
  wire tmp40865;
  wire tmp40866;
  wire tmp40867;
  wire tmp40868;
  wire tmp40869;
  wire tmp40870;
  wire tmp40871;
  wire tmp40872;
  wire tmp40873;
  wire tmp40874;
  wire tmp40875;
  wire tmp40876;
  wire tmp40877;
  wire tmp40878;
  wire tmp40879;
  wire tmp40880;
  wire tmp40881;
  wire tmp40882;
  wire tmp40883;
  wire tmp40884;
  wire tmp40885;
  wire tmp40886;
  wire tmp40887;
  wire tmp40888;
  wire tmp40889;
  wire tmp40890;
  wire tmp40891;
  wire tmp40892;
  wire tmp40893;
  wire tmp40894;
  wire tmp40895;
  wire tmp40896;
  wire tmp40897;
  wire tmp40898;
  wire tmp40899;
  wire tmp40900;
  wire tmp40901;
  wire tmp40902;
  wire tmp40903;
  wire tmp40904;
  wire tmp40905;
  wire tmp40906;
  wire tmp40907;
  wire tmp40908;
  wire tmp40909;
  wire tmp40910;
  wire tmp40911;
  wire tmp40912;
  wire tmp40913;
  wire tmp40914;
  wire tmp40915;
  wire tmp40916;
  wire tmp40917;
  wire tmp40918;
  wire tmp40919;
  wire tmp40920;
  wire tmp40921;
  wire tmp40922;
  wire tmp40923;
  wire tmp40924;
  wire tmp40925;
  wire tmp40926;
  wire tmp40927;
  wire tmp40928;
  wire tmp40929;
  wire tmp40930;
  wire tmp40931;
  wire tmp40932;
  wire tmp40933;
  wire tmp40934;
  wire tmp40935;
  wire tmp40936;
  wire tmp40937;
  wire tmp40938;
  wire tmp40939;
  wire tmp40940;
  wire tmp40941;
  wire tmp40942;
  wire tmp40943;
  wire tmp40944;
  wire tmp40945;
  wire tmp40946;
  wire tmp40947;
  wire tmp40948;
  wire tmp40949;
  wire tmp40950;
  wire tmp40951;
  wire tmp40952;
  wire tmp40953;
  wire tmp40954;
  wire tmp40955;
  wire tmp40956;
  wire tmp40957;
  wire tmp40958;
  wire tmp40959;
  wire tmp40960;
  wire tmp40961;
  wire tmp40962;
  wire tmp40963;
  wire tmp40964;
  wire tmp40965;
  wire tmp40966;
  wire tmp40967;
  wire tmp40968;
  wire tmp40969;
  wire tmp40970;
  wire tmp40971;
  wire tmp40972;
  wire tmp40973;
  wire tmp40974;
  wire tmp40975;
  wire tmp40976;
  wire tmp40977;
  wire tmp40978;
  wire tmp40979;
  wire tmp40980;
  wire tmp40981;
  wire tmp40982;
  wire tmp40983;
  wire tmp40984;
  wire tmp40985;
  wire tmp40986;
  wire tmp40987;
  wire tmp40988;
  wire tmp40989;
  wire tmp40990;
  wire tmp40991;
  wire tmp40992;
  wire tmp40993;
  wire tmp40994;
  wire tmp40995;
  wire tmp40996;
  wire tmp40997;
  wire tmp40998;
  wire tmp40999;
  wire tmp41000;
  wire tmp41001;
  wire tmp41002;
  wire tmp41003;
  wire tmp41004;
  wire tmp41005;
  wire tmp41006;
  wire tmp41007;
  wire tmp41008;
  wire tmp41009;
  wire tmp41010;
  wire tmp41011;
  wire tmp41012;
  wire tmp41013;
  wire tmp41014;
  wire tmp41015;
  wire tmp41016;
  wire tmp41017;
  wire tmp41018;
  wire tmp41019;
  wire tmp41020;
  wire tmp41021;
  wire tmp41022;
  wire tmp41023;
  wire tmp41024;
  wire tmp41025;
  wire tmp41026;
  wire tmp41027;
  wire tmp41028;
  wire tmp41029;
  wire tmp41030;
  wire tmp41031;
  wire tmp41032;
  wire tmp41033;
  wire tmp41034;
  wire tmp41035;
  wire tmp41036;
  wire tmp41037;
  wire tmp41038;
  wire tmp41039;
  wire tmp41040;
  wire tmp41041;
  wire tmp41042;
  wire tmp41043;
  wire tmp41044;
  wire tmp41045;
  wire tmp41046;
  wire tmp41047;
  wire tmp41048;
  wire tmp41049;
  wire tmp41050;
  wire tmp41051;
  wire tmp41052;
  wire tmp41053;
  wire tmp41054;
  wire tmp41055;
  wire tmp41056;
  wire tmp41057;
  wire tmp41058;
  wire tmp41059;
  wire tmp41060;
  wire tmp41061;
  wire tmp41062;
  wire tmp41063;
  wire tmp41064;
  wire tmp41065;
  wire tmp41066;
  wire tmp41067;
  wire tmp41068;
  wire tmp41069;
  wire tmp41070;
  wire tmp41071;
  wire tmp41072;
  wire tmp41073;
  wire tmp41074;
  wire tmp41075;
  wire tmp41076;
  wire tmp41077;
  wire tmp41078;
  wire tmp41079;
  wire tmp41080;
  wire tmp41081;
  wire tmp41082;
  wire tmp41083;
  wire tmp41084;
  wire tmp41085;
  wire tmp41086;
  wire tmp41087;
  wire tmp41088;
  wire tmp41089;
  wire tmp41090;
  wire tmp41091;
  wire tmp41092;
  wire tmp41093;
  wire tmp41094;
  wire tmp41095;
  wire tmp41096;
  wire tmp41097;
  wire tmp41098;
  wire tmp41099;
  wire tmp41100;
  wire tmp41101;
  wire tmp41102;
  wire tmp41103;
  wire tmp41104;
  wire tmp41105;
  wire tmp41106;
  wire tmp41107;
  wire tmp41108;
  wire tmp41109;
  wire tmp41110;
  wire tmp41111;
  wire tmp41112;
  wire tmp41113;
  wire tmp41114;
  wire tmp41115;
  wire tmp41116;
  wire tmp41117;
  wire tmp41118;
  wire tmp41119;
  wire tmp41120;
  wire tmp41121;
  wire tmp41122;
  wire tmp41123;
  wire tmp41124;
  wire tmp41125;
  wire tmp41126;
  wire tmp41127;
  wire tmp41128;
  wire tmp41129;
  wire tmp41130;
  wire tmp41131;
  wire tmp41132;
  wire tmp41133;
  wire tmp41134;
  wire tmp41135;
  wire tmp41136;
  wire tmp41137;
  wire tmp41138;
  wire tmp41139;
  wire tmp41140;
  wire tmp41141;
  wire tmp41142;
  wire tmp41143;
  wire tmp41144;
  wire tmp41145;
  wire tmp41146;
  wire tmp41147;
  wire tmp41148;
  wire tmp41149;
  wire tmp41150;
  wire tmp41151;
  wire tmp41152;
  wire tmp41153;
  wire tmp41154;
  wire tmp41155;
  wire tmp41156;
  wire tmp41157;
  wire tmp41158;
  wire tmp41159;
  wire tmp41160;
  wire tmp41161;
  wire tmp41162;
  wire tmp41163;
  wire tmp41164;
  wire tmp41165;
  wire tmp41166;
  wire tmp41167;
  wire tmp41168;
  wire tmp41169;
  wire tmp41170;
  wire tmp41171;
  wire tmp41172;
  wire tmp41173;
  wire tmp41174;
  wire tmp41175;
  wire tmp41176;
  wire tmp41177;
  wire tmp41178;
  wire tmp41179;
  wire tmp41180;
  wire tmp41181;
  wire tmp41182;
  wire tmp41183;
  wire tmp41184;
  wire tmp41185;
  wire tmp41186;
  wire tmp41187;
  wire tmp41188;
  wire tmp41189;
  wire tmp41190;
  wire tmp41191;
  wire tmp41192;
  wire tmp41193;
  wire tmp41194;
  wire tmp41195;
  wire tmp41196;
  wire tmp41197;
  wire tmp41198;
  wire tmp41199;
  wire tmp41200;
  wire tmp41201;
  wire tmp41202;
  wire tmp41203;
  wire tmp41204;
  wire tmp41205;
  wire tmp41206;
  wire tmp41207;
  wire tmp41208;
  wire tmp41209;
  wire tmp41210;
  wire tmp41211;
  wire tmp41212;
  wire tmp41213;
  wire tmp41214;
  wire tmp41215;
  wire tmp41216;
  wire tmp41217;
  wire tmp41218;
  wire tmp41219;
  wire tmp41220;
  wire tmp41221;
  wire tmp41222;
  wire tmp41223;
  wire tmp41224;
  wire tmp41225;
  wire tmp41226;
  wire tmp41227;
  wire tmp41228;
  wire tmp41229;
  wire tmp41230;
  wire tmp41231;
  wire tmp41232;
  wire tmp41233;
  wire tmp41234;
  wire tmp41235;
  wire tmp41236;
  wire tmp41237;
  wire tmp41238;
  wire tmp41239;
  wire tmp41240;
  wire tmp41241;
  wire tmp41242;
  wire tmp41243;
  wire tmp41244;
  wire tmp41245;
  wire tmp41246;
  wire tmp41247;
  wire tmp41248;
  wire tmp41249;
  wire tmp41250;
  wire tmp41251;
  wire tmp41252;
  wire tmp41253;
  wire tmp41254;
  wire tmp41255;
  wire tmp41256;
  wire tmp41257;
  wire tmp41258;
  wire tmp41259;
  wire tmp41260;
  wire tmp41261;
  wire tmp41262;
  wire tmp41263;
  wire tmp41264;
  wire tmp41265;
  wire tmp41266;
  wire tmp41267;
  wire tmp41268;
  wire tmp41269;
  wire tmp41270;
  wire tmp41271;
  wire tmp41272;
  wire tmp41273;
  wire tmp41274;
  wire tmp41275;
  wire tmp41276;
  wire tmp41277;
  wire tmp41278;
  wire tmp41279;
  wire tmp41280;
  wire tmp41281;
  wire tmp41282;
  wire tmp41283;
  wire tmp41284;
  wire tmp41285;
  wire tmp41286;
  wire tmp41287;
  wire tmp41288;
  wire tmp41289;
  wire tmp41290;
  wire tmp41291;
  wire tmp41292;
  wire tmp41293;
  wire tmp41294;
  wire tmp41295;
  wire tmp41296;
  wire tmp41297;
  wire tmp41298;
  wire tmp41299;
  wire tmp41300;
  wire tmp41301;
  wire tmp41302;
  wire tmp41303;
  wire tmp41304;
  wire tmp41305;
  wire tmp41306;
  wire tmp41307;
  wire tmp41308;
  wire tmp41309;
  wire tmp41310;
  wire tmp41311;
  wire tmp41312;
  wire tmp41313;
  wire tmp41314;
  wire tmp41315;
  wire tmp41316;
  wire tmp41317;
  wire tmp41318;
  wire tmp41319;
  wire tmp41320;
  wire tmp41321;
  wire tmp41322;
  wire tmp41323;
  wire tmp41324;
  wire tmp41325;
  wire tmp41326;
  wire tmp41327;
  wire tmp41328;
  wire tmp41329;
  wire tmp41330;
  wire tmp41331;
  wire tmp41332;
  wire tmp41333;
  wire tmp41334;
  wire tmp41335;
  wire tmp41336;
  wire tmp41337;
  wire tmp41338;
  wire tmp41339;
  wire tmp41340;
  wire tmp41341;
  wire tmp41342;
  wire tmp41343;
  wire tmp41344;
  wire tmp41345;
  wire tmp41346;
  wire tmp41347;
  wire tmp41348;
  wire tmp41349;
  wire tmp41350;
  wire tmp41351;
  wire tmp41352;
  wire tmp41353;
  wire tmp41354;
  wire tmp41355;
  wire tmp41356;
  wire tmp41357;
  wire tmp41358;
  wire tmp41359;
  wire tmp41360;
  wire tmp41361;
  wire tmp41362;
  wire tmp41363;
  wire tmp41364;
  wire tmp41365;
  wire tmp41366;
  wire tmp41367;
  wire tmp41368;
  wire tmp41369;
  wire tmp41370;
  wire tmp41371;
  wire tmp41372;
  wire tmp41373;
  wire tmp41374;
  wire tmp41375;
  wire tmp41376;
  wire tmp41377;
  wire tmp41378;
  wire tmp41379;
  wire tmp41380;
  wire tmp41381;
  wire tmp41382;
  wire tmp41383;
  wire tmp41384;
  wire tmp41385;
  wire tmp41386;
  wire tmp41387;
  wire tmp41388;
  wire tmp41389;
  wire tmp41390;
  wire tmp41391;
  wire tmp41392;
  wire tmp41393;
  wire tmp41394;
  wire tmp41395;
  wire tmp41396;
  wire tmp41397;
  wire tmp41398;
  wire tmp41399;
  wire tmp41400;
  wire tmp41401;
  wire tmp41402;
  wire tmp41403;
  wire tmp41404;
  wire tmp41405;
  wire tmp41406;
  wire tmp41407;
  wire tmp41408;
  wire tmp41409;
  wire tmp41410;
  wire tmp41411;
  wire tmp41412;
  wire tmp41413;
  wire tmp41414;
  wire tmp41415;
  wire tmp41416;
  wire tmp41417;
  wire tmp41418;
  wire tmp41419;
  wire tmp41420;
  wire tmp41421;
  wire tmp41422;
  wire tmp41423;
  wire tmp41424;
  wire tmp41425;
  wire tmp41426;
  wire tmp41427;
  wire tmp41428;
  wire tmp41429;
  wire tmp41430;
  wire tmp41431;
  wire tmp41432;
  wire tmp41433;
  wire tmp41434;
  wire tmp41435;
  wire tmp41436;
  wire tmp41437;
  wire tmp41438;
  wire tmp41439;
  wire tmp41440;
  wire tmp41441;
  wire tmp41442;
  wire tmp41443;
  wire tmp41444;
  wire tmp41445;
  wire tmp41446;
  wire tmp41447;
  wire tmp41448;
  wire tmp41449;
  wire tmp41450;
  wire tmp41451;
  wire tmp41452;
  wire tmp41453;
  wire tmp41454;
  wire tmp41455;
  wire tmp41456;
  wire tmp41457;
  wire tmp41458;
  wire tmp41459;
  wire tmp41460;
  wire tmp41461;
  wire tmp41462;
  wire tmp41463;
  wire tmp41464;
  wire tmp41465;
  wire tmp41466;
  wire tmp41467;
  wire tmp41468;
  wire tmp41469;
  wire tmp41470;
  wire tmp41471;
  wire tmp41472;
  wire tmp41473;
  wire tmp41474;
  wire tmp41475;
  wire tmp41476;
  wire tmp41477;
  wire tmp41478;
  wire tmp41479;
  wire tmp41480;
  wire tmp41481;
  wire tmp41482;
  wire tmp41483;
  wire tmp41484;
  wire tmp41485;
  wire tmp41486;
  wire tmp41487;
  wire tmp41488;
  wire tmp41489;
  wire tmp41490;
  wire tmp41491;
  wire tmp41492;
  wire tmp41493;
  wire tmp41494;
  wire tmp41495;
  wire tmp41496;
  wire tmp41497;
  wire tmp41498;
  wire tmp41499;
  wire tmp41500;
  wire tmp41501;
  wire tmp41502;
  wire tmp41503;
  wire tmp41504;
  wire tmp41505;
  wire tmp41506;
  wire tmp41507;
  wire tmp41508;
  wire tmp41509;
  wire tmp41510;
  wire tmp41511;
  wire tmp41512;
  wire tmp41513;
  wire tmp41514;
  wire tmp41515;
  wire tmp41516;
  wire tmp41517;
  wire tmp41518;
  wire tmp41519;
  wire tmp41520;
  wire tmp41521;
  wire tmp41522;
  wire tmp41523;
  wire tmp41524;
  wire tmp41525;
  wire tmp41526;
  wire tmp41527;
  wire tmp41528;
  wire tmp41529;
  wire tmp41530;
  wire tmp41531;
  wire tmp41532;
  wire tmp41533;
  wire tmp41534;
  wire tmp41535;
  wire tmp41536;
  wire tmp41537;
  wire tmp41538;
  wire tmp41539;
  wire tmp41540;
  wire tmp41541;
  wire tmp41542;
  wire tmp41543;
  wire tmp41544;
  wire tmp41545;
  wire tmp41546;
  wire tmp41547;
  wire tmp41548;
  wire tmp41549;
  wire tmp41550;
  wire tmp41551;
  wire tmp41552;
  wire tmp41553;
  wire tmp41554;
  wire tmp41555;
  wire tmp41556;
  wire tmp41557;
  wire tmp41558;
  wire tmp41559;
  wire tmp41560;
  wire tmp41561;
  wire tmp41562;
  wire tmp41563;
  wire tmp41564;
  wire tmp41565;
  wire tmp41566;
  wire tmp41567;
  wire tmp41568;
  wire tmp41569;
  wire tmp41570;
  wire tmp41571;
  wire tmp41572;
  wire tmp41573;
  wire tmp41574;
  wire tmp41575;
  wire tmp41576;
  wire tmp41577;
  wire tmp41578;
  wire tmp41579;
  wire tmp41580;
  wire tmp41581;
  wire tmp41582;
  wire tmp41583;
  wire tmp41584;
  wire tmp41585;
  wire tmp41586;
  wire tmp41587;
  wire tmp41588;
  wire tmp41589;
  wire tmp41590;
  wire tmp41591;
  wire tmp41592;
  wire tmp41593;
  wire tmp41594;
  wire tmp41595;
  wire tmp41596;
  wire tmp41597;
  wire tmp41598;
  wire tmp41599;
  wire tmp41600;
  wire tmp41601;
  wire tmp41602;
  wire tmp41603;
  wire tmp41604;
  wire tmp41605;
  wire tmp41606;
  wire tmp41607;
  wire tmp41608;
  wire tmp41609;
  wire tmp41610;
  wire tmp41611;
  wire tmp41612;
  wire tmp41613;
  wire tmp41614;
  wire tmp41615;
  wire tmp41616;
  wire tmp41617;
  wire tmp41618;
  wire tmp41619;
  wire tmp41620;
  wire tmp41621;
  wire tmp41622;
  wire tmp41623;
  wire tmp41624;
  wire tmp41625;
  wire tmp41626;
  wire tmp41627;
  wire tmp41628;
  wire tmp41629;
  wire tmp41630;
  wire tmp41631;
  wire tmp41632;
  wire tmp41633;
  wire tmp41634;
  wire tmp41635;
  wire tmp41636;
  wire tmp41637;
  wire tmp41638;
  wire tmp41639;
  wire tmp41640;
  wire tmp41641;
  wire tmp41642;
  wire tmp41643;
  wire tmp41644;
  wire tmp41645;
  wire tmp41646;
  wire tmp41647;
  wire tmp41648;
  wire tmp41649;
  wire tmp41650;
  wire tmp41651;
  wire tmp41652;
  wire tmp41653;
  wire tmp41654;
  wire tmp41655;
  wire tmp41656;
  wire tmp41657;
  wire tmp41658;
  wire tmp41659;
  wire tmp41660;
  wire tmp41661;
  wire tmp41662;
  wire tmp41663;
  wire tmp41664;
  wire tmp41665;
  wire tmp41666;
  wire tmp41667;
  wire tmp41668;
  wire tmp41669;
  wire tmp41670;
  wire tmp41671;
  wire tmp41672;
  wire tmp41673;
  wire tmp41674;
  wire tmp41675;
  wire tmp41676;
  wire tmp41677;
  wire tmp41678;
  wire tmp41679;
  wire tmp41680;
  wire tmp41681;
  wire tmp41682;
  wire tmp41683;
  wire tmp41684;
  wire tmp41685;
  wire tmp41686;
  wire tmp41687;
  wire tmp41688;
  wire tmp41689;
  wire tmp41690;
  wire tmp41691;
  wire tmp41692;
  wire tmp41693;
  wire tmp41694;
  wire tmp41695;
  wire tmp41696;
  wire tmp41697;
  wire tmp41698;
  wire tmp41699;
  wire tmp41700;
  wire tmp41701;
  wire tmp41702;
  wire tmp41703;
  wire tmp41704;
  wire tmp41705;
  wire tmp41706;
  wire tmp41707;
  wire tmp41708;
  wire tmp41709;
  wire tmp41710;
  wire tmp41711;
  wire tmp41712;
  wire tmp41713;
  wire tmp41714;
  wire tmp41715;
  wire tmp41716;
  wire tmp41717;
  wire tmp41718;
  wire tmp41719;
  wire tmp41720;
  wire tmp41721;
  wire tmp41722;
  wire tmp41723;
  wire tmp41724;
  wire tmp41725;
  wire tmp41726;
  wire tmp41727;
  wire tmp41728;
  wire tmp41729;
  wire tmp41730;
  wire tmp41731;
  wire tmp41732;
  wire tmp41733;
  wire tmp41734;
  wire tmp41735;
  wire tmp41736;
  wire tmp41737;
  wire tmp41738;
  wire tmp41739;
  wire tmp41740;
  wire tmp41741;
  wire tmp41742;
  wire tmp41743;
  wire tmp41744;
  wire tmp41745;
  wire tmp41746;
  wire tmp41747;
  wire tmp41748;
  wire tmp41749;
  wire tmp41750;
  wire tmp41751;
  wire tmp41752;
  wire tmp41753;
  wire tmp41754;
  wire tmp41755;
  wire tmp41756;
  wire tmp41757;
  wire tmp41758;
  wire tmp41759;
  wire tmp41760;
  wire tmp41761;
  wire tmp41762;
  wire tmp41763;
  wire tmp41764;
  wire tmp41765;
  wire tmp41766;
  wire tmp41767;
  wire tmp41768;
  wire tmp41769;
  wire tmp41770;
  wire tmp41771;
  wire tmp41772;
  wire tmp41773;
  wire tmp41774;
  wire tmp41775;
  wire tmp41776;
  wire tmp41777;
  wire tmp41778;
  wire tmp41779;
  wire tmp41780;
  wire tmp41781;
  wire tmp41782;
  wire tmp41783;
  wire tmp41784;
  wire tmp41785;
  wire tmp41786;
  wire tmp41787;
  wire tmp41788;
  wire tmp41789;
  wire tmp41790;
  wire tmp41791;
  wire tmp41792;
  wire tmp41793;
  wire tmp41794;
  wire tmp41795;
  wire tmp41796;
  wire tmp41797;
  wire tmp41798;
  wire tmp41799;
  wire tmp41800;
  wire tmp41801;
  wire tmp41802;
  wire tmp41803;
  wire tmp41804;
  wire tmp41805;
  wire tmp41806;
  wire tmp41807;
  wire tmp41808;
  wire tmp41809;
  wire tmp41810;
  wire tmp41811;
  wire tmp41812;
  wire tmp41813;
  wire tmp41814;
  wire tmp41815;
  wire tmp41816;
  wire tmp41817;
  wire tmp41818;
  wire tmp41819;
  wire tmp41820;
  wire tmp41821;
  wire tmp41822;
  wire tmp41823;
  wire tmp41824;
  wire tmp41825;
  wire tmp41826;
  wire tmp41827;
  wire tmp41828;
  wire tmp41829;
  wire tmp41830;
  wire tmp41831;
  wire tmp41832;
  wire tmp41833;
  wire tmp41834;
  wire tmp41835;
  wire tmp41836;
  wire tmp41837;
  wire tmp41838;
  wire tmp41839;
  wire tmp41840;
  wire tmp41841;
  wire tmp41842;
  wire tmp41843;
  wire tmp41844;
  wire tmp41845;
  wire tmp41846;
  wire tmp41847;
  wire tmp41848;
  wire tmp41849;
  wire tmp41850;
  wire tmp41851;
  wire tmp41852;
  wire tmp41853;
  wire tmp41854;
  wire tmp41855;
  wire tmp41856;
  wire tmp41857;
  wire tmp41858;
  wire tmp41859;
  wire tmp41860;
  wire tmp41861;
  wire tmp41862;
  wire tmp41863;
  wire tmp41864;
  wire tmp41865;
  wire tmp41866;
  wire tmp41867;
  wire tmp41868;
  wire tmp41869;
  wire tmp41870;
  wire tmp41871;
  wire tmp41872;
  wire tmp41873;
  wire tmp41874;
  wire tmp41875;
  wire tmp41876;
  wire tmp41877;
  wire tmp41878;
  wire tmp41879;
  wire tmp41880;
  wire tmp41881;
  wire tmp41882;
  wire tmp41883;
  wire tmp41884;
  wire tmp41885;
  wire tmp41886;
  wire tmp41887;
  wire tmp41888;
  wire tmp41889;
  wire tmp41890;
  wire tmp41891;
  wire tmp41892;
  wire tmp41893;
  wire tmp41894;
  wire tmp41895;
  wire tmp41896;
  wire tmp41897;
  wire tmp41898;
  wire tmp41899;
  wire tmp41900;
  wire tmp41901;
  wire tmp41902;
  wire tmp41903;
  wire tmp41904;
  wire tmp41905;
  wire tmp41906;
  wire tmp41907;
  wire tmp41908;
  wire tmp41909;
  wire tmp41910;
  wire tmp41911;
  wire tmp41912;
  wire tmp41913;
  wire tmp41914;
  wire tmp41915;
  wire tmp41916;
  wire tmp41917;
  wire tmp41918;
  wire tmp41919;
  wire tmp41920;
  wire tmp41921;
  wire tmp41922;
  wire tmp41923;
  wire tmp41924;
  wire tmp41925;
  wire tmp41926;
  wire tmp41927;
  wire tmp41928;
  wire tmp41929;
  wire tmp41930;
  wire tmp41931;
  wire tmp41932;
  wire tmp41933;
  wire tmp41934;
  wire tmp41935;
  wire tmp41936;
  wire tmp41937;
  wire tmp41938;
  wire tmp41939;
  wire tmp41940;
  wire tmp41941;
  wire tmp41942;
  wire tmp41943;
  wire tmp41944;
  wire tmp41945;
  wire tmp41946;
  wire tmp41947;
  wire tmp41948;
  wire tmp41949;
  wire tmp41950;
  wire tmp41951;
  wire tmp41952;
  wire tmp41953;
  wire tmp41954;
  wire tmp41955;
  wire tmp41956;
  wire tmp41957;
  wire tmp41958;
  wire tmp41959;
  wire tmp41960;
  wire tmp41961;
  wire tmp41962;
  wire tmp41963;
  wire tmp41964;
  wire tmp41965;
  wire tmp41966;
  wire tmp41967;
  wire tmp41968;
  wire tmp41969;
  wire tmp41970;
  wire tmp41971;
  wire tmp41972;
  wire tmp41973;
  wire tmp41974;
  wire tmp41975;
  wire tmp41976;
  wire tmp41977;
  wire tmp41978;
  wire tmp41979;
  wire tmp41980;
  wire tmp41981;
  wire tmp41982;
  wire tmp41983;
  wire tmp41984;
  wire tmp41985;
  wire tmp41986;
  wire tmp41987;
  wire tmp41988;
  wire tmp41989;
  wire tmp41990;
  wire tmp41991;
  wire tmp41992;
  wire tmp41993;
  wire tmp41994;
  wire tmp41995;
  wire tmp41996;
  wire tmp41997;
  wire tmp41998;
  wire tmp41999;
  wire tmp42000;
  wire tmp42001;
  wire tmp42002;
  wire tmp42003;
  wire tmp42004;
  wire tmp42005;
  wire tmp42006;
  wire tmp42007;
  wire tmp42008;
  wire tmp42009;
  wire tmp42010;
  wire tmp42011;
  wire tmp42012;
  wire tmp42013;
  wire tmp42014;
  wire tmp42015;
  wire tmp42016;
  wire tmp42017;
  wire tmp42018;
  wire tmp42019;
  wire tmp42020;
  wire tmp42021;
  wire tmp42022;
  wire tmp42023;
  wire tmp42024;
  wire tmp42025;
  wire tmp42026;
  wire tmp42027;
  wire tmp42028;
  wire tmp42029;
  wire tmp42030;
  wire tmp42031;
  wire tmp42032;
  wire tmp42033;
  wire tmp42034;
  wire tmp42035;
  wire tmp42036;
  wire tmp42037;
  wire tmp42038;
  wire tmp42039;
  wire tmp42040;
  wire tmp42041;
  wire tmp42042;
  wire tmp42043;
  wire tmp42044;
  wire tmp42045;
  wire tmp42046;
  wire tmp42047;
  wire tmp42048;
  wire tmp42049;
  wire tmp42050;
  wire tmp42051;
  wire tmp42052;
  wire tmp42053;
  wire tmp42054;
  wire tmp42055;
  wire tmp42056;
  wire tmp42057;
  wire tmp42058;
  wire tmp42059;
  wire tmp42060;
  wire tmp42061;
  wire tmp42062;
  wire tmp42063;
  wire tmp42064;
  wire tmp42065;
  wire tmp42066;
  wire tmp42067;
  wire tmp42068;
  wire tmp42069;
  wire tmp42070;
  wire tmp42071;
  wire tmp42072;
  wire tmp42073;
  wire tmp42074;
  wire tmp42075;
  wire tmp42076;
  wire tmp42077;
  wire tmp42078;
  wire tmp42079;
  wire tmp42080;
  wire tmp42081;
  wire tmp42082;
  wire tmp42083;
  wire tmp42084;
  wire tmp42085;
  wire tmp42086;
  wire tmp42087;
  wire tmp42088;
  wire tmp42089;
  wire tmp42090;
  wire tmp42091;
  wire tmp42092;
  wire tmp42093;
  wire tmp42094;
  wire tmp42095;
  wire tmp42096;
  wire tmp42097;
  wire tmp42098;
  wire tmp42099;
  wire tmp42100;
  wire tmp42101;
  wire tmp42102;
  wire tmp42103;
  wire tmp42104;
  wire tmp42105;
  wire tmp42106;
  wire tmp42107;
  wire tmp42108;
  wire tmp42109;
  wire tmp42110;
  wire tmp42111;
  wire tmp42112;
  wire tmp42113;
  wire tmp42114;
  wire tmp42115;
  wire tmp42116;
  wire tmp42117;
  wire tmp42118;
  wire tmp42119;
  wire tmp42120;
  wire tmp42121;
  wire tmp42122;
  wire tmp42123;
  wire tmp42124;
  wire tmp42125;
  wire tmp42126;
  wire tmp42127;
  wire tmp42128;
  wire tmp42129;
  wire tmp42130;
  wire tmp42131;
  wire tmp42132;
  wire tmp42133;
  wire tmp42134;
  wire tmp42135;
  wire tmp42136;
  wire tmp42137;
  wire tmp42138;
  wire tmp42139;
  wire tmp42140;
  wire tmp42141;
  wire tmp42142;
  wire tmp42143;
  wire tmp42144;
  wire tmp42145;
  wire tmp42146;
  wire tmp42147;
  wire tmp42148;
  wire tmp42149;
  wire tmp42150;
  wire tmp42151;
  wire tmp42152;
  wire tmp42153;
  wire tmp42154;
  wire tmp42155;
  wire tmp42156;
  wire tmp42157;
  wire tmp42158;
  wire tmp42159;
  wire tmp42160;
  wire tmp42161;
  wire tmp42162;
  wire tmp42163;
  wire tmp42164;
  wire tmp42165;
  wire tmp42166;
  wire tmp42167;
  wire tmp42168;
  wire tmp42169;
  wire tmp42170;
  wire tmp42171;
  wire tmp42172;
  wire tmp42173;
  wire tmp42174;
  wire tmp42175;
  wire tmp42176;
  wire tmp42177;
  wire tmp42178;
  wire tmp42179;
  wire tmp42180;
  wire tmp42181;
  wire tmp42182;
  wire tmp42183;
  wire tmp42184;
  wire tmp42185;
  wire tmp42186;
  wire tmp42187;
  wire tmp42188;
  wire tmp42189;
  wire tmp42190;
  wire tmp42191;
  wire tmp42192;
  wire tmp42193;
  wire tmp42194;
  wire tmp42195;
  wire tmp42196;
  wire tmp42197;
  wire tmp42198;
  wire tmp42199;
  wire tmp42200;
  wire tmp42201;
  wire tmp42202;
  wire tmp42203;
  wire tmp42204;
  wire tmp42205;
  wire tmp42206;
  wire tmp42207;
  wire tmp42208;
  wire tmp42209;
  wire tmp42210;
  wire tmp42211;
  wire tmp42212;
  wire tmp42213;
  wire tmp42214;
  wire tmp42215;
  wire tmp42216;
  wire tmp42217;
  wire tmp42218;
  wire tmp42219;
  wire tmp42220;
  wire tmp42221;
  wire tmp42222;
  wire tmp42223;
  wire tmp42224;
  wire tmp42225;
  wire tmp42226;
  wire tmp42227;
  wire tmp42228;
  wire tmp42229;
  wire tmp42230;
  wire tmp42231;
  wire tmp42232;
  wire tmp42233;
  wire tmp42234;
  wire tmp42235;
  wire tmp42236;
  wire tmp42237;
  wire tmp42238;
  wire tmp42239;
  wire tmp42240;
  wire tmp42241;
  wire tmp42242;
  wire tmp42243;
  wire tmp42244;
  wire tmp42245;
  wire tmp42246;
  wire tmp42247;
  wire tmp42248;
  wire tmp42249;
  wire tmp42250;
  wire tmp42251;
  wire tmp42252;
  wire tmp42253;
  wire tmp42254;
  wire tmp42255;
  wire tmp42256;
  wire tmp42257;
  wire tmp42258;
  wire tmp42259;
  wire tmp42260;
  wire tmp42261;
  wire tmp42262;
  wire tmp42263;
  wire tmp42264;
  wire tmp42265;
  wire tmp42266;
  wire tmp42267;
  wire tmp42268;
  wire tmp42269;
  wire tmp42270;
  wire tmp42271;
  wire tmp42272;
  wire tmp42273;
  wire tmp42274;
  wire tmp42275;
  wire tmp42276;
  wire tmp42277;
  wire tmp42278;
  wire tmp42279;
  wire tmp42280;
  wire tmp42281;
  wire tmp42282;
  wire tmp42283;
  wire tmp42284;
  wire tmp42285;
  wire tmp42286;
  wire tmp42287;
  wire tmp42288;
  wire tmp42289;
  wire tmp42290;
  wire tmp42291;
  wire tmp42292;
  wire tmp42293;
  wire tmp42294;
  wire tmp42295;
  wire tmp42296;
  wire tmp42297;
  wire tmp42298;
  wire tmp42299;
  wire tmp42300;
  wire tmp42301;
  wire tmp42302;
  wire tmp42303;
  wire tmp42304;
  wire tmp42305;
  wire tmp42306;
  wire tmp42307;
  wire tmp42308;
  wire tmp42309;
  wire tmp42310;
  wire tmp42311;
  wire tmp42312;
  wire tmp42313;
  wire tmp42314;
  wire tmp42315;
  wire tmp42316;
  wire tmp42317;
  wire tmp42318;
  wire tmp42319;
  wire tmp42320;
  wire tmp42321;
  wire tmp42322;
  wire tmp42323;
  wire tmp42324;
  wire tmp42325;
  wire tmp42326;
  wire tmp42327;
  wire tmp42328;
  wire tmp42329;
  wire tmp42330;
  wire tmp42331;
  wire tmp42332;
  wire tmp42333;
  wire tmp42334;
  wire tmp42335;
  wire tmp42336;
  wire tmp42337;
  wire tmp42338;
  wire tmp42339;
  wire tmp42340;
  wire tmp42341;
  wire tmp42342;
  wire tmp42343;
  wire tmp42344;
  wire tmp42345;
  wire tmp42346;
  wire tmp42347;
  wire tmp42348;
  wire tmp42349;
  wire tmp42350;
  wire tmp42351;
  wire tmp42352;
  wire tmp42353;
  wire tmp42354;
  wire tmp42355;
  wire tmp42356;
  wire tmp42357;
  wire tmp42358;
  wire tmp42359;
  wire tmp42360;
  wire tmp42361;
  wire tmp42362;
  wire tmp42363;
  wire tmp42364;
  wire tmp42365;
  wire tmp42366;
  wire tmp42367;
  wire tmp42368;
  wire tmp42369;
  wire tmp42370;
  wire tmp42371;
  wire tmp42372;
  wire tmp42373;
  wire tmp42374;
  wire tmp42375;
  wire tmp42376;
  wire tmp42377;
  wire tmp42378;
  wire tmp42379;
  wire tmp42380;
  wire tmp42381;
  wire tmp42382;
  wire tmp42383;
  wire tmp42384;
  wire tmp42385;
  wire tmp42386;
  wire tmp42387;
  wire tmp42388;
  wire tmp42389;
  wire tmp42390;
  wire tmp42391;
  wire tmp42392;
  wire tmp42393;
  wire tmp42394;
  wire tmp42395;
  wire tmp42396;
  wire tmp42397;
  wire tmp42398;
  wire tmp42399;
  wire tmp42400;
  wire tmp42401;
  wire tmp42402;
  wire tmp42403;
  wire tmp42404;
  wire tmp42405;
  wire tmp42406;
  wire tmp42407;
  wire tmp42408;
  wire tmp42409;
  wire tmp42410;
  wire tmp42411;
  wire tmp42412;
  wire tmp42413;
  wire tmp42414;
  wire tmp42415;
  wire tmp42416;
  wire tmp42417;
  wire tmp42418;
  wire tmp42419;
  wire tmp42420;
  wire tmp42421;
  wire tmp42422;
  wire tmp42423;
  wire tmp42424;
  wire tmp42425;
  wire tmp42426;
  wire tmp42427;
  wire tmp42428;
  wire tmp42429;
  wire tmp42430;
  wire tmp42431;
  wire tmp42432;
  wire tmp42433;
  wire tmp42434;
  wire tmp42435;
  wire tmp42436;
  wire tmp42437;
  wire tmp42438;
  wire tmp42439;
  wire tmp42440;
  wire tmp42441;
  wire tmp42442;
  wire tmp42443;
  wire tmp42444;
  wire tmp42445;
  wire tmp42446;
  wire tmp42447;
  wire tmp42448;
  wire tmp42449;
  wire tmp42450;
  wire tmp42451;
  wire tmp42452;
  wire tmp42453;
  wire tmp42454;
  wire tmp42455;
  wire tmp42456;
  wire tmp42457;
  wire tmp42458;
  wire tmp42459;
  wire tmp42460;
  wire tmp42461;
  wire tmp42462;
  wire tmp42463;
  wire tmp42464;
  wire tmp42465;
  wire tmp42466;
  wire tmp42467;
  wire tmp42468;
  wire tmp42469;
  wire tmp42470;
  wire tmp42471;
  wire tmp42472;
  wire tmp42473;
  wire tmp42474;
  wire tmp42475;
  wire tmp42476;
  wire tmp42477;
  wire tmp42478;
  wire tmp42479;
  wire tmp42480;
  wire tmp42481;
  wire tmp42482;
  wire tmp42483;
  wire tmp42484;
  wire tmp42485;
  wire tmp42486;
  wire tmp42487;
  wire tmp42488;
  wire tmp42489;
  wire tmp42490;
  wire tmp42491;
  wire tmp42492;
  wire tmp42493;
  wire tmp42494;
  wire tmp42495;
  wire tmp42496;
  wire tmp42497;
  wire tmp42498;
  wire tmp42499;
  wire tmp42500;
  wire tmp42501;
  wire tmp42502;
  wire tmp42503;
  wire tmp42504;
  wire tmp42505;
  wire tmp42506;
  wire tmp42507;
  wire tmp42508;
  wire tmp42509;
  wire tmp42510;
  wire tmp42511;
  wire tmp42512;
  wire tmp42513;
  wire tmp42514;
  wire tmp42515;
  wire tmp42516;
  wire tmp42517;
  wire tmp42518;
  wire tmp42519;
  wire tmp42520;
  wire tmp42521;
  wire tmp42522;
  wire tmp42523;
  wire tmp42524;
  wire tmp42525;
  wire tmp42526;
  wire tmp42527;
  wire tmp42528;
  wire tmp42529;
  wire tmp42530;
  wire tmp42531;
  wire tmp42532;
  wire tmp42533;
  wire tmp42534;
  wire tmp42535;
  wire tmp42536;
  wire tmp42537;
  wire tmp42538;
  wire tmp42539;
  wire tmp42540;
  wire tmp42541;
  wire tmp42542;
  wire tmp42543;
  wire tmp42544;
  wire tmp42545;
  wire tmp42546;
  wire tmp42547;
  wire tmp42548;
  wire tmp42549;
  wire tmp42550;
  wire tmp42551;
  wire tmp42552;
  wire tmp42553;
  wire tmp42554;
  wire tmp42555;
  wire tmp42556;
  wire tmp42557;
  wire tmp42558;
  wire tmp42559;
  wire tmp42560;
  wire tmp42561;
  wire tmp42562;
  wire tmp42563;
  wire tmp42564;
  wire tmp42565;
  wire tmp42566;
  wire tmp42567;
  wire tmp42568;
  wire tmp42569;
  wire tmp42570;
  wire tmp42571;
  wire tmp42572;
  wire tmp42573;
  wire tmp42574;
  wire tmp42575;
  wire tmp42576;
  wire tmp42577;
  wire tmp42578;
  wire tmp42579;
  wire tmp42580;
  wire tmp42581;
  wire tmp42582;
  wire tmp42583;
  wire tmp42584;
  wire tmp42585;
  wire tmp42586;
  wire tmp42587;
  wire tmp42588;
  wire tmp42589;
  wire tmp42590;
  wire tmp42591;
  wire tmp42592;
  wire tmp42593;
  wire tmp42594;
  wire tmp42595;
  wire tmp42596;
  wire tmp42597;
  wire tmp42598;
  wire tmp42599;
  wire tmp42600;
  wire tmp42601;
  wire tmp42602;
  wire tmp42603;
  wire tmp42604;
  wire tmp42605;
  wire tmp42606;
  wire tmp42607;
  wire tmp42608;
  wire tmp42609;
  wire tmp42610;
  wire tmp42611;
  wire tmp42612;
  wire tmp42613;
  wire tmp42614;
  wire tmp42615;
  wire tmp42616;
  wire tmp42617;
  wire tmp42618;
  wire tmp42619;
  wire tmp42620;
  wire tmp42621;
  wire tmp42622;
  wire tmp42623;
  wire tmp42624;
  wire tmp42625;
  wire tmp42626;
  wire tmp42627;
  wire tmp42628;
  wire tmp42629;
  wire tmp42630;
  wire tmp42631;
  wire tmp42632;
  wire tmp42633;
  wire tmp42634;
  wire tmp42635;
  wire tmp42636;
  wire tmp42637;
  wire tmp42638;
  wire tmp42639;
  wire tmp42640;
  wire tmp42641;
  wire tmp42642;
  wire tmp42643;
  wire tmp42644;
  wire tmp42645;
  wire tmp42646;
  wire tmp42647;
  wire tmp42648;
  wire tmp42649;
  wire tmp42650;
  wire tmp42651;
  wire tmp42652;
  wire tmp42653;
  wire tmp42654;
  wire tmp42655;
  wire tmp42656;
  wire tmp42657;
  wire tmp42658;
  wire tmp42659;
  wire tmp42660;
  wire tmp42661;
  wire tmp42662;
  wire tmp42663;
  wire tmp42664;
  wire tmp42665;
  wire tmp42666;
  wire tmp42667;
  wire tmp42668;
  wire tmp42669;
  wire tmp42670;
  wire tmp42671;
  wire tmp42672;
  wire tmp42673;
  wire tmp42674;
  wire tmp42675;
  wire tmp42676;
  wire tmp42677;
  wire tmp42678;
  wire tmp42679;
  wire tmp42680;
  wire tmp42681;
  wire tmp42682;
  wire tmp42683;
  wire tmp42684;
  wire tmp42685;
  wire tmp42686;
  wire tmp42687;
  wire tmp42688;
  wire tmp42689;
  wire tmp42690;
  wire tmp42691;
  wire tmp42692;
  wire tmp42693;
  wire tmp42694;
  wire tmp42695;
  wire tmp42696;
  wire tmp42697;
  wire tmp42698;
  wire tmp42699;
  wire tmp42700;
  wire tmp42701;
  wire tmp42702;
  wire tmp42703;
  wire tmp42704;
  wire tmp42705;
  wire tmp42706;
  wire tmp42707;
  wire tmp42708;
  wire tmp42709;
  wire tmp42710;
  wire tmp42711;
  wire tmp42712;
  wire tmp42713;
  wire tmp42714;
  wire tmp42715;
  wire tmp42716;
  wire tmp42717;
  wire tmp42718;
  wire tmp42719;
  wire tmp42720;
  wire tmp42721;
  wire tmp42722;
  wire tmp42723;
  wire tmp42724;
  wire tmp42725;
  wire tmp42726;
  wire tmp42727;
  wire tmp42728;
  wire tmp42729;
  wire tmp42730;
  wire tmp42731;
  wire tmp42732;
  wire tmp42733;
  wire tmp42734;
  wire tmp42735;
  wire tmp42736;
  wire tmp42737;
  wire tmp42738;
  wire tmp42739;
  wire tmp42740;
  wire tmp42741;
  wire tmp42742;
  wire tmp42743;
  wire tmp42744;
  wire tmp42745;
  wire tmp42746;
  wire tmp42747;
  wire tmp42748;
  wire tmp42749;
  wire tmp42750;
  wire tmp42751;
  wire tmp42752;
  wire tmp42753;
  wire tmp42754;
  wire tmp42755;
  wire tmp42756;
  wire tmp42757;
  wire tmp42758;
  wire tmp42759;
  wire tmp42760;
  wire tmp42761;
  wire tmp42762;
  wire tmp42763;
  wire tmp42764;
  wire tmp42765;
  wire tmp42766;
  wire tmp42767;
  wire tmp42768;
  wire tmp42769;
  wire tmp42770;
  wire tmp42771;
  wire tmp42772;
  wire tmp42773;
  wire tmp42774;
  wire tmp42775;
  wire tmp42776;
  wire tmp42777;
  wire tmp42778;
  wire tmp42779;
  wire tmp42780;
  wire tmp42781;
  wire tmp42782;
  wire tmp42783;
  wire tmp42784;
  wire tmp42785;
  wire tmp42786;
  wire tmp42787;
  wire tmp42788;
  wire tmp42789;
  wire tmp42790;
  wire tmp42791;
  wire tmp42792;
  wire tmp42793;
  wire tmp42794;
  wire tmp42795;
  wire tmp42796;
  wire tmp42797;
  wire tmp42798;
  wire tmp42799;
  wire tmp42800;
  wire tmp42801;
  wire tmp42802;
  wire tmp42803;
  wire tmp42804;
  wire tmp42805;
  wire tmp42806;
  wire tmp42807;
  wire tmp42808;
  wire tmp42809;
  wire tmp42810;
  wire tmp42811;
  wire tmp42812;
  wire tmp42813;
  wire tmp42814;
  wire tmp42815;
  wire tmp42816;
  wire tmp42817;
  wire tmp42818;
  wire tmp42819;
  wire tmp42820;
  wire tmp42821;
  wire tmp42822;
  wire tmp42823;
  wire tmp42824;
  wire tmp42825;
  wire tmp42826;
  wire tmp42827;
  wire tmp42828;
  wire tmp42829;
  wire tmp42830;
  wire tmp42831;
  wire tmp42832;
  wire tmp42833;
  wire tmp42834;
  wire tmp42835;
  wire tmp42836;
  wire tmp42837;
  wire tmp42838;
  wire tmp42839;
  wire tmp42840;
  wire tmp42841;
  wire tmp42842;
  wire tmp42843;
  wire tmp42844;
  wire tmp42845;
  wire tmp42846;
  wire tmp42847;
  wire tmp42848;
  wire tmp42849;
  wire tmp42850;
  wire tmp42851;
  wire tmp42852;
  wire tmp42853;
  wire tmp42854;
  wire tmp42855;
  wire tmp42856;
  wire tmp42857;
  wire tmp42858;
  wire tmp42859;
  wire tmp42860;
  wire tmp42861;
  wire tmp42862;
  wire tmp42863;
  wire tmp42864;
  wire tmp42865;
  wire tmp42866;
  wire tmp42867;
  wire tmp42868;
  wire tmp42869;
  wire tmp42870;
  wire tmp42871;
  wire tmp42872;
  wire tmp42873;
  wire tmp42874;
  wire tmp42875;
  wire tmp42876;
  wire tmp42877;
  wire tmp42878;
  wire tmp42879;
  wire tmp42880;
  wire tmp42881;
  wire tmp42882;
  wire tmp42883;
  wire tmp42884;
  wire tmp42885;
  wire tmp42886;
  wire tmp42887;
  wire tmp42888;
  wire tmp42889;
  wire tmp42890;
  wire tmp42891;
  wire tmp42892;
  wire tmp42893;
  wire tmp42894;
  wire tmp42895;
  wire tmp42896;
  wire tmp42897;
  wire tmp42898;
  wire tmp42899;
  wire tmp42900;
  wire tmp42901;
  wire tmp42902;
  wire tmp42903;
  wire tmp42904;
  wire tmp42905;
  wire tmp42906;
  wire tmp42907;
  wire tmp42908;
  wire tmp42909;
  wire tmp42910;
  wire tmp42911;
  wire tmp42912;
  wire tmp42913;
  wire tmp42914;
  wire tmp42915;
  wire tmp42916;
  wire tmp42917;
  wire tmp42918;
  wire tmp42919;
  wire tmp42920;
  wire tmp42921;
  wire tmp42922;
  wire tmp42923;
  wire tmp42924;
  wire tmp42925;
  wire tmp42926;
  wire tmp42927;
  wire tmp42928;
  wire tmp42929;
  wire tmp42930;
  wire tmp42931;
  wire tmp42932;
  wire tmp42933;
  wire tmp42934;
  wire tmp42935;
  wire tmp42936;
  wire tmp42937;
  wire tmp42938;
  wire tmp42939;
  wire tmp42940;
  wire tmp42941;
  wire tmp42942;
  wire tmp42943;
  wire tmp42944;
  wire tmp42945;
  wire tmp42946;
  wire tmp42947;
  wire tmp42948;
  wire tmp42949;
  wire tmp42950;
  wire tmp42951;
  wire tmp42952;
  wire tmp42953;
  wire tmp42954;
  wire tmp42955;
  wire tmp42956;
  wire tmp42957;
  wire tmp42958;
  wire tmp42959;
  wire tmp42960;
  wire tmp42961;
  wire tmp42962;
  wire tmp42963;
  wire tmp42964;
  wire tmp42965;
  wire tmp42966;
  wire tmp42967;
  wire tmp42968;
  wire tmp42969;
  wire tmp42970;
  wire tmp42971;
  wire tmp42972;
  wire tmp42973;
  wire tmp42974;
  wire tmp42975;
  wire tmp42976;
  wire tmp42977;
  wire tmp42978;
  wire tmp42979;
  wire tmp42980;
  wire tmp42981;
  wire tmp42982;
  wire tmp42983;
  wire tmp42984;
  wire tmp42985;
  wire tmp42986;
  wire tmp42987;
  wire tmp42988;
  wire tmp42989;
  wire tmp42990;
  wire tmp42991;
  wire tmp42992;
  wire tmp42993;
  wire tmp42994;
  wire tmp42995;
  wire tmp42996;
  wire tmp42997;
  wire tmp42998;
  wire tmp42999;
  wire tmp43000;
  wire tmp43001;
  wire tmp43002;
  wire tmp43003;
  wire tmp43004;
  wire tmp43005;
  wire tmp43006;
  wire tmp43007;
  wire tmp43008;
  wire tmp43009;
  wire tmp43010;
  wire tmp43011;
  wire tmp43012;
  wire tmp43013;
  wire tmp43014;
  wire tmp43015;
  wire tmp43016;
  wire tmp43017;
  wire tmp43018;
  wire tmp43019;
  wire tmp43020;
  wire tmp43021;
  wire tmp43022;
  wire tmp43023;
  wire tmp43024;
  wire tmp43025;
  wire tmp43026;
  wire tmp43027;
  wire tmp43028;
  wire tmp43029;
  wire tmp43030;
  wire tmp43031;
  wire tmp43032;
  wire tmp43033;
  wire tmp43034;
  wire tmp43035;
  wire tmp43036;
  wire tmp43037;
  wire tmp43038;
  wire tmp43039;
  wire tmp43040;
  wire tmp43041;
  wire tmp43042;
  wire tmp43043;
  wire tmp43044;
  wire tmp43045;
  wire tmp43046;
  wire tmp43047;
  wire tmp43048;
  wire tmp43049;
  wire tmp43050;
  wire tmp43051;
  wire tmp43052;
  wire tmp43053;
  wire tmp43054;
  wire tmp43055;
  wire tmp43056;
  wire tmp43057;
  wire tmp43058;
  wire tmp43059;
  wire tmp43060;
  wire tmp43061;
  wire tmp43062;
  wire tmp43063;
  wire tmp43064;
  wire tmp43065;
  wire tmp43066;
  wire tmp43067;
  wire tmp43068;
  wire tmp43069;
  wire tmp43070;
  wire tmp43071;
  wire tmp43072;
  wire tmp43073;
  wire tmp43074;
  wire tmp43075;
  wire tmp43076;
  wire tmp43077;
  wire tmp43078;
  wire tmp43079;
  wire tmp43080;
  wire tmp43081;
  wire tmp43082;
  wire tmp43083;
  wire tmp43084;
  wire tmp43085;
  wire tmp43086;
  wire tmp43087;
  wire tmp43088;
  wire tmp43089;
  wire tmp43090;
  wire tmp43091;
  wire tmp43092;
  wire tmp43093;
  wire tmp43094;
  wire tmp43095;
  wire tmp43096;
  wire tmp43097;
  wire tmp43098;
  wire tmp43099;
  wire tmp43100;
  wire tmp43101;
  wire tmp43102;
  wire tmp43103;
  wire tmp43104;
  wire tmp43105;
  wire tmp43106;
  wire tmp43107;
  wire tmp43108;
  wire tmp43109;
  wire tmp43110;
  wire tmp43111;
  wire tmp43112;
  wire tmp43113;
  wire tmp43114;
  wire tmp43115;
  wire tmp43116;
  wire tmp43117;
  wire tmp43118;
  wire tmp43119;
  wire tmp43120;
  wire tmp43121;
  wire tmp43122;
  wire tmp43123;
  wire tmp43124;
  wire tmp43125;
  wire tmp43126;
  wire tmp43127;
  wire tmp43128;
  wire tmp43129;
  wire tmp43130;
  wire tmp43131;
  wire tmp43132;
  wire tmp43133;
  wire tmp43134;
  wire tmp43135;
  wire tmp43136;
  wire tmp43137;
  wire tmp43138;
  wire tmp43139;
  wire tmp43140;
  wire tmp43141;
  wire tmp43142;
  wire tmp43143;
  wire tmp43144;
  wire tmp43145;
  wire tmp43146;
  wire tmp43147;
  wire tmp43148;
  wire tmp43149;
  wire tmp43150;
  wire tmp43151;
  wire tmp43152;
  wire tmp43153;
  wire tmp43154;
  wire tmp43155;
  wire tmp43156;
  wire tmp43157;
  wire tmp43158;
  wire tmp43159;
  wire tmp43160;
  wire tmp43161;
  wire tmp43162;
  wire tmp43163;
  wire tmp43164;
  wire tmp43165;
  wire tmp43166;
  wire tmp43167;
  wire tmp43168;
  wire tmp43169;
  wire tmp43170;
  wire tmp43171;
  wire tmp43172;
  wire tmp43173;
  wire tmp43174;
  wire tmp43175;
  wire tmp43176;
  wire tmp43177;
  wire tmp43178;
  wire tmp43179;
  wire tmp43180;
  wire tmp43181;
  wire tmp43182;
  wire tmp43183;
  wire tmp43184;
  wire tmp43185;
  wire tmp43186;
  wire tmp43187;
  wire tmp43188;
  wire tmp43189;
  wire tmp43190;
  wire tmp43191;
  wire tmp43192;
  wire tmp43193;
  wire tmp43194;
  wire tmp43195;
  wire tmp43196;
  wire tmp43197;
  wire tmp43198;
  wire tmp43199;
  wire tmp43200;
  wire tmp43201;
  wire tmp43202;
  wire tmp43203;
  wire tmp43204;
  wire tmp43205;
  wire tmp43206;
  wire tmp43207;
  wire tmp43208;
  wire tmp43209;
  wire tmp43210;
  wire tmp43211;
  wire tmp43212;
  wire tmp43213;
  wire tmp43214;
  wire tmp43215;
  wire tmp43216;
  wire tmp43217;
  wire tmp43218;
  wire tmp43219;
  wire tmp43220;
  wire tmp43221;
  wire tmp43222;
  wire tmp43223;
  wire tmp43224;
  wire tmp43225;
  wire tmp43226;
  wire tmp43227;
  wire tmp43228;
  wire tmp43229;
  wire tmp43230;
  wire tmp43231;
  wire tmp43232;
  wire tmp43233;
  wire tmp43234;
  wire tmp43235;
  wire tmp43236;
  wire tmp43237;
  wire tmp43238;
  wire tmp43239;
  wire tmp43240;
  wire tmp43241;
  wire tmp43242;
  wire tmp43243;
  wire tmp43244;
  wire tmp43245;
  wire tmp43246;
  wire tmp43247;
  wire tmp43248;
  wire tmp43249;
  wire tmp43250;
  wire tmp43251;
  wire tmp43252;
  wire tmp43253;
  wire tmp43254;
  wire tmp43255;
  wire tmp43256;
  wire tmp43257;
  wire tmp43258;
  wire tmp43259;
  wire tmp43260;
  wire tmp43261;
  wire tmp43262;
  wire tmp43263;
  wire tmp43264;
  wire tmp43265;
  wire tmp43266;
  wire tmp43267;
  wire tmp43268;
  wire tmp43269;
  wire tmp43270;
  wire tmp43271;
  wire tmp43272;
  wire tmp43273;
  wire tmp43274;
  wire tmp43275;
  wire tmp43276;
  wire tmp43277;
  wire tmp43278;
  wire tmp43279;
  wire tmp43280;
  wire tmp43281;
  wire tmp43282;
  wire tmp43283;
  wire tmp43284;
  wire tmp43285;
  wire tmp43286;
  wire tmp43287;
  wire tmp43288;
  wire tmp43289;
  wire tmp43290;
  wire tmp43291;
  wire tmp43292;
  wire tmp43293;
  wire tmp43294;
  wire tmp43295;
  wire tmp43296;
  wire tmp43297;
  wire tmp43298;
  wire tmp43299;
  wire tmp43300;
  wire tmp43301;
  wire tmp43302;
  wire tmp43303;
  wire tmp43304;
  wire tmp43305;
  wire tmp43306;
  wire tmp43307;
  wire tmp43308;
  wire tmp43309;
  wire tmp43310;
  wire tmp43311;
  wire tmp43312;
  wire tmp43313;
  wire tmp43314;
  wire tmp43315;
  wire tmp43316;
  wire tmp43317;
  wire tmp43318;
  wire tmp43319;
  wire tmp43320;
  wire tmp43321;
  wire tmp43322;
  wire tmp43323;
  wire tmp43324;
  wire tmp43325;
  wire tmp43326;
  wire tmp43327;
  wire tmp43328;
  wire tmp43329;
  wire tmp43330;
  wire tmp43331;
  wire tmp43332;
  wire tmp43333;
  wire tmp43334;
  wire tmp43335;
  wire tmp43336;
  wire tmp43337;
  wire tmp43338;
  wire tmp43339;
  wire tmp43340;
  wire tmp43341;
  wire tmp43342;
  wire tmp43343;
  wire tmp43344;
  wire tmp43345;
  wire tmp43346;
  wire tmp43347;
  wire tmp43348;
  wire tmp43349;
  wire tmp43350;
  wire tmp43351;
  wire tmp43352;
  wire tmp43353;
  wire tmp43354;
  wire tmp43355;
  wire tmp43356;
  wire tmp43357;
  wire tmp43358;
  wire tmp43359;
  wire tmp43360;
  wire tmp43361;
  wire tmp43362;
  wire tmp43363;
  wire tmp43364;
  wire tmp43365;
  wire tmp43366;
  wire tmp43367;
  wire tmp43368;
  wire tmp43369;
  wire tmp43370;
  wire tmp43371;
  wire tmp43372;
  wire tmp43373;
  wire tmp43374;
  wire tmp43375;
  wire tmp43376;
  wire tmp43377;
  wire tmp43378;
  wire tmp43379;
  wire tmp43380;
  wire tmp43381;
  wire tmp43382;
  wire tmp43383;
  wire tmp43384;
  wire tmp43385;
  wire tmp43386;
  wire tmp43387;
  wire tmp43388;
  wire tmp43389;
  wire tmp43390;
  wire tmp43391;
  wire tmp43392;
  wire tmp43393;
  wire tmp43394;
  wire tmp43395;
  wire tmp43396;
  wire tmp43397;
  wire tmp43398;
  wire tmp43399;
  wire tmp43400;
  wire tmp43401;
  wire tmp43402;
  wire tmp43403;
  wire tmp43404;
  wire tmp43405;
  wire tmp43406;
  wire tmp43407;
  wire tmp43408;
  wire tmp43409;
  wire tmp43410;
  wire tmp43411;
  wire tmp43412;
  wire tmp43413;
  wire tmp43414;
  wire tmp43415;
  wire tmp43416;
  wire tmp43417;
  wire tmp43418;
  wire tmp43419;
  wire tmp43420;
  wire tmp43421;
  wire tmp43422;
  wire tmp43423;
  wire tmp43424;
  wire tmp43425;
  wire tmp43426;
  wire tmp43427;
  wire tmp43428;
  wire tmp43429;
  wire tmp43430;
  wire tmp43431;
  wire tmp43432;
  wire tmp43433;
  wire tmp43434;
  wire tmp43435;
  wire tmp43436;
  wire tmp43437;
  wire tmp43438;
  wire tmp43439;
  wire tmp43440;
  wire tmp43441;
  wire tmp43442;
  wire tmp43443;
  wire tmp43444;
  wire tmp43445;
  wire tmp43446;
  wire tmp43447;
  wire tmp43448;
  wire tmp43449;
  wire tmp43450;
  wire tmp43451;
  wire tmp43452;
  wire tmp43453;
  wire tmp43454;
  wire tmp43455;
  wire tmp43456;
  wire tmp43457;
  wire tmp43458;
  wire tmp43459;
  wire tmp43460;
  wire tmp43461;
  wire tmp43462;
  wire tmp43463;
  wire tmp43464;
  wire tmp43465;
  wire tmp43466;
  wire tmp43467;
  wire tmp43468;
  wire tmp43469;
  wire tmp43470;
  wire tmp43471;
  wire tmp43472;
  wire tmp43473;
  wire tmp43474;
  wire tmp43475;
  wire tmp43476;
  wire tmp43477;
  wire tmp43478;
  wire tmp43479;
  wire tmp43480;
  wire tmp43481;
  wire tmp43482;
  wire tmp43483;
  wire tmp43484;
  wire tmp43485;
  wire tmp43486;
  wire tmp43487;
  wire tmp43488;
  wire tmp43489;
  wire tmp43490;
  wire tmp43491;
  wire tmp43492;
  wire tmp43493;
  wire tmp43494;
  wire tmp43495;
  wire tmp43496;
  wire tmp43497;
  wire tmp43498;
  wire tmp43499;
  wire tmp43500;
  wire tmp43501;
  wire tmp43502;
  wire tmp43503;
  wire tmp43504;
  wire tmp43505;
  wire tmp43506;
  wire tmp43507;
  wire tmp43508;
  wire tmp43509;
  wire tmp43510;
  wire tmp43511;
  wire tmp43512;
  wire tmp43513;
  wire tmp43514;
  wire tmp43515;
  wire tmp43516;
  wire tmp43517;
  wire tmp43518;
  wire tmp43519;
  wire tmp43520;
  wire tmp43521;
  wire tmp43522;
  wire tmp43523;
  wire tmp43524;
  wire tmp43525;
  wire tmp43526;
  wire tmp43527;
  wire tmp43528;
  wire tmp43529;
  wire tmp43530;
  wire tmp43531;
  wire tmp43532;
  wire tmp43533;
  wire tmp43534;
  wire tmp43535;
  wire tmp43536;
  wire tmp43537;
  wire tmp43538;
  wire tmp43539;
  wire tmp43540;
  wire tmp43541;
  wire tmp43542;
  wire tmp43543;
  wire tmp43544;
  wire tmp43545;
  wire tmp43546;
  wire tmp43547;
  wire tmp43548;
  wire tmp43549;
  wire tmp43550;
  wire tmp43551;
  wire tmp43552;
  wire tmp43553;
  wire tmp43554;
  wire tmp43555;
  wire tmp43556;
  wire tmp43557;
  wire tmp43558;
  wire tmp43559;
  wire tmp43560;
  wire tmp43561;
  wire tmp43562;
  wire tmp43563;
  wire tmp43564;
  wire tmp43565;
  wire tmp43566;
  wire tmp43567;
  wire tmp43568;
  wire tmp43569;
  wire tmp43570;
  wire tmp43571;
  wire tmp43572;
  wire tmp43573;
  wire tmp43574;
  wire tmp43575;
  wire tmp43576;
  wire tmp43577;
  wire tmp43578;
  wire tmp43579;
  wire tmp43580;
  wire tmp43581;
  wire tmp43582;
  wire tmp43583;
  wire tmp43584;
  wire tmp43585;
  wire tmp43586;
  wire tmp43587;
  wire tmp43588;
  wire tmp43589;
  wire tmp43590;
  wire tmp43591;
  wire tmp43592;
  wire tmp43593;
  wire tmp43594;
  wire tmp43595;
  wire tmp43596;
  wire tmp43597;
  wire tmp43598;
  wire tmp43599;
  wire tmp43600;
  wire tmp43601;
  wire tmp43602;
  wire tmp43603;
  wire tmp43604;
  wire tmp43605;
  wire tmp43606;
  wire tmp43607;
  wire tmp43608;
  wire tmp43609;
  wire tmp43610;
  wire tmp43611;
  wire tmp43612;
  wire tmp43613;
  wire tmp43614;
  wire tmp43615;
  wire tmp43616;
  wire tmp43617;
  wire tmp43618;
  wire tmp43619;
  wire tmp43620;
  wire tmp43621;
  wire tmp43622;
  wire tmp43623;
  wire tmp43624;
  wire tmp43625;
  wire tmp43626;
  wire tmp43627;
  wire tmp43628;
  wire tmp43629;
  wire tmp43630;
  wire tmp43631;
  wire tmp43632;
  wire tmp43633;
  wire tmp43634;
  wire tmp43635;
  wire tmp43636;
  wire tmp43637;
  wire tmp43638;
  wire tmp43639;
  wire tmp43640;
  wire tmp43641;
  wire tmp43642;
  wire tmp43643;
  wire tmp43644;
  wire tmp43645;
  wire tmp43646;
  wire tmp43647;
  wire tmp43648;
  wire tmp43649;
  wire tmp43650;
  wire tmp43651;
  wire tmp43652;
  wire tmp43653;
  wire tmp43654;
  wire tmp43655;
  wire tmp43656;
  wire tmp43657;
  wire tmp43658;
  wire tmp43659;
  wire tmp43660;
  wire tmp43661;
  wire tmp43662;
  wire tmp43663;
  wire tmp43664;
  wire tmp43665;
  wire tmp43666;
  wire tmp43667;
  wire tmp43668;
  wire tmp43669;
  wire tmp43670;
  wire tmp43671;
  wire tmp43672;
  wire tmp43673;
  wire tmp43674;
  wire tmp43675;
  wire tmp43676;
  wire tmp43677;
  wire tmp43678;
  wire tmp43679;
  wire tmp43680;
  wire tmp43681;
  wire tmp43682;
  wire tmp43683;
  wire tmp43684;
  wire tmp43685;
  wire tmp43686;
  wire tmp43687;
  wire tmp43688;
  wire tmp43689;
  wire tmp43690;
  wire tmp43691;
  wire tmp43692;
  wire tmp43693;
  wire tmp43694;
  wire tmp43695;
  wire tmp43696;
  wire tmp43697;
  wire tmp43698;
  wire tmp43699;
  wire tmp43700;
  wire tmp43701;
  wire tmp43702;
  wire tmp43703;
  wire tmp43704;
  wire tmp43705;
  wire tmp43706;
  wire tmp43707;
  wire tmp43708;
  wire tmp43709;
  wire tmp43710;
  wire tmp43711;
  wire tmp43712;
  wire tmp43713;
  wire tmp43714;
  wire tmp43715;
  wire tmp43716;
  wire tmp43717;
  wire tmp43718;
  wire tmp43719;
  wire tmp43720;
  wire tmp43721;
  wire tmp43722;
  wire tmp43723;
  wire tmp43724;
  wire tmp43725;
  wire tmp43726;
  wire tmp43727;
  wire tmp43728;
  wire tmp43729;
  wire tmp43730;
  wire tmp43731;
  wire tmp43732;
  wire tmp43733;
  wire tmp43734;
  wire tmp43735;
  wire tmp43736;
  wire tmp43737;
  wire tmp43738;
  wire tmp43739;
  wire tmp43740;
  wire tmp43741;
  wire tmp43742;
  wire tmp43743;
  wire tmp43744;
  wire tmp43745;
  wire tmp43746;
  wire tmp43747;
  wire tmp43748;
  wire tmp43749;
  wire tmp43750;
  wire tmp43751;
  wire tmp43752;
  wire tmp43753;
  wire tmp43754;
  wire tmp43755;
  wire tmp43756;
  wire tmp43757;
  wire tmp43758;
  wire tmp43759;
  wire tmp43760;
  wire tmp43761;
  wire tmp43762;
  wire tmp43763;
  wire tmp43764;
  wire tmp43765;
  wire tmp43766;
  wire tmp43767;
  wire tmp43768;
  wire tmp43769;
  wire tmp43770;
  wire tmp43771;
  wire tmp43772;
  wire tmp43773;
  wire tmp43774;
  wire tmp43775;
  wire tmp43776;
  wire tmp43777;
  wire tmp43778;
  wire tmp43779;
  wire tmp43780;
  wire tmp43781;
  wire tmp43782;
  wire tmp43783;
  wire tmp43784;
  wire tmp43785;
  wire tmp43786;
  wire tmp43787;
  wire tmp43788;
  wire tmp43789;
  wire tmp43790;
  wire tmp43791;
  wire tmp43792;
  wire tmp43793;
  wire tmp43794;
  wire tmp43795;
  wire tmp43796;
  wire tmp43797;
  wire tmp43798;
  wire tmp43799;
  wire tmp43800;
  wire tmp43801;
  wire tmp43802;
  wire tmp43803;
  wire tmp43804;
  wire tmp43805;
  wire tmp43806;
  wire tmp43807;
  wire tmp43808;
  wire tmp43809;
  wire tmp43810;
  wire tmp43811;
  wire tmp43812;
  wire tmp43813;
  wire tmp43814;
  wire tmp43815;
  wire tmp43816;
  wire tmp43817;
  wire tmp43818;
  wire tmp43819;
  wire tmp43820;
  wire tmp43821;
  wire tmp43822;
  wire tmp43823;
  wire tmp43824;
  wire tmp43825;
  wire tmp43826;
  wire tmp43827;
  wire tmp43828;
  wire tmp43829;
  wire tmp43830;
  wire tmp43831;
  wire tmp43832;
  wire tmp43833;
  wire tmp43834;
  wire tmp43835;
  wire tmp43836;
  wire tmp43837;
  wire tmp43838;
  wire tmp43839;
  wire tmp43840;
  wire tmp43841;
  wire tmp43842;
  wire tmp43843;
  wire tmp43844;
  wire tmp43845;
  wire tmp43846;
  wire tmp43847;
  wire tmp43848;
  wire tmp43849;
  wire tmp43850;
  wire tmp43851;
  wire tmp43852;
  wire tmp43853;
  wire tmp43854;
  wire tmp43855;
  wire tmp43856;
  wire tmp43857;
  wire tmp43858;
  wire tmp43859;
  wire tmp43860;
  wire tmp43861;
  wire tmp43862;
  wire tmp43863;
  wire tmp43864;
  wire tmp43865;
  wire tmp43866;
  wire tmp43867;
  wire tmp43868;
  wire tmp43869;
  wire tmp43870;
  wire tmp43871;
  wire tmp43872;
  wire tmp43873;
  wire tmp43874;
  wire tmp43875;
  wire tmp43876;
  wire tmp43877;
  wire tmp43878;
  wire tmp43879;
  wire tmp43880;
  wire tmp43881;
  wire tmp43882;
  wire tmp43883;
  wire tmp43884;
  wire tmp43885;
  wire tmp43886;
  wire tmp43887;
  wire tmp43888;
  wire tmp43889;
  wire tmp43890;
  wire tmp43891;
  wire tmp43892;
  wire tmp43893;
  wire tmp43894;
  wire tmp43895;
  wire tmp43896;
  wire tmp43897;
  wire tmp43898;
  wire tmp43899;
  wire tmp43900;
  wire tmp43901;
  wire tmp43902;
  wire tmp43903;
  wire tmp43904;
  wire tmp43905;
  wire tmp43906;
  wire tmp43907;
  wire tmp43908;
  wire tmp43909;
  wire tmp43910;
  wire tmp43911;
  wire tmp43912;
  wire tmp43913;
  wire tmp43914;
  wire tmp43915;
  wire tmp43916;
  wire tmp43917;
  wire tmp43918;
  wire tmp43919;
  wire tmp43920;
  wire tmp43921;
  wire tmp43922;
  wire tmp43923;
  wire tmp43924;
  wire tmp43925;
  wire tmp43926;
  wire tmp43927;
  wire tmp43928;
  wire tmp43929;
  wire tmp43930;
  wire tmp43931;
  wire tmp43932;
  wire tmp43933;
  wire tmp43934;
  wire tmp43935;
  wire tmp43936;
  wire tmp43937;
  wire tmp43938;
  wire tmp43939;
  wire tmp43940;
  wire tmp43941;
  wire tmp43942;
  wire tmp43943;
  wire tmp43944;
  wire tmp43945;
  wire tmp43946;
  wire tmp43947;
  wire tmp43948;
  wire tmp43949;
  wire tmp43950;
  wire tmp43951;
  wire tmp43952;
  wire tmp43953;
  wire tmp43954;
  wire tmp43955;
  wire tmp43956;
  wire tmp43957;
  wire tmp43958;
  wire tmp43959;
  wire tmp43960;
  wire tmp43961;
  wire tmp43962;
  wire tmp43963;
  wire tmp43964;
  wire tmp43965;
  wire tmp43966;
  wire tmp43967;
  wire tmp43968;
  wire tmp43969;
  wire tmp43970;
  wire tmp43971;
  wire tmp43972;
  wire tmp43973;
  wire tmp43974;
  wire tmp43975;
  wire tmp43976;
  wire tmp43977;
  wire tmp43978;
  wire tmp43979;
  wire tmp43980;
  wire tmp43981;
  wire tmp43982;
  wire tmp43983;
  wire tmp43984;
  wire tmp43985;
  wire tmp43986;
  wire tmp43987;
  wire tmp43988;
  wire tmp43989;
  wire tmp43990;
  wire tmp43991;
  wire tmp43992;
  wire tmp43993;
  wire tmp43994;
  wire tmp43995;
  wire tmp43996;
  wire tmp43997;
  wire tmp43998;
  wire tmp43999;
  wire tmp44000;
  wire tmp44001;
  wire tmp44002;
  wire tmp44003;
  wire tmp44004;
  wire tmp44005;
  wire tmp44006;
  wire tmp44007;
  wire tmp44008;
  wire tmp44009;
  wire tmp44010;
  wire tmp44011;
  wire tmp44012;
  wire tmp44013;
  wire tmp44014;
  wire tmp44015;
  wire tmp44016;
  wire tmp44017;
  wire tmp44018;
  wire tmp44019;
  wire tmp44020;
  wire tmp44021;
  wire tmp44022;
  wire tmp44023;
  wire tmp44024;
  wire tmp44025;
  wire tmp44026;
  wire tmp44027;
  wire tmp44028;
  wire tmp44029;
  wire tmp44030;
  wire tmp44031;
  wire tmp44032;
  wire tmp44033;
  wire tmp44034;
  wire tmp44035;
  wire tmp44036;
  wire tmp44037;
  wire tmp44038;
  wire tmp44039;
  wire tmp44040;
  wire tmp44041;
  wire tmp44042;
  wire tmp44043;
  wire tmp44044;
  wire tmp44045;
  wire tmp44046;
  wire tmp44047;
  wire tmp44048;
  wire tmp44049;
  wire tmp44050;
  wire tmp44051;
  wire tmp44052;
  wire tmp44053;
  wire tmp44054;
  wire tmp44055;
  wire tmp44056;
  wire tmp44057;
  wire tmp44058;
  wire tmp44059;
  wire tmp44060;
  wire tmp44061;
  wire tmp44062;
  wire tmp44063;
  wire tmp44064;
  wire tmp44065;
  wire tmp44066;
  wire tmp44067;
  wire tmp44068;
  wire tmp44069;
  wire tmp44070;
  wire tmp44071;
  wire tmp44072;
  wire tmp44073;
  wire tmp44074;
  wire tmp44075;
  wire tmp44076;
  wire tmp44077;
  wire tmp44078;
  wire tmp44079;
  wire tmp44080;
  wire tmp44081;
  wire tmp44082;
  wire tmp44083;
  wire tmp44084;
  wire tmp44085;
  wire tmp44086;
  wire tmp44087;
  wire tmp44088;
  wire tmp44089;
  wire tmp44090;
  wire tmp44091;
  wire tmp44092;
  wire tmp44093;
  wire tmp44094;
  wire tmp44095;
  wire tmp44096;
  wire tmp44097;
  wire tmp44098;
  wire tmp44099;
  wire tmp44100;
  wire tmp44101;
  wire tmp44102;
  wire tmp44103;
  wire tmp44104;
  wire tmp44105;
  wire tmp44106;
  wire tmp44107;
  wire tmp44108;
  wire tmp44109;
  wire tmp44110;
  wire tmp44111;
  wire tmp44112;
  wire tmp44113;
  wire tmp44114;
  wire tmp44115;
  wire tmp44116;
  wire tmp44117;
  wire tmp44118;
  wire tmp44119;
  wire tmp44120;
  wire tmp44121;
  wire tmp44122;
  wire tmp44123;
  wire tmp44124;
  wire tmp44125;
  wire tmp44126;
  wire tmp44127;
  wire tmp44128;
  wire tmp44129;
  wire tmp44130;
  wire tmp44131;
  wire tmp44132;
  wire tmp44133;
  wire tmp44134;
  wire tmp44135;
  wire tmp44136;
  wire tmp44137;
  wire tmp44138;
  wire tmp44139;
  wire tmp44140;
  wire tmp44141;
  wire tmp44142;
  wire tmp44143;
  wire tmp44144;
  wire tmp44145;
  wire tmp44146;
  wire tmp44147;
  wire tmp44148;
  wire tmp44149;
  wire tmp44150;
  wire tmp44151;
  wire tmp44152;
  wire tmp44153;
  wire tmp44154;
  wire tmp44155;
  wire tmp44156;
  wire tmp44157;
  wire tmp44158;
  wire tmp44159;
  wire tmp44160;
  wire tmp44161;
  wire tmp44162;
  wire tmp44163;
  wire tmp44164;
  wire tmp44165;
  wire tmp44166;
  wire tmp44167;
  wire tmp44168;
  wire tmp44169;
  wire tmp44170;
  wire tmp44171;
  wire tmp44172;
  wire tmp44173;
  wire tmp44174;
  wire tmp44175;
  wire tmp44176;
  wire tmp44177;
  wire tmp44178;
  wire tmp44179;
  wire tmp44180;
  wire tmp44181;
  wire tmp44182;
  wire tmp44183;
  wire tmp44184;
  wire tmp44185;
  wire tmp44186;
  wire tmp44187;
  wire tmp44188;
  wire tmp44189;
  wire tmp44190;
  wire tmp44191;
  wire tmp44192;
  wire tmp44193;
  wire tmp44194;
  wire tmp44195;
  wire tmp44196;
  wire tmp44197;
  wire tmp44198;
  wire tmp44199;
  wire tmp44200;
  wire tmp44201;
  wire tmp44202;
  wire tmp44203;
  wire tmp44204;
  wire tmp44205;
  wire tmp44206;
  wire tmp44207;
  wire tmp44208;
  wire tmp44209;
  wire tmp44210;
  wire tmp44211;
  wire tmp44212;
  wire tmp44213;
  wire tmp44214;
  wire tmp44215;
  wire tmp44216;
  wire tmp44217;
  wire tmp44218;
  wire tmp44219;
  wire tmp44220;
  wire tmp44221;
  wire tmp44222;
  wire tmp44223;
  wire tmp44224;
  wire tmp44225;
  wire tmp44226;
  wire tmp44227;
  wire tmp44228;
  wire tmp44229;
  wire tmp44230;
  wire tmp44231;
  wire tmp44232;
  wire tmp44233;
  wire tmp44234;
  wire tmp44235;
  wire tmp44236;
  wire tmp44237;
  wire tmp44238;
  wire tmp44239;
  wire tmp44240;
  wire tmp44241;
  wire tmp44242;
  wire tmp44243;
  wire tmp44244;
  wire tmp44245;
  wire tmp44246;
  wire tmp44247;
  wire tmp44248;
  wire tmp44249;
  wire tmp44250;
  wire tmp44251;
  wire tmp44252;
  wire tmp44253;
  wire tmp44254;
  wire tmp44255;
  wire tmp44256;
  wire tmp44257;
  wire tmp44258;
  wire tmp44259;
  wire tmp44260;
  wire tmp44261;
  wire tmp44262;
  wire tmp44263;
  wire tmp44264;
  wire tmp44265;
  wire tmp44266;
  wire tmp44267;
  wire tmp44268;
  wire tmp44269;
  wire tmp44270;
  wire tmp44271;
  wire tmp44272;
  wire tmp44273;
  wire tmp44274;
  wire tmp44275;
  wire tmp44276;
  wire tmp44277;
  wire tmp44278;
  wire tmp44279;
  wire tmp44280;
  wire tmp44281;
  wire tmp44282;
  wire tmp44283;
  wire tmp44284;
  wire tmp44285;
  wire tmp44286;
  wire tmp44287;
  wire tmp44288;
  wire tmp44289;
  wire tmp44290;
  wire tmp44291;
  wire tmp44292;
  wire tmp44293;
  wire tmp44294;
  wire tmp44295;
  wire tmp44296;
  wire tmp44297;
  wire tmp44298;
  wire tmp44299;
  wire tmp44300;
  wire tmp44301;
  wire tmp44302;
  wire tmp44303;
  wire tmp44304;
  wire tmp44305;
  wire tmp44306;
  wire tmp44307;
  wire tmp44308;
  wire tmp44309;
  wire tmp44310;
  wire tmp44311;
  wire tmp44312;
  wire tmp44313;
  wire tmp44314;
  wire tmp44315;
  wire tmp44316;
  wire tmp44317;
  wire tmp44318;
  wire tmp44319;
  wire tmp44320;
  wire tmp44321;
  wire tmp44322;
  wire tmp44323;
  wire tmp44324;
  wire tmp44325;
  wire tmp44326;
  wire tmp44327;
  wire tmp44328;
  wire tmp44329;
  wire tmp44330;
  wire tmp44331;
  wire tmp44332;
  wire tmp44333;
  wire tmp44334;
  wire tmp44335;
  wire tmp44336;
  wire tmp44337;
  wire tmp44338;
  wire tmp44339;
  wire tmp44340;
  wire tmp44341;
  wire tmp44342;
  wire tmp44343;
  wire tmp44344;
  wire tmp44345;
  wire tmp44346;
  wire tmp44347;
  wire tmp44348;
  wire tmp44349;
  wire tmp44350;
  wire tmp44351;
  wire tmp44352;
  wire tmp44353;
  wire tmp44354;
  wire tmp44355;
  wire tmp44356;
  wire tmp44357;
  wire tmp44358;
  wire tmp44359;
  wire tmp44360;
  wire tmp44361;
  wire tmp44362;
  wire tmp44363;
  wire tmp44364;
  wire tmp44365;
  wire tmp44366;
  wire tmp44367;
  wire tmp44368;
  wire tmp44369;
  wire tmp44370;
  wire tmp44371;
  wire tmp44372;
  wire tmp44373;
  wire tmp44374;
  wire tmp44375;
  wire tmp44376;
  wire tmp44377;
  wire tmp44378;
  wire tmp44379;
  wire tmp44380;
  wire tmp44381;
  wire tmp44382;
  wire tmp44383;
  wire tmp44384;
  wire tmp44385;
  wire tmp44386;
  wire tmp44387;
  wire tmp44388;
  wire tmp44389;
  wire tmp44390;
  wire tmp44391;
  wire tmp44392;
  wire tmp44393;
  wire tmp44394;
  wire tmp44395;
  wire tmp44396;
  wire tmp44397;
  wire tmp44398;
  wire tmp44399;
  wire tmp44400;
  wire tmp44401;
  wire tmp44402;
  wire tmp44403;
  wire tmp44404;
  wire tmp44405;
  wire tmp44406;
  wire tmp44407;
  wire tmp44408;
  wire tmp44409;
  wire tmp44410;
  wire tmp44411;
  wire tmp44412;
  wire tmp44413;
  wire tmp44414;
  wire tmp44415;
  wire tmp44416;
  wire tmp44417;
  wire tmp44418;
  wire tmp44419;
  wire tmp44420;
  wire tmp44421;
  wire tmp44422;
  wire tmp44423;
  wire tmp44424;
  wire tmp44425;
  wire tmp44426;
  wire tmp44427;
  wire tmp44428;
  wire tmp44429;
  wire tmp44430;
  wire tmp44431;
  wire tmp44432;
  wire tmp44433;
  wire tmp44434;
  wire tmp44435;
  wire tmp44436;
  wire tmp44437;
  wire tmp44438;
  wire tmp44439;
  wire tmp44440;
  wire tmp44441;
  wire tmp44442;
  wire tmp44443;
  wire tmp44444;
  wire tmp44445;
  wire tmp44446;
  wire tmp44447;
  wire tmp44448;
  wire tmp44449;
  wire tmp44450;
  wire tmp44451;
  wire tmp44452;
  wire tmp44453;
  wire tmp44454;
  wire tmp44455;
  wire tmp44456;
  wire tmp44457;
  wire tmp44458;
  wire tmp44459;
  wire tmp44460;
  wire tmp44461;
  wire tmp44462;
  wire tmp44463;
  wire tmp44464;
  wire tmp44465;
  wire tmp44466;
  wire tmp44467;
  wire tmp44468;
  wire tmp44469;
  wire tmp44470;
  wire tmp44471;
  wire tmp44472;
  wire tmp44473;
  wire tmp44474;
  wire tmp44475;
  wire tmp44476;
  wire tmp44477;
  wire tmp44478;
  wire tmp44479;
  wire tmp44480;
  wire tmp44481;
  wire tmp44482;
  wire tmp44483;
  wire tmp44484;
  wire tmp44485;
  wire tmp44486;
  wire tmp44487;
  wire tmp44488;
  wire tmp44489;
  wire tmp44490;
  wire tmp44491;
  wire tmp44492;
  wire tmp44493;
  wire tmp44494;
  wire tmp44495;
  wire tmp44496;
  wire tmp44497;
  wire tmp44498;
  wire tmp44499;
  wire tmp44500;
  wire tmp44501;
  wire tmp44502;
  wire tmp44503;
  wire tmp44504;
  wire tmp44505;
  wire tmp44506;
  wire tmp44507;
  wire tmp44508;
  wire tmp44509;
  wire tmp44510;
  wire tmp44511;
  wire tmp44512;
  wire tmp44513;
  wire tmp44514;
  wire tmp44515;
  wire tmp44516;
  wire tmp44517;
  wire tmp44518;
  wire tmp44519;
  wire tmp44520;
  wire tmp44521;
  wire tmp44522;
  wire tmp44523;
  wire tmp44524;
  wire tmp44525;
  wire tmp44526;
  wire tmp44527;
  wire tmp44528;
  wire tmp44529;
  wire tmp44530;
  wire tmp44531;
  wire tmp44532;
  wire tmp44533;
  wire tmp44534;
  wire tmp44535;
  wire tmp44536;
  wire tmp44537;
  wire tmp44538;
  wire tmp44539;
  wire tmp44540;
  wire tmp44541;
  wire tmp44542;
  wire tmp44543;
  wire tmp44544;
  wire tmp44545;
  wire tmp44546;
  wire tmp44547;
  wire tmp44548;
  wire tmp44549;
  wire tmp44550;
  wire tmp44551;
  wire tmp44552;
  wire tmp44553;
  wire tmp44554;
  wire tmp44555;
  wire tmp44556;
  wire tmp44557;
  wire tmp44558;
  wire tmp44559;
  wire tmp44560;
  wire tmp44561;
  wire tmp44562;
  wire tmp44563;
  wire tmp44564;
  wire tmp44565;
  wire tmp44566;
  wire tmp44567;
  wire tmp44568;
  wire tmp44569;
  wire tmp44570;
  wire tmp44571;
  wire tmp44572;
  wire tmp44573;
  wire tmp44574;
  wire tmp44575;
  wire tmp44576;
  wire tmp44577;
  wire tmp44578;
  wire tmp44579;
  wire tmp44580;
  wire tmp44581;
  wire tmp44582;
  wire tmp44583;
  wire tmp44584;
  wire tmp44585;
  wire tmp44586;
  wire tmp44587;
  wire tmp44588;
  wire tmp44589;
  wire tmp44590;
  wire tmp44591;
  wire tmp44592;
  wire tmp44593;
  wire tmp44594;
  wire tmp44595;
  wire tmp44596;
  wire tmp44597;
  wire tmp44598;
  wire tmp44599;
  wire tmp44600;
  wire tmp44601;
  wire tmp44602;
  wire tmp44603;
  wire tmp44604;
  wire tmp44605;
  wire tmp44606;
  wire tmp44607;
  wire tmp44608;
  wire tmp44609;
  wire tmp44610;
  wire tmp44611;
  wire tmp44612;
  wire tmp44613;
  wire tmp44614;
  wire tmp44615;
  wire tmp44616;
  wire tmp44617;
  wire tmp44618;
  wire tmp44619;
  wire tmp44620;
  wire tmp44621;
  wire tmp44622;
  wire tmp44623;
  wire tmp44624;
  wire tmp44625;
  wire tmp44626;
  wire tmp44627;
  wire tmp44628;
  wire tmp44629;
  wire tmp44630;
  wire tmp44631;
  wire tmp44632;
  wire tmp44633;
  wire tmp44634;
  wire tmp44635;
  wire tmp44636;
  wire tmp44637;
  wire tmp44638;
  wire tmp44639;
  wire tmp44640;
  wire tmp44641;
  wire tmp44642;
  wire tmp44643;
  wire tmp44644;
  wire tmp44645;
  wire tmp44646;
  wire tmp44647;
  wire tmp44648;
  wire tmp44649;
  wire tmp44650;
  wire tmp44651;
  wire tmp44652;
  wire tmp44653;
  wire tmp44654;
  wire tmp44655;
  wire tmp44656;
  wire tmp44657;
  wire tmp44658;
  wire tmp44659;
  wire tmp44660;
  wire tmp44661;
  wire tmp44662;
  wire tmp44663;
  wire tmp44664;
  wire tmp44665;
  wire tmp44666;
  wire tmp44667;
  wire tmp44668;
  wire tmp44669;
  wire tmp44670;
  wire tmp44671;
  wire tmp44672;
  wire tmp44673;
  wire tmp44674;
  wire tmp44675;
  wire tmp44676;
  wire tmp44677;
  wire tmp44678;
  wire tmp44679;
  wire tmp44680;
  wire tmp44681;
  wire tmp44682;
  wire tmp44683;
  wire tmp44684;
  wire tmp44685;
  wire tmp44686;
  wire tmp44687;
  wire tmp44688;
  wire tmp44689;
  wire tmp44690;
  wire tmp44691;
  wire tmp44692;
  wire tmp44693;
  wire tmp44694;
  wire tmp44695;
  wire tmp44696;
  wire tmp44697;
  wire tmp44698;
  wire tmp44699;
  wire tmp44700;
  wire tmp44701;
  wire tmp44702;
  wire tmp44703;
  wire tmp44704;
  wire tmp44705;
  wire tmp44706;
  wire tmp44707;
  wire tmp44708;
  wire tmp44709;
  wire tmp44710;
  wire tmp44711;
  wire tmp44712;
  wire tmp44713;
  wire tmp44714;
  wire tmp44715;
  wire tmp44716;
  wire tmp44717;
  wire tmp44718;
  wire tmp44719;
  wire tmp44720;
  wire tmp44721;
  wire tmp44722;
  wire tmp44723;
  wire tmp44724;
  wire tmp44725;
  wire tmp44726;
  wire tmp44727;
  wire tmp44728;
  wire tmp44729;
  wire tmp44730;
  wire tmp44731;
  wire tmp44732;
  wire tmp44733;
  wire tmp44734;
  wire tmp44735;
  wire tmp44736;
  wire tmp44737;
  wire tmp44738;
  wire tmp44739;
  wire tmp44740;
  wire tmp44741;
  wire tmp44742;
  wire tmp44743;
  wire tmp44744;
  wire tmp44745;
  wire tmp44746;
  wire tmp44747;
  wire tmp44748;
  wire tmp44749;
  wire tmp44750;
  wire tmp44751;
  wire tmp44752;
  wire tmp44753;
  wire tmp44754;
  wire tmp44755;
  wire tmp44756;
  wire tmp44757;
  wire tmp44758;
  wire tmp44759;
  wire tmp44760;
  wire tmp44761;
  wire tmp44762;
  wire tmp44763;
  wire tmp44764;
  wire tmp44765;
  wire tmp44766;
  wire tmp44767;
  wire tmp44768;
  wire tmp44769;
  wire tmp44770;
  wire tmp44771;
  wire tmp44772;
  wire tmp44773;
  wire tmp44774;
  wire tmp44775;
  wire tmp44776;
  wire tmp44777;
  wire tmp44778;
  wire tmp44779;
  wire tmp44780;
  wire tmp44781;
  wire tmp44782;
  wire tmp44783;
  wire tmp44784;
  wire tmp44785;
  wire tmp44786;
  wire tmp44787;
  wire tmp44788;
  wire tmp44789;
  wire tmp44790;
  wire tmp44791;
  wire tmp44792;
  wire tmp44793;
  wire tmp44794;
  wire tmp44795;
  wire tmp44796;
  wire tmp44797;
  wire tmp44798;
  wire tmp44799;
  wire tmp44800;
  wire tmp44801;
  wire tmp44802;
  wire tmp44803;
  wire tmp44804;
  wire tmp44805;
  wire tmp44806;
  wire tmp44807;
  wire tmp44808;
  wire tmp44809;
  wire tmp44810;
  wire tmp44811;
  wire tmp44812;
  wire tmp44813;
  wire tmp44814;
  wire tmp44815;
  wire tmp44816;
  wire tmp44817;
  wire tmp44818;
  wire tmp44819;
  wire tmp44820;
  wire tmp44821;
  wire tmp44822;
  wire tmp44823;
  wire tmp44824;
  wire tmp44825;
  wire tmp44826;
  wire tmp44827;
  wire tmp44828;
  wire tmp44829;
  wire tmp44830;
  wire tmp44831;
  wire tmp44832;
  wire tmp44833;
  wire tmp44834;
  wire tmp44835;
  wire tmp44836;
  wire tmp44837;
  wire tmp44838;
  wire tmp44839;
  wire tmp44840;
  wire tmp44841;
  wire tmp44842;
  wire tmp44843;
  wire tmp44844;
  wire tmp44845;
  wire tmp44846;
  wire tmp44847;
  wire tmp44848;
  wire tmp44849;
  wire tmp44850;
  wire tmp44851;
  wire tmp44852;
  wire tmp44853;
  wire tmp44854;
  wire tmp44855;
  wire tmp44856;
  wire tmp44857;
  wire tmp44858;
  wire tmp44859;
  wire tmp44860;
  wire tmp44861;
  wire tmp44862;
  wire tmp44863;
  wire tmp44864;
  wire tmp44865;
  wire tmp44866;
  wire tmp44867;
  wire tmp44868;
  wire tmp44869;
  wire tmp44870;
  wire tmp44871;
  wire tmp44872;
  wire tmp44873;
  wire tmp44874;
  wire tmp44875;
  wire tmp44876;
  wire tmp44877;
  wire tmp44878;
  wire tmp44879;
  wire tmp44880;
  wire tmp44881;
  wire tmp44882;
  wire tmp44883;
  wire tmp44884;
  wire tmp44885;
  wire tmp44886;
  wire tmp44887;
  wire tmp44888;
  wire tmp44889;
  wire tmp44890;
  wire tmp44891;
  wire tmp44892;
  wire tmp44893;
  wire tmp44894;
  wire tmp44895;
  wire tmp44896;
  wire tmp44897;
  wire tmp44898;
  wire tmp44899;
  wire tmp44900;
  wire tmp44901;
  wire tmp44902;
  wire tmp44903;
  wire tmp44904;
  wire tmp44905;
  wire tmp44906;
  wire tmp44907;
  wire tmp44908;
  wire tmp44909;
  wire tmp44910;
  wire tmp44911;
  wire tmp44912;
  wire tmp44913;
  wire tmp44914;
  wire tmp44915;
  wire tmp44916;
  wire tmp44917;
  wire tmp44918;
  wire tmp44919;
  wire tmp44920;
  wire tmp44921;
  wire tmp44922;
  wire tmp44923;
  wire tmp44924;
  wire tmp44925;
  wire tmp44926;
  wire tmp44927;
  wire tmp44928;
  wire tmp44929;
  wire tmp44930;
  wire tmp44931;
  wire tmp44932;
  wire tmp44933;
  wire tmp44934;
  wire tmp44935;
  wire tmp44936;
  wire tmp44937;
  wire tmp44938;
  wire tmp44939;
  wire tmp44940;
  wire tmp44941;
  wire tmp44942;
  wire tmp44943;
  wire tmp44944;
  wire tmp44945;
  wire tmp44946;
  wire tmp44947;
  wire tmp44948;
  wire tmp44949;
  wire tmp44950;
  wire tmp44951;
  wire tmp44952;
  wire tmp44953;
  wire tmp44954;
  wire tmp44955;
  wire tmp44956;
  wire tmp44957;
  wire tmp44958;
  wire tmp44959;
  wire tmp44960;
  wire tmp44961;
  wire tmp44962;
  wire tmp44963;
  wire tmp44964;
  wire tmp44965;
  wire tmp44966;
  wire tmp44967;
  wire tmp44968;
  wire tmp44969;
  wire tmp44970;
  wire tmp44971;
  wire tmp44972;
  wire tmp44973;
  wire tmp44974;
  wire tmp44975;
  wire tmp44976;
  wire tmp44977;
  wire tmp44978;
  wire tmp44979;
  wire tmp44980;
  wire tmp44981;
  wire tmp44982;
  wire tmp44983;
  wire tmp44984;
  wire tmp44985;
  wire tmp44986;
  wire tmp44987;
  wire tmp44988;
  wire tmp44989;
  wire tmp44990;
  wire tmp44991;
  wire tmp44992;
  wire tmp44993;
  wire tmp44994;
  wire tmp44995;
  wire tmp44996;
  wire tmp44997;
  wire tmp44998;
  wire tmp44999;
  wire tmp45000;
  wire tmp45001;
  wire tmp45002;
  wire tmp45003;
  wire tmp45004;
  wire tmp45005;
  wire tmp45006;
  wire tmp45007;
  wire tmp45008;
  wire tmp45009;
  wire tmp45010;
  wire tmp45011;
  wire tmp45012;
  wire tmp45013;
  wire tmp45014;
  wire tmp45015;
  wire tmp45016;
  wire tmp45017;
  wire tmp45018;
  wire tmp45019;
  wire tmp45020;
  wire tmp45021;
  wire tmp45022;
  wire tmp45023;
  wire tmp45024;
  wire tmp45025;
  wire tmp45026;
  wire tmp45027;
  wire tmp45028;
  wire tmp45029;
  wire tmp45030;
  wire tmp45031;
  wire tmp45032;
  wire tmp45033;
  wire tmp45034;
  wire tmp45035;
  wire tmp45036;
  wire tmp45037;
  wire tmp45038;
  wire tmp45039;
  wire tmp45040;
  wire tmp45041;
  wire tmp45042;
  wire tmp45043;
  wire tmp45044;
  wire tmp45045;
  wire tmp45046;
  wire tmp45047;
  wire tmp45048;
  wire tmp45049;
  wire tmp45050;
  wire tmp45051;
  wire tmp45052;
  wire tmp45053;
  wire tmp45054;
  wire tmp45055;
  wire tmp45056;
  wire tmp45057;
  wire tmp45058;
  wire tmp45059;
  wire tmp45060;
  wire tmp45061;
  wire tmp45062;
  wire tmp45063;
  wire tmp45064;
  wire tmp45065;
  wire tmp45066;
  wire tmp45067;
  wire tmp45068;
  wire tmp45069;
  wire tmp45070;
  wire tmp45071;
  wire tmp45072;
  wire tmp45073;
  wire tmp45074;
  wire tmp45075;
  wire tmp45076;
  wire tmp45077;
  wire tmp45078;
  wire tmp45079;
  wire tmp45080;
  wire tmp45081;
  wire tmp45082;
  wire tmp45083;
  wire tmp45084;
  wire tmp45085;
  wire tmp45086;
  wire tmp45087;
  wire tmp45088;
  wire tmp45089;
  wire tmp45090;
  wire tmp45091;
  wire tmp45092;
  wire tmp45093;
  wire tmp45094;
  wire tmp45095;
  wire tmp45096;
  wire tmp45097;
  wire tmp45098;
  wire tmp45099;
  wire tmp45100;
  wire tmp45101;
  wire tmp45102;
  wire tmp45103;
  wire tmp45104;
  wire tmp45105;
  wire tmp45106;
  wire tmp45107;
  wire tmp45108;
  wire tmp45109;
  wire tmp45110;
  wire tmp45111;
  wire tmp45112;
  wire tmp45113;
  wire tmp45114;
  wire tmp45115;
  wire tmp45116;
  wire tmp45117;
  wire tmp45118;
  wire tmp45119;
  wire tmp45120;
  wire tmp45121;
  wire tmp45122;
  wire tmp45123;
  wire tmp45124;
  wire tmp45125;
  wire tmp45126;
  wire tmp45127;
  wire tmp45128;
  wire tmp45129;
  wire tmp45130;
  wire tmp45131;
  wire tmp45132;
  wire tmp45133;
  wire tmp45134;
  wire tmp45135;
  wire tmp45136;
  wire tmp45137;
  wire tmp45138;
  wire tmp45139;
  wire tmp45140;
  wire tmp45141;
  wire tmp45142;
  wire tmp45143;
  wire tmp45144;
  wire tmp45145;
  wire tmp45146;
  wire tmp45147;
  wire tmp45148;
  wire tmp45149;
  wire tmp45150;
  wire tmp45151;
  wire tmp45152;
  wire tmp45153;
  wire tmp45154;
  wire tmp45155;
  wire tmp45156;
  wire tmp45157;
  wire tmp45158;
  wire tmp45159;
  wire tmp45160;
  wire tmp45161;
  wire tmp45162;
  wire tmp45163;
  wire tmp45164;
  wire tmp45165;
  wire tmp45166;
  wire tmp45167;
  wire tmp45168;
  wire tmp45169;
  wire tmp45170;
  wire tmp45171;
  wire tmp45172;
  wire tmp45173;
  wire tmp45174;
  wire tmp45175;
  wire tmp45176;
  wire tmp45177;
  wire tmp45178;
  wire tmp45179;
  wire tmp45180;
  wire tmp45181;
  wire tmp45182;
  wire tmp45183;
  wire tmp45184;
  wire tmp45185;
  wire tmp45186;
  wire tmp45187;
  wire tmp45188;
  wire tmp45189;
  wire tmp45190;
  wire tmp45191;
  wire tmp45192;
  wire tmp45193;
  wire tmp45194;
  wire tmp45195;
  wire tmp45196;
  wire tmp45197;
  wire tmp45198;
  wire tmp45199;
  wire tmp45200;
  wire tmp45201;
  wire tmp45202;
  wire tmp45203;
  wire tmp45204;
  wire tmp45205;
  wire tmp45206;
  wire tmp45207;
  wire tmp45208;
  wire tmp45209;
  wire tmp45210;
  wire tmp45211;
  wire tmp45212;
  wire tmp45213;
  wire tmp45214;
  wire tmp45215;
  wire tmp45216;
  wire tmp45217;
  wire tmp45218;
  wire tmp45219;
  wire tmp45220;
  wire tmp45221;
  wire tmp45222;
  wire tmp45223;
  wire tmp45224;
  wire tmp45225;
  wire tmp45226;
  wire tmp45227;
  wire tmp45228;
  wire tmp45229;
  wire tmp45230;
  wire tmp45231;
  wire tmp45232;
  wire tmp45233;
  wire tmp45234;
  wire tmp45235;
  wire tmp45236;
  wire tmp45237;
  wire tmp45238;
  wire tmp45239;
  wire tmp45240;
  wire tmp45241;
  wire tmp45242;
  wire tmp45243;
  wire tmp45244;
  wire tmp45245;
  wire tmp45246;
  wire tmp45247;
  wire tmp45248;
  wire tmp45249;
  wire tmp45250;
  wire tmp45251;
  wire tmp45252;
  wire tmp45253;
  wire tmp45254;
  wire tmp45255;
  wire tmp45256;
  wire tmp45257;
  wire tmp45258;
  wire tmp45259;
  wire tmp45260;
  wire tmp45261;
  wire tmp45262;
  wire tmp45263;
  wire tmp45264;
  wire tmp45265;
  wire tmp45266;
  wire tmp45267;
  wire tmp45268;
  wire tmp45269;
  wire tmp45270;
  wire tmp45271;
  wire tmp45272;
  wire tmp45273;
  wire tmp45274;
  wire tmp45275;
  wire tmp45276;
  wire tmp45277;
  wire tmp45278;
  wire tmp45279;
  wire tmp45280;
  wire tmp45281;
  wire tmp45282;
  wire tmp45283;
  wire tmp45284;
  wire tmp45285;
  wire tmp45286;
  wire tmp45287;
  wire tmp45288;
  wire tmp45289;
  wire tmp45290;
  wire tmp45291;
  wire tmp45292;
  wire tmp45293;
  wire tmp45294;
  wire tmp45295;
  wire tmp45296;
  wire tmp45297;
  wire tmp45298;
  wire tmp45299;
  wire tmp45300;
  wire tmp45301;
  wire tmp45302;
  wire tmp45303;
  wire tmp45304;
  wire tmp45305;
  wire tmp45306;
  wire tmp45307;
  wire tmp45308;
  wire tmp45309;
  wire tmp45310;
  wire tmp45311;
  wire tmp45312;
  wire tmp45313;
  wire tmp45314;
  wire tmp45315;
  wire tmp45316;
  wire tmp45317;
  wire tmp45318;
  wire tmp45319;
  wire tmp45320;
  wire tmp45321;
  wire tmp45322;
  wire tmp45323;
  wire tmp45324;
  wire tmp45325;
  wire tmp45326;
  wire tmp45327;
  wire tmp45328;
  wire tmp45329;
  wire tmp45330;
  wire tmp45331;
  wire tmp45332;
  wire tmp45333;
  wire tmp45334;
  wire tmp45335;
  wire tmp45336;
  wire tmp45337;
  wire tmp45338;
  wire tmp45339;
  wire tmp45340;
  wire tmp45341;
  wire tmp45342;
  wire tmp45343;
  wire tmp45344;
  wire tmp45345;
  wire tmp45346;
  wire tmp45347;
  wire tmp45348;
  wire tmp45349;
  wire tmp45350;
  wire tmp45351;
  wire tmp45352;
  wire tmp45353;
  wire tmp45354;
  wire tmp45355;
  wire tmp45356;
  wire tmp45357;
  wire tmp45358;
  wire tmp45359;
  wire tmp45360;
  wire tmp45361;
  wire tmp45362;
  wire tmp45363;
  wire tmp45364;
  wire tmp45365;
  wire tmp45366;
  wire tmp45367;
  wire tmp45368;
  wire tmp45369;
  wire tmp45370;
  wire tmp45371;
  wire tmp45372;
  wire tmp45373;
  wire tmp45374;
  wire tmp45375;
  wire tmp45376;
  wire tmp45377;
  wire tmp45378;
  wire tmp45379;
  wire tmp45380;
  wire tmp45381;
  wire tmp45382;
  wire tmp45383;
  wire tmp45384;
  wire tmp45385;
  wire tmp45386;
  wire tmp45387;
  wire tmp45388;
  wire tmp45389;
  wire tmp45390;
  wire tmp45391;
  wire tmp45392;
  wire tmp45393;
  wire tmp45394;
  wire tmp45395;
  wire tmp45396;
  wire tmp45397;
  wire tmp45398;
  wire tmp45399;
  wire tmp45400;
  wire tmp45401;
  wire tmp45402;
  wire tmp45403;
  wire tmp45404;
  wire tmp45405;
  wire tmp45406;
  wire tmp45407;
  wire tmp45408;
  wire tmp45409;
  wire tmp45410;
  wire tmp45411;
  wire tmp45412;
  wire tmp45413;
  wire tmp45414;
  wire tmp45415;
  wire tmp45416;
  wire tmp45417;
  wire tmp45418;
  wire tmp45419;
  wire tmp45420;
  wire tmp45421;
  wire tmp45422;
  wire tmp45423;
  wire tmp45424;
  wire tmp45425;
  wire tmp45426;
  wire tmp45427;
  wire tmp45428;
  wire tmp45429;
  wire tmp45430;
  wire tmp45431;
  wire tmp45432;
  wire tmp45433;
  wire tmp45434;
  wire tmp45435;
  wire tmp45436;
  wire tmp45437;
  wire tmp45438;
  wire tmp45439;
  wire tmp45440;
  wire tmp45441;
  wire tmp45442;
  wire tmp45443;
  wire tmp45444;
  wire tmp45445;
  wire tmp45446;
  wire tmp45447;
  wire tmp45448;
  wire tmp45449;
  wire tmp45450;
  wire tmp45451;
  wire tmp45452;
  wire tmp45453;
  wire tmp45454;
  wire tmp45455;
  wire tmp45456;
  wire tmp45457;
  wire tmp45458;
  wire tmp45459;
  wire tmp45460;
  wire tmp45461;
  wire tmp45462;
  wire tmp45463;
  wire tmp45464;
  wire tmp45465;
  wire tmp45466;
  wire tmp45467;
  wire tmp45468;
  wire tmp45469;
  wire tmp45470;
  wire tmp45471;
  wire tmp45472;
  wire tmp45473;
  wire tmp45474;
  wire tmp45475;
  wire tmp45476;
  wire tmp45477;
  wire tmp45478;
  wire tmp45479;
  wire tmp45480;
  wire tmp45481;
  wire tmp45482;
  wire tmp45483;
  wire tmp45484;
  wire tmp45485;
  wire tmp45486;
  wire tmp45487;
  wire tmp45488;
  wire tmp45489;
  wire tmp45490;
  wire tmp45491;
  wire tmp45492;
  wire tmp45493;
  wire tmp45494;
  wire tmp45495;
  wire tmp45496;
  wire tmp45497;
  wire tmp45498;
  wire tmp45499;
  wire tmp45500;
  wire tmp45501;
  wire tmp45502;
  wire tmp45503;
  wire tmp45504;
  wire tmp45505;
  wire tmp45506;
  wire tmp45507;
  wire tmp45508;
  wire tmp45509;
  wire tmp45510;
  wire tmp45511;
  wire tmp45512;
  wire tmp45513;
  wire tmp45514;
  wire tmp45515;
  wire tmp45516;
  wire tmp45517;
  wire tmp45518;
  wire tmp45519;
  wire tmp45520;
  wire tmp45521;
  wire tmp45522;
  wire tmp45523;
  wire tmp45524;
  wire tmp45525;
  wire tmp45526;
  wire tmp45527;
  wire tmp45528;
  wire tmp45529;
  wire tmp45530;
  wire tmp45531;
  wire tmp45532;
  wire tmp45533;
  wire tmp45534;
  wire tmp45535;
  wire tmp45536;
  wire tmp45537;
  wire tmp45538;
  wire tmp45539;
  wire tmp45540;
  wire tmp45541;
  wire tmp45542;
  wire tmp45543;
  wire tmp45544;
  wire tmp45545;
  wire tmp45546;
  wire tmp45547;
  wire tmp45548;
  wire tmp45549;
  wire tmp45550;
  wire tmp45551;
  wire tmp45552;
  wire tmp45553;
  wire tmp45554;
  wire tmp45555;
  wire tmp45556;
  wire tmp45557;
  wire tmp45558;
  wire tmp45559;
  wire tmp45560;
  wire tmp45561;
  wire tmp45562;
  wire tmp45563;
  wire tmp45564;
  wire tmp45565;
  wire tmp45566;
  wire tmp45567;
  wire tmp45568;
  wire tmp45569;
  wire tmp45570;
  wire tmp45571;
  wire tmp45572;
  wire tmp45573;
  wire tmp45574;
  wire tmp45575;
  wire tmp45576;
  wire tmp45577;
  wire tmp45578;
  wire tmp45579;
  wire tmp45580;
  wire tmp45581;
  wire tmp45582;
  wire tmp45583;
  wire tmp45584;
  wire tmp45585;
  wire tmp45586;
  wire tmp45587;
  wire tmp45588;
  wire tmp45589;
  wire tmp45590;
  wire tmp45591;
  wire tmp45592;
  wire tmp45593;
  wire tmp45594;
  wire tmp45595;
  wire tmp45596;
  wire tmp45597;
  wire tmp45598;
  wire tmp45599;
  wire tmp45600;
  wire tmp45601;
  wire tmp45602;
  wire tmp45603;
  wire tmp45604;
  wire tmp45605;
  wire tmp45606;
  wire tmp45607;
  wire tmp45608;
  wire tmp45609;
  wire tmp45610;
  wire tmp45611;
  wire tmp45612;
  wire tmp45613;
  wire tmp45614;
  wire tmp45615;
  wire tmp45616;
  wire tmp45617;
  wire tmp45618;
  wire tmp45619;
  wire tmp45620;
  wire tmp45621;
  wire tmp45622;
  wire tmp45623;
  wire tmp45624;
  wire tmp45625;
  wire tmp45626;
  wire tmp45627;
  wire tmp45628;
  wire tmp45629;
  wire tmp45630;
  wire tmp45631;
  wire tmp45632;
  wire tmp45633;
  wire tmp45634;
  wire tmp45635;
  wire tmp45636;
  wire tmp45637;
  wire tmp45638;
  wire tmp45639;
  wire tmp45640;
  wire tmp45641;
  wire tmp45642;
  wire tmp45643;
  wire tmp45644;
  wire tmp45645;
  wire tmp45646;
  wire tmp45647;
  wire tmp45648;
  wire tmp45649;
  wire tmp45650;
  wire tmp45651;
  wire tmp45652;
  wire tmp45653;
  wire tmp45654;
  wire tmp45655;
  wire tmp45656;
  wire tmp45657;
  wire tmp45658;
  wire tmp45659;
  wire tmp45660;
  wire tmp45661;
  wire tmp45662;
  wire tmp45663;
  wire tmp45664;
  wire tmp45665;
  wire tmp45666;
  wire tmp45667;
  wire tmp45668;
  wire tmp45669;
  wire tmp45670;
  wire tmp45671;
  wire tmp45672;
  wire tmp45673;
  wire tmp45674;
  wire tmp45675;
  wire tmp45676;
  wire tmp45677;
  wire tmp45678;
  wire tmp45679;
  wire tmp45680;
  wire tmp45681;
  wire tmp45682;
  wire tmp45683;
  wire tmp45684;
  wire tmp45685;
  wire tmp45686;
  wire tmp45687;
  wire tmp45688;
  wire tmp45689;
  wire tmp45690;
  wire tmp45691;
  wire tmp45692;
  wire tmp45693;
  wire tmp45694;
  wire tmp45695;
  wire tmp45696;
  wire tmp45697;
  wire tmp45698;
  wire tmp45699;
  wire tmp45700;
  wire tmp45701;
  wire tmp45702;
  wire tmp45703;
  wire tmp45704;
  wire tmp45705;
  wire tmp45706;
  wire tmp45707;
  wire tmp45708;
  wire tmp45709;
  wire tmp45710;
  wire tmp45711;
  wire tmp45712;
  wire tmp45713;
  wire tmp45714;
  wire tmp45715;
  wire tmp45716;
  wire tmp45717;
  wire tmp45718;
  wire tmp45719;
  wire tmp45720;
  wire tmp45721;
  wire tmp45722;
  wire tmp45723;
  wire tmp45724;
  wire tmp45725;
  wire tmp45726;
  wire tmp45727;
  wire tmp45728;
  wire tmp45729;
  wire tmp45730;
  wire tmp45731;
  wire tmp45732;
  wire tmp45733;
  wire tmp45734;
  wire tmp45735;
  wire tmp45736;
  wire tmp45737;
  wire tmp45738;
  wire tmp45739;
  wire tmp45740;
  wire tmp45741;
  wire tmp45742;
  wire tmp45743;
  wire tmp45744;
  wire tmp45745;
  wire tmp45746;
  wire tmp45747;
  wire tmp45748;
  wire tmp45749;
  wire tmp45750;
  wire tmp45751;
  wire tmp45752;
  wire tmp45753;
  wire tmp45754;
  wire tmp45755;
  wire tmp45756;
  wire tmp45757;
  wire tmp45758;
  wire tmp45759;
  wire tmp45760;
  wire tmp45761;
  wire tmp45762;
  wire tmp45763;
  wire tmp45764;
  wire tmp45765;
  wire tmp45766;
  wire tmp45767;
  wire tmp45768;
  wire tmp45769;
  wire tmp45770;
  wire tmp45771;
  wire tmp45772;
  wire tmp45773;
  wire tmp45774;
  wire tmp45775;
  wire tmp45776;
  wire tmp45777;
  wire tmp45778;
  wire tmp45779;
  wire tmp45780;
  wire tmp45781;
  wire tmp45782;
  wire tmp45783;
  wire tmp45784;
  wire tmp45785;
  wire tmp45786;
  wire tmp45787;
  wire tmp45788;
  wire tmp45789;
  wire tmp45790;
  wire tmp45791;
  wire tmp45792;
  wire tmp45793;
  wire tmp45794;
  wire tmp45795;
  wire tmp45796;
  wire tmp45797;
  wire tmp45798;
  wire tmp45799;
  wire tmp45800;
  wire tmp45801;
  wire tmp45802;
  wire tmp45803;
  wire tmp45804;
  wire tmp45805;
  wire tmp45806;
  wire tmp45807;
  wire tmp45808;
  wire tmp45809;
  wire tmp45810;
  wire tmp45811;
  wire tmp45812;
  wire tmp45813;
  wire tmp45814;
  wire tmp45815;
  wire tmp45816;
  wire tmp45817;
  wire tmp45818;
  wire tmp45819;
  wire tmp45820;
  wire tmp45821;
  wire tmp45822;
  wire tmp45823;
  wire tmp45824;
  wire tmp45825;
  wire tmp45826;
  wire tmp45827;
  wire tmp45828;
  wire tmp45829;
  wire tmp45830;
  wire tmp45831;
  wire tmp45832;
  wire tmp45833;
  wire tmp45834;
  wire tmp45835;
  wire tmp45836;
  wire tmp45837;
  wire tmp45838;
  wire tmp45839;
  wire tmp45840;
  wire tmp45841;
  wire tmp45842;
  wire tmp45843;
  wire tmp45844;
  wire tmp45845;
  wire tmp45846;
  wire tmp45847;
  wire tmp45848;
  wire tmp45849;
  wire tmp45850;
  wire tmp45851;
  wire tmp45852;
  wire tmp45853;
  wire tmp45854;
  wire tmp45855;
  wire tmp45856;
  wire tmp45857;
  wire tmp45858;
  wire tmp45859;
  wire tmp45860;
  wire tmp45861;
  wire tmp45862;
  wire tmp45863;
  wire tmp45864;
  wire tmp45865;
  wire tmp45866;
  wire tmp45867;
  wire tmp45868;
  wire tmp45869;
  wire tmp45870;
  wire tmp45871;
  wire tmp45872;
  wire tmp45873;
  wire tmp45874;
  wire tmp45875;
  wire tmp45876;
  wire tmp45877;
  wire tmp45878;
  wire tmp45879;
  wire tmp45880;
  wire tmp45881;
  wire tmp45882;
  wire tmp45883;
  wire tmp45884;
  wire tmp45885;
  wire tmp45886;
  wire tmp45887;
  wire tmp45888;
  wire tmp45889;
  wire tmp45890;
  wire tmp45891;
  wire tmp45892;
  wire tmp45893;
  wire tmp45894;
  wire tmp45895;
  wire tmp45896;
  wire tmp45897;
  wire tmp45898;
  wire tmp45899;
  wire tmp45900;
  wire tmp45901;
  wire tmp45902;
  wire tmp45903;
  wire tmp45904;
  wire tmp45905;
  wire tmp45906;
  wire tmp45907;
  wire tmp45908;
  wire tmp45909;
  wire tmp45910;
  wire tmp45911;
  wire tmp45912;
  wire tmp45913;
  wire tmp45914;
  wire tmp45915;
  wire tmp45916;
  wire tmp45917;
  wire tmp45918;
  wire tmp45919;
  wire tmp45920;
  wire tmp45921;
  wire tmp45922;
  wire tmp45923;
  wire tmp45924;
  wire tmp45925;
  wire tmp45926;
  wire tmp45927;
  wire tmp45928;
  wire tmp45929;
  wire tmp45930;
  wire tmp45931;
  wire tmp45932;
  wire tmp45933;
  wire tmp45934;
  wire tmp45935;
  wire tmp45936;
  wire tmp45937;
  wire tmp45938;
  wire tmp45939;
  wire tmp45940;
  wire tmp45941;
  wire tmp45942;
  wire tmp45943;
  wire tmp45944;
  wire tmp45945;
  wire tmp45946;
  wire tmp45947;
  wire tmp45948;
  wire tmp45949;
  wire tmp45950;
  wire tmp45951;
  wire tmp45952;
  wire tmp45953;
  wire tmp45954;
  wire tmp45955;
  wire tmp45956;
  wire tmp45957;
  wire tmp45958;
  wire tmp45959;
  wire tmp45960;
  wire tmp45961;
  wire tmp45962;
  wire tmp45963;
  wire tmp45964;
  wire tmp45965;
  wire tmp45966;
  wire tmp45967;
  wire tmp45968;
  wire tmp45969;
  wire tmp45970;
  wire tmp45971;
  wire tmp45972;
  wire tmp45973;
  wire tmp45974;
  wire tmp45975;
  wire tmp45976;
  wire tmp45977;
  wire tmp45978;
  wire tmp45979;
  wire tmp45980;
  wire tmp45981;
  wire tmp45982;
  wire tmp45983;
  wire tmp45984;
  wire tmp45985;
  wire tmp45986;
  wire tmp45987;
  wire tmp45988;
  wire tmp45989;
  wire tmp45990;
  wire tmp45991;
  wire tmp45992;
  wire tmp45993;
  wire tmp45994;
  wire tmp45995;
  wire tmp45996;
  wire tmp45997;
  wire tmp45998;
  wire tmp45999;
  wire tmp46000;
  wire tmp46001;
  wire tmp46002;
  wire tmp46003;
  wire tmp46004;
  wire tmp46005;
  wire tmp46006;
  wire tmp46007;
  wire tmp46008;
  wire tmp46009;
  wire tmp46010;
  wire tmp46011;
  wire tmp46012;
  wire tmp46013;
  wire tmp46014;
  wire tmp46015;
  wire tmp46016;
  wire tmp46017;
  wire tmp46018;
  wire tmp46019;
  wire tmp46020;
  wire tmp46021;
  wire tmp46022;
  wire tmp46023;
  wire tmp46024;
  wire tmp46025;
  wire tmp46026;
  wire tmp46027;
  wire tmp46028;
  wire tmp46029;
  wire tmp46030;
  wire tmp46031;
  wire tmp46032;
  wire tmp46033;
  wire tmp46034;
  wire tmp46035;
  wire tmp46036;
  wire tmp46037;
  wire tmp46038;
  wire tmp46039;
  wire tmp46040;
  wire tmp46041;
  wire tmp46042;
  wire tmp46043;
  wire tmp46044;
  wire tmp46045;
  wire tmp46046;
  wire tmp46047;
  wire tmp46048;
  wire tmp46049;
  wire tmp46050;
  wire tmp46051;
  wire tmp46052;
  wire tmp46053;
  wire tmp46054;
  wire tmp46055;
  wire tmp46056;
  wire tmp46057;
  wire tmp46058;
  wire tmp46059;
  wire tmp46060;
  wire tmp46061;
  wire tmp46062;
  wire tmp46063;
  wire tmp46064;
  wire tmp46065;
  wire tmp46066;
  wire tmp46067;
  wire tmp46068;
  wire tmp46069;
  wire tmp46070;
  wire tmp46071;
  wire tmp46072;
  wire tmp46073;
  wire tmp46074;
  wire tmp46075;
  wire tmp46076;
  wire tmp46077;
  wire tmp46078;
  wire tmp46079;
  wire tmp46080;
  wire tmp46081;
  wire tmp46082;
  wire tmp46083;
  wire tmp46084;
  wire tmp46085;
  wire tmp46086;
  wire tmp46087;
  wire tmp46088;
  wire tmp46089;
  wire tmp46090;
  wire tmp46091;
  wire tmp46092;
  wire tmp46093;
  wire tmp46094;
  wire tmp46095;
  wire tmp46096;
  wire tmp46097;
  wire tmp46098;
  wire tmp46099;
  wire tmp46100;
  wire tmp46101;
  wire tmp46102;
  wire tmp46103;
  wire tmp46104;
  wire tmp46105;
  wire tmp46106;
  wire tmp46107;
  wire tmp46108;
  wire tmp46109;
  wire tmp46110;
  wire tmp46111;
  wire tmp46112;
  wire tmp46113;
  wire tmp46114;
  wire tmp46115;
  wire tmp46116;
  wire tmp46117;
  wire tmp46118;
  wire tmp46119;
  wire tmp46120;
  wire tmp46121;
  wire tmp46122;
  wire tmp46123;
  wire tmp46124;
  wire tmp46125;
  wire tmp46126;
  wire tmp46127;
  wire tmp46128;
  wire tmp46129;
  wire tmp46130;
  wire tmp46131;
  wire tmp46132;
  wire tmp46133;
  wire tmp46134;
  wire tmp46135;
  wire tmp46136;
  wire tmp46137;
  wire tmp46138;
  wire tmp46139;
  wire tmp46140;
  wire tmp46141;
  wire tmp46142;
  wire tmp46143;
  wire tmp46144;
  wire tmp46145;
  wire tmp46146;
  wire tmp46147;
  wire tmp46148;
  wire tmp46149;
  wire tmp46150;
  wire tmp46151;
  wire tmp46152;
  wire tmp46153;
  wire tmp46154;
  wire tmp46155;
  wire tmp46156;
  wire tmp46157;
  wire tmp46158;
  wire tmp46159;
  wire tmp46160;
  wire tmp46161;
  wire tmp46162;
  wire tmp46163;
  wire tmp46164;
  wire tmp46165;
  wire tmp46166;
  wire tmp46167;
  wire tmp46168;
  wire tmp46169;
  wire tmp46170;
  wire tmp46171;
  wire tmp46172;
  wire tmp46173;
  wire tmp46174;
  wire tmp46175;

  reg s0;
  reg s1;
  reg s2;
  reg s3;
  reg s4;
  reg s5;
  reg s6;
  reg s7;
  reg s8;
  reg s9;
  reg s10;
  reg s11;
  reg s12;
  reg s13;
  reg s14;
  reg s15;
  reg s16;
  reg s17;
  reg s18;

  assign tmp17 = l4 ? 1 : 0;
  assign tmp16 = ~(l3 ? tmp17 : 1);
  assign tmp15 = l2 ? 1 : tmp16;
  assign tmp19 = l3 ? 1 : 0;
  assign tmp21 = ~(l4 ? 1 : 0);
  assign tmp20 = ~(l3 ? 1 : tmp21);
  assign tmp18 = ~(l2 ? tmp19 : tmp20);
  assign tmp14 = l1 ? tmp15 : tmp18;
  assign tmp24 = l2 ? tmp19 : 0;
  assign tmp23 = l1 ? 1 : tmp24;
  assign tmp26 = l2 ? 1 : tmp21;
  assign tmp25 = ~(l1 ? tmp26 : tmp18);
  assign tmp22 = ~(s0 ? tmp23 : tmp25);
  assign tmp13 = s1 ? tmp14 : tmp22;
  assign tmp31 = l2 ? 1 : 0;
  assign tmp33 = ~(l3 ? 1 : 0);
  assign tmp32 = ~(l2 ? 1 : tmp33);
  assign tmp30 = l1 ? tmp31 : tmp32;
  assign tmp35 = l2 ? tmp17 : tmp20;
  assign tmp34 = ~(l1 ? tmp17 : tmp35);
  assign tmp29 = s0 ? tmp30 : tmp34;
  assign tmp38 = ~(l2 ? tmp19 : tmp33);
  assign tmp37 = l1 ? tmp15 : tmp38;
  assign tmp36 = s0 ? tmp37 : tmp34;
  assign tmp28 = s1 ? tmp29 : tmp36;
  assign tmp41 = ~(l1 ? 1 : tmp31);
  assign tmp40 = s0 ? tmp37 : tmp41;
  assign tmp43 = l1 ? tmp17 : tmp35;
  assign tmp45 = l2 ? tmp19 : tmp20;
  assign tmp44 = l1 ? tmp17 : tmp45;
  assign tmp42 = ~(s0 ? tmp43 : tmp44);
  assign tmp39 = s1 ? tmp40 : tmp42;
  assign tmp27 = s2 ? tmp28 : tmp39;
  assign tmp12 = s3 ? tmp13 : tmp27;
  assign tmp50 = l1 ? tmp31 : tmp18;
  assign tmp49 = s0 ? tmp50 : tmp41;
  assign tmp51 = ~(s0 ? tmp44 : tmp43);
  assign tmp48 = s1 ? tmp49 : tmp51;
  assign tmp54 = ~(l1 ? 1 : 0);
  assign tmp53 = s0 ? tmp14 : tmp54;
  assign tmp55 = ~(l1 ? 1 : tmp19);
  assign tmp52 = s1 ? tmp53 : tmp55;
  assign tmp47 = s2 ? tmp48 : tmp52;
  assign tmp57 = s1 ? tmp23 : 0;
  assign tmp59 = ~(s0 ? 1 : tmp34);
  assign tmp58 = s1 ? tmp43 : tmp59;
  assign tmp56 = ~(s2 ? tmp57 : tmp58);
  assign tmp46 = s3 ? tmp47 : tmp56;
  assign tmp11 = s4 ? tmp12 : tmp46;
  assign tmp66 = l1 ? tmp26 : tmp18;
  assign tmp65 = s0 ? tmp66 : tmp41;
  assign tmp64 = s1 ? tmp65 : tmp30;
  assign tmp69 = ~(l3 ? 1 : tmp17);
  assign tmp68 = l1 ? tmp26 : tmp69;
  assign tmp70 = ~(s0 ? tmp43 : tmp31);
  assign tmp67 = s1 ? tmp68 : tmp70;
  assign tmp63 = s2 ? tmp64 : tmp67;
  assign tmp74 = l2 ? 1 : tmp19;
  assign tmp73 = l1 ? tmp74 : tmp38;
  assign tmp72 = s1 ? tmp73 : tmp21;
  assign tmp75 = s1 ? 1 : tmp21;
  assign tmp71 = s2 ? tmp72 : tmp75;
  assign tmp62 = s3 ? tmp63 : tmp71;
  assign tmp81 = l2 ? tmp19 : tmp17;
  assign tmp80 = ~(l1 ? tmp17 : tmp81);
  assign tmp79 = s0 ? 1 : tmp80;
  assign tmp83 = l1 ? 1 : 0;
  assign tmp82 = ~(s0 ? 1 : tmp83);
  assign tmp78 = s1 ? tmp79 : tmp82;
  assign tmp84 = l1 ? tmp31 : tmp69;
  assign tmp77 = s2 ? tmp78 : tmp84;
  assign tmp88 = l1 ? tmp74 : tmp26;
  assign tmp87 = s0 ? tmp84 : tmp88;
  assign tmp86 = s1 ? tmp87 : tmp21;
  assign tmp85 = s2 ? tmp86 : 1;
  assign tmp76 = s3 ? tmp77 : tmp85;
  assign tmp61 = s4 ? tmp62 : tmp76;
  assign tmp93 = s0 ? tmp17 : 0;
  assign tmp92 = s1 ? tmp93 : 0;
  assign tmp94 = ~(l1 ? tmp31 : 0);
  assign tmp91 = s2 ? tmp92 : tmp94;
  assign tmp97 = l1 ? tmp31 : tmp21;
  assign tmp96 = s1 ? 1 : tmp97;
  assign tmp95 = ~(s2 ? 1 : tmp96);
  assign tmp90 = s3 ? tmp91 : tmp95;
  assign tmp99 = s2 ? 1 : tmp68;
  assign tmp102 = ~(l2 ? 1 : tmp21);
  assign tmp101 = ~(l1 ? tmp17 : tmp102);
  assign tmp100 = s1 ? 1 : tmp101;
  assign tmp98 = ~(s3 ? tmp99 : tmp100);
  assign tmp89 = ~(s4 ? tmp90 : tmp98);
  assign tmp60 = s5 ? tmp61 : tmp89;
  assign tmp10 = ~(s6 ? tmp11 : tmp60);
  assign tmp9 = s7 ? 1 : tmp10;
  assign tmp110 = l3 ? tmp17 : 1;
  assign tmp109 = l2 ? tmp17 : tmp110;
  assign tmp108 = l1 ? tmp109 : tmp45;
  assign tmp111 = s0 ? tmp23 : tmp44;
  assign tmp107 = s1 ? tmp108 : tmp111;
  assign tmp116 = l2 ? tmp17 : 1;
  assign tmp117 = l2 ? tmp19 : tmp33;
  assign tmp115 = l1 ? tmp116 : tmp117;
  assign tmp120 = l3 ? tmp17 : 0;
  assign tmp119 = l2 ? tmp120 : tmp20;
  assign tmp118 = l1 ? tmp17 : tmp119;
  assign tmp114 = s0 ? tmp115 : tmp118;
  assign tmp122 = l1 ? tmp109 : tmp117;
  assign tmp121 = s0 ? tmp122 : tmp118;
  assign tmp113 = s1 ? tmp114 : tmp121;
  assign tmp124 = s0 ? tmp122 : tmp23;
  assign tmp125 = s0 ? tmp118 : tmp44;
  assign tmp123 = s1 ? tmp124 : tmp125;
  assign tmp112 = s2 ? tmp113 : tmp123;
  assign tmp106 = s3 ? tmp107 : tmp112;
  assign tmp130 = l1 ? tmp116 : tmp45;
  assign tmp131 = l1 ? 1 : tmp31;
  assign tmp129 = s0 ? tmp130 : tmp131;
  assign tmp132 = s0 ? tmp44 : tmp118;
  assign tmp128 = s1 ? tmp129 : tmp132;
  assign tmp134 = s0 ? tmp108 : tmp83;
  assign tmp135 = l1 ? 1 : tmp19;
  assign tmp133 = s1 ? tmp134 : tmp135;
  assign tmp127 = s2 ? tmp128 : tmp133;
  assign tmp139 = ~(l1 ? tmp17 : tmp119);
  assign tmp138 = ~(s0 ? 1 : tmp139);
  assign tmp137 = s1 ? tmp118 : tmp138;
  assign tmp136 = s2 ? tmp57 : tmp137;
  assign tmp126 = s3 ? tmp127 : tmp136;
  assign tmp105 = s4 ? tmp106 : tmp126;
  assign tmp145 = s0 ? tmp44 : tmp131;
  assign tmp144 = s1 ? tmp145 : tmp115;
  assign tmp147 = l1 ? tmp17 : tmp81;
  assign tmp148 = s0 ? tmp118 : tmp23;
  assign tmp146 = s1 ? tmp147 : tmp148;
  assign tmp143 = s2 ? tmp144 : tmp146;
  assign tmp152 = l2 ? tmp17 : tmp33;
  assign tmp151 = l1 ? tmp152 : tmp117;
  assign tmp154 = l2 ? tmp120 : tmp17;
  assign tmp153 = l1 ? tmp17 : tmp154;
  assign tmp150 = s1 ? tmp151 : tmp153;
  assign tmp156 = ~(l1 ? tmp17 : tmp154);
  assign tmp155 = ~(s1 ? 1 : tmp156);
  assign tmp149 = s2 ? tmp150 : tmp155;
  assign tmp142 = s3 ? tmp143 : tmp149;
  assign tmp159 = ~(l1 ? tmp116 : tmp81);
  assign tmp158 = s2 ? tmp78 : tmp159;
  assign tmp164 = ~(l2 ? tmp19 : tmp17);
  assign tmp163 = l1 ? tmp31 : tmp164;
  assign tmp165 = ~(l1 ? tmp152 : tmp102);
  assign tmp162 = s0 ? tmp163 : tmp165;
  assign tmp161 = s1 ? tmp162 : tmp21;
  assign tmp160 = s2 ? tmp161 : 1;
  assign tmp157 = ~(s3 ? tmp158 : tmp160);
  assign tmp141 = s4 ? tmp142 : tmp157;
  assign tmp170 = s0 ? tmp153 : 0;
  assign tmp169 = s1 ? tmp170 : 0;
  assign tmp173 = ~(l2 ? tmp19 : 1);
  assign tmp172 = l1 ? tmp31 : tmp173;
  assign tmp174 = l1 ? tmp31 : 0;
  assign tmp171 = ~(s1 ? tmp172 : tmp174);
  assign tmp168 = s2 ? tmp169 : tmp171;
  assign tmp167 = s3 ? tmp168 : tmp95;
  assign tmp177 = l1 ? tmp26 : tmp164;
  assign tmp176 = s2 ? 1 : tmp177;
  assign tmp175 = ~(s3 ? tmp176 : tmp100);
  assign tmp166 = s4 ? tmp167 : tmp175;
  assign tmp140 = s5 ? tmp141 : tmp166;
  assign tmp104 = s6 ? tmp105 : tmp140;
  assign tmp103 = s7 ? 1 : tmp104;
  assign tmp8 = s8 ? tmp9 : tmp103;
  assign tmp185 = ~(l2 ? tmp19 : 0);
  assign tmp184 = l1 ? tmp15 : tmp185;
  assign tmp187 = l1 ? tmp31 : tmp185;
  assign tmp188 = l1 ? tmp26 : tmp185;
  assign tmp186 = s0 ? tmp187 : tmp188;
  assign tmp183 = s1 ? tmp184 : tmp186;
  assign tmp193 = ~(l2 ? tmp120 : 0);
  assign tmp192 = l1 ? tmp26 : tmp193;
  assign tmp191 = s0 ? tmp187 : tmp192;
  assign tmp194 = s0 ? tmp184 : tmp192;
  assign tmp190 = s1 ? tmp191 : tmp194;
  assign tmp196 = s0 ? tmp184 : tmp187;
  assign tmp197 = s0 ? tmp192 : tmp188;
  assign tmp195 = s1 ? tmp196 : tmp197;
  assign tmp189 = s2 ? tmp190 : tmp195;
  assign tmp182 = s3 ? tmp183 : tmp189;
  assign tmp203 = ~(l2 ? 1 : 0);
  assign tmp202 = l1 ? tmp31 : tmp203;
  assign tmp201 = s0 ? tmp187 : tmp202;
  assign tmp204 = s0 ? tmp188 : tmp192;
  assign tmp200 = s1 ? tmp201 : tmp204;
  assign tmp207 = l1 ? tmp31 : 1;
  assign tmp206 = s0 ? tmp184 : tmp207;
  assign tmp208 = l1 ? tmp31 : tmp33;
  assign tmp205 = s1 ? tmp206 : tmp208;
  assign tmp199 = s2 ? tmp200 : tmp205;
  assign tmp210 = s1 ? tmp187 : 1;
  assign tmp212 = s0 ? 1 : tmp192;
  assign tmp211 = s1 ? tmp192 : tmp212;
  assign tmp209 = s2 ? tmp210 : tmp211;
  assign tmp198 = s3 ? tmp199 : tmp209;
  assign tmp181 = s4 ? tmp182 : tmp198;
  assign tmp218 = s0 ? tmp188 : tmp41;
  assign tmp217 = s1 ? tmp218 : tmp187;
  assign tmp221 = l1 ? 1 : tmp185;
  assign tmp220 = s0 ? tmp192 : tmp221;
  assign tmp219 = s1 ? tmp188 : tmp220;
  assign tmp216 = s2 ? tmp217 : tmp219;
  assign tmp224 = l1 ? tmp74 : tmp185;
  assign tmp226 = l2 ? tmp120 : 0;
  assign tmp225 = ~(l1 ? tmp17 : tmp226);
  assign tmp223 = s1 ? tmp224 : tmp225;
  assign tmp228 = ~(l2 ? tmp120 : tmp17);
  assign tmp227 = s1 ? 1 : tmp228;
  assign tmp222 = s2 ? tmp223 : tmp227;
  assign tmp215 = s3 ? tmp216 : tmp222;
  assign tmp232 = s0 ? 1 : tmp188;
  assign tmp233 = s0 ? tmp174 : tmp207;
  assign tmp231 = s1 ? tmp232 : tmp233;
  assign tmp230 = s2 ? tmp231 : tmp187;
  assign tmp237 = l1 ? tmp74 : 1;
  assign tmp236 = s0 ? tmp187 : tmp237;
  assign tmp235 = s1 ? tmp236 : tmp21;
  assign tmp234 = s2 ? tmp235 : 1;
  assign tmp229 = s3 ? tmp230 : tmp234;
  assign tmp214 = s4 ? tmp215 : tmp229;
  assign tmp243 = l1 ? tmp17 : tmp226;
  assign tmp242 = s0 ? tmp243 : 0;
  assign tmp241 = s1 ? tmp242 : 0;
  assign tmp244 = ~(s1 ? tmp208 : tmp31);
  assign tmp240 = s2 ? tmp241 : tmp244;
  assign tmp246 = s1 ? 1 : tmp207;
  assign tmp245 = ~(s2 ? 1 : tmp246);
  assign tmp239 = s3 ? tmp240 : tmp245;
  assign tmp248 = s2 ? 1 : tmp188;
  assign tmp250 = ~(l1 ? tmp17 : 0);
  assign tmp249 = s1 ? 1 : tmp250;
  assign tmp247 = ~(s3 ? tmp248 : tmp249);
  assign tmp238 = ~(s4 ? tmp239 : tmp247);
  assign tmp213 = s5 ? tmp214 : tmp238;
  assign tmp180 = ~(s6 ? tmp181 : tmp213);
  assign tmp179 = s7 ? 1 : tmp180;
  assign tmp178 = s8 ? tmp103 : tmp179;
  assign tmp7 = s9 ? tmp8 : tmp178;
  assign tmp258 = s0 ? tmp187 : tmp66;
  assign tmp257 = s1 ? tmp14 : tmp258;
  assign tmp262 = l1 ? tmp31 : tmp38;
  assign tmp264 = ~(l2 ? tmp120 : tmp20);
  assign tmp263 = l1 ? tmp26 : tmp264;
  assign tmp261 = s0 ? tmp262 : tmp263;
  assign tmp265 = s0 ? tmp37 : tmp263;
  assign tmp260 = s1 ? tmp261 : tmp265;
  assign tmp267 = s0 ? tmp37 : tmp187;
  assign tmp268 = s0 ? tmp263 : tmp66;
  assign tmp266 = s1 ? tmp267 : tmp268;
  assign tmp259 = s2 ? tmp260 : tmp266;
  assign tmp256 = s3 ? tmp257 : tmp259;
  assign tmp272 = s0 ? tmp50 : tmp202;
  assign tmp273 = s0 ? tmp66 : tmp263;
  assign tmp271 = s1 ? tmp272 : tmp273;
  assign tmp275 = s0 ? tmp14 : tmp207;
  assign tmp274 = s1 ? tmp275 : tmp208;
  assign tmp270 = s2 ? tmp271 : tmp274;
  assign tmp278 = s0 ? 1 : tmp263;
  assign tmp277 = s1 ? tmp263 : tmp278;
  assign tmp276 = s2 ? tmp210 : tmp277;
  assign tmp269 = s3 ? tmp270 : tmp276;
  assign tmp255 = s4 ? tmp256 : tmp269;
  assign tmp283 = s1 ? tmp65 : tmp262;
  assign tmp285 = s0 ? tmp263 : tmp221;
  assign tmp284 = s1 ? tmp177 : tmp285;
  assign tmp282 = s2 ? tmp283 : tmp284;
  assign tmp287 = s1 ? tmp73 : tmp156;
  assign tmp286 = s2 ? tmp287 : tmp227;
  assign tmp281 = s3 ? tmp282 : tmp286;
  assign tmp291 = s0 ? 1 : tmp177;
  assign tmp290 = s1 ? tmp291 : tmp233;
  assign tmp289 = s2 ? tmp290 : tmp163;
  assign tmp294 = s0 ? tmp163 : tmp88;
  assign tmp293 = s1 ? tmp294 : tmp21;
  assign tmp292 = s2 ? tmp293 : 1;
  assign tmp288 = s3 ? tmp289 : tmp292;
  assign tmp280 = s4 ? tmp281 : tmp288;
  assign tmp295 = ~(s4 ? tmp167 : tmp175);
  assign tmp279 = s5 ? tmp280 : tmp295;
  assign tmp254 = ~(s6 ? tmp255 : tmp279);
  assign tmp253 = s7 ? 1 : tmp254;
  assign tmp252 = s8 ? tmp253 : 1;
  assign tmp298 = s6 ? tmp11 : tmp60;
  assign tmp299 = s6 ? tmp181 : tmp213;
  assign tmp297 = s7 ? tmp298 : tmp299;
  assign tmp300 = ~(s7 ? tmp104 : tmp254);
  assign tmp296 = ~(s8 ? tmp297 : tmp300);
  assign tmp251 = s9 ? tmp252 : tmp296;
  assign tmp6 = s10 ? tmp7 : tmp251;
  assign tmp312 = ~(l3 ? tmp17 : 0);
  assign tmp311 = l2 ? 1 : tmp312;
  assign tmp313 = ~(l2 ? tmp19 : tmp120);
  assign tmp310 = l1 ? tmp311 : tmp313;
  assign tmp316 = l2 ? tmp19 : 1;
  assign tmp315 = l1 ? tmp19 : tmp316;
  assign tmp317 = ~(l1 ? tmp311 : tmp33);
  assign tmp314 = ~(s0 ? tmp315 : tmp317);
  assign tmp309 = s1 ? tmp310 : tmp314;
  assign tmp322 = l2 ? 1 : tmp33;
  assign tmp323 = ~(l2 ? 1 : tmp19);
  assign tmp321 = l1 ? tmp322 : tmp323;
  assign tmp324 = ~(l2 ? tmp17 : tmp120);
  assign tmp320 = s0 ? tmp321 : tmp324;
  assign tmp326 = l1 ? tmp311 : tmp33;
  assign tmp325 = s0 ? tmp326 : tmp324;
  assign tmp319 = s1 ? tmp320 : tmp325;
  assign tmp328 = s0 ? tmp326 : 0;
  assign tmp330 = l2 ? tmp17 : tmp120;
  assign tmp331 = ~(l1 ? tmp311 : tmp313);
  assign tmp329 = ~(s0 ? tmp330 : tmp331);
  assign tmp327 = s1 ? tmp328 : tmp329;
  assign tmp318 = s2 ? tmp319 : tmp327;
  assign tmp308 = s3 ? tmp309 : tmp318;
  assign tmp336 = l1 ? tmp322 : tmp33;
  assign tmp337 = ~(l1 ? tmp19 : 1);
  assign tmp335 = s0 ? tmp336 : tmp337;
  assign tmp338 = s0 ? tmp310 : tmp324;
  assign tmp334 = s1 ? tmp335 : tmp338;
  assign tmp340 = s0 ? tmp310 : 0;
  assign tmp339 = s1 ? tmp340 : tmp33;
  assign tmp333 = s2 ? tmp334 : tmp339;
  assign tmp342 = s1 ? tmp315 : 0;
  assign tmp344 = ~(s0 ? 1 : tmp324);
  assign tmp343 = s1 ? tmp330 : tmp344;
  assign tmp341 = ~(s2 ? tmp342 : tmp343);
  assign tmp332 = s3 ? tmp333 : tmp341;
  assign tmp307 = s4 ? tmp308 : tmp332;
  assign tmp349 = s1 ? tmp328 : tmp321;
  assign tmp351 = l1 ? tmp311 : tmp185;
  assign tmp352 = ~(s0 ? tmp330 : 1);
  assign tmp350 = s1 ? tmp351 : tmp352;
  assign tmp348 = s2 ? tmp349 : tmp350;
  assign tmp355 = l1 ? 1 : tmp33;
  assign tmp356 = ~(l2 ? tmp17 : 0);
  assign tmp354 = s1 ? tmp355 : tmp356;
  assign tmp357 = s1 ? 1 : tmp324;
  assign tmp353 = s2 ? tmp354 : tmp357;
  assign tmp347 = s3 ? tmp348 : tmp353;
  assign tmp361 = s0 ? 1 : tmp351;
  assign tmp363 = l1 ? tmp19 : 1;
  assign tmp362 = ~(s0 ? tmp363 : 0);
  assign tmp360 = s1 ? tmp361 : tmp362;
  assign tmp364 = l1 ? tmp322 : tmp185;
  assign tmp359 = s2 ? tmp360 : tmp364;
  assign tmp367 = s0 ? tmp221 : 1;
  assign tmp366 = s1 ? tmp367 : 1;
  assign tmp365 = s2 ? tmp366 : 1;
  assign tmp358 = s3 ? tmp359 : tmp365;
  assign tmp346 = s4 ? tmp347 : tmp358;
  assign tmp373 = l2 ? tmp17 : 0;
  assign tmp372 = s0 ? tmp373 : 0;
  assign tmp371 = s1 ? tmp372 : 0;
  assign tmp375 = l1 ? 1 : tmp203;
  assign tmp374 = ~(s1 ? tmp375 : 1);
  assign tmp370 = s2 ? tmp371 : tmp374;
  assign tmp369 = s3 ? tmp370 : 0;
  assign tmp377 = s2 ? 1 : tmp221;
  assign tmp376 = ~(s3 ? tmp377 : 1);
  assign tmp368 = ~(s4 ? tmp369 : tmp376);
  assign tmp345 = s5 ? tmp346 : tmp368;
  assign tmp306 = ~(s6 ? tmp307 : tmp345);
  assign tmp305 = s7 ? 1 : tmp306;
  assign tmp384 = l2 ? tmp19 : tmp120;
  assign tmp383 = l1 ? tmp330 : tmp384;
  assign tmp386 = l1 ? tmp74 : tmp316;
  assign tmp387 = l1 ? tmp330 : tmp19;
  assign tmp385 = s0 ? tmp386 : tmp387;
  assign tmp382 = s1 ? tmp383 : tmp385;
  assign tmp392 = l2 ? tmp17 : tmp19;
  assign tmp391 = l1 ? tmp392 : tmp19;
  assign tmp393 = l1 ? tmp330 : tmp120;
  assign tmp390 = s0 ? tmp391 : tmp393;
  assign tmp394 = s0 ? tmp387 : tmp393;
  assign tmp389 = s1 ? tmp390 : tmp394;
  assign tmp397 = l1 ? 1 : tmp316;
  assign tmp396 = s0 ? tmp387 : tmp397;
  assign tmp398 = s0 ? tmp393 : tmp383;
  assign tmp395 = s1 ? tmp396 : tmp398;
  assign tmp388 = s2 ? tmp389 : tmp395;
  assign tmp381 = s3 ? tmp382 : tmp388;
  assign tmp402 = s0 ? tmp391 : tmp237;
  assign tmp403 = s0 ? tmp383 : tmp393;
  assign tmp401 = s1 ? tmp402 : tmp403;
  assign tmp405 = s0 ? tmp383 : 1;
  assign tmp406 = l1 ? tmp74 : tmp19;
  assign tmp404 = s1 ? tmp405 : tmp406;
  assign tmp400 = s2 ? tmp401 : tmp404;
  assign tmp408 = s1 ? tmp386 : 0;
  assign tmp411 = ~(l1 ? tmp330 : tmp120);
  assign tmp410 = ~(s0 ? 1 : tmp411);
  assign tmp409 = s1 ? tmp393 : tmp410;
  assign tmp407 = s2 ? tmp408 : tmp409;
  assign tmp399 = s3 ? tmp400 : tmp407;
  assign tmp380 = s4 ? tmp381 : tmp399;
  assign tmp417 = s0 ? tmp387 : 1;
  assign tmp416 = s1 ? tmp417 : tmp391;
  assign tmp420 = l1 ? tmp373 : tmp120;
  assign tmp419 = s0 ? tmp420 : tmp397;
  assign tmp418 = s1 ? tmp387 : tmp419;
  assign tmp415 = s2 ? tmp416 : tmp418;
  assign tmp423 = l1 ? tmp373 : tmp19;
  assign tmp424 = ~(l1 ? 1 : tmp312);
  assign tmp422 = s1 ? tmp423 : tmp424;
  assign tmp425 = ~(s1 ? 1 : tmp411);
  assign tmp421 = s2 ? tmp422 : tmp425;
  assign tmp414 = s3 ? tmp415 : tmp421;
  assign tmp430 = ~(l1 ? tmp330 : tmp24);
  assign tmp429 = s0 ? 1 : tmp430;
  assign tmp431 = ~(s0 ? tmp237 : tmp174);
  assign tmp428 = s1 ? tmp429 : tmp431;
  assign tmp432 = ~(l1 ? tmp392 : tmp19);
  assign tmp427 = s2 ? tmp428 : tmp432;
  assign tmp436 = ~(l1 ? tmp373 : 0);
  assign tmp435 = s0 ? tmp355 : tmp436;
  assign tmp434 = s1 ? tmp435 : 1;
  assign tmp433 = s2 ? tmp434 : 1;
  assign tmp426 = ~(s3 ? tmp427 : tmp433);
  assign tmp413 = s4 ? tmp414 : tmp426;
  assign tmp442 = l1 ? 1 : tmp312;
  assign tmp441 = s0 ? tmp442 : 1;
  assign tmp440 = s1 ? tmp441 : 1;
  assign tmp443 = s1 ? tmp355 : 1;
  assign tmp439 = s2 ? tmp440 : tmp443;
  assign tmp438 = s3 ? tmp439 : 1;
  assign tmp445 = s2 ? 1 : tmp355;
  assign tmp444 = s3 ? tmp445 : 1;
  assign tmp437 = ~(s4 ? tmp438 : tmp444);
  assign tmp412 = s5 ? tmp413 : tmp437;
  assign tmp379 = s6 ? tmp380 : tmp412;
  assign tmp378 = s7 ? 1 : tmp379;
  assign tmp304 = s8 ? tmp305 : tmp378;
  assign tmp452 = l1 ? tmp311 : tmp164;
  assign tmp451 = s1 ? tmp452 : tmp314;
  assign tmp456 = l1 ? tmp322 : tmp173;
  assign tmp457 = ~(l1 ? tmp120 : tmp154);
  assign tmp455 = s0 ? tmp456 : tmp457;
  assign tmp459 = l1 ? tmp311 : tmp173;
  assign tmp458 = s0 ? tmp459 : tmp457;
  assign tmp454 = s1 ? tmp455 : tmp458;
  assign tmp461 = s0 ? tmp459 : tmp173;
  assign tmp463 = l1 ? tmp120 : tmp154;
  assign tmp464 = l1 ? tmp120 : tmp81;
  assign tmp462 = ~(s0 ? tmp463 : tmp464);
  assign tmp460 = s1 ? tmp461 : tmp462;
  assign tmp453 = s2 ? tmp454 : tmp460;
  assign tmp450 = s3 ? tmp451 : tmp453;
  assign tmp468 = ~(s0 ? tmp464 : tmp463);
  assign tmp467 = s1 ? tmp335 : tmp468;
  assign tmp470 = s0 ? tmp452 : tmp174;
  assign tmp469 = s1 ? tmp470 : tmp33;
  assign tmp466 = s2 ? tmp467 : tmp469;
  assign tmp473 = ~(s0 ? 1 : tmp457);
  assign tmp472 = s1 ? tmp463 : tmp473;
  assign tmp471 = ~(s2 ? tmp342 : tmp472);
  assign tmp465 = s3 ? tmp466 : tmp471;
  assign tmp449 = s4 ? tmp450 : tmp465;
  assign tmp478 = s1 ? tmp328 : tmp456;
  assign tmp481 = l1 ? 1 : tmp228;
  assign tmp480 = s0 ? tmp481 : tmp173;
  assign tmp479 = s1 ? tmp351 : tmp480;
  assign tmp477 = s2 ? tmp478 : tmp479;
  assign tmp484 = l1 ? 1 : tmp173;
  assign tmp485 = l1 ? 1 : tmp193;
  assign tmp483 = s1 ? tmp484 : tmp485;
  assign tmp487 = ~(l1 ? tmp120 : tmp226);
  assign tmp486 = s1 ? 1 : tmp487;
  assign tmp482 = s2 ? tmp483 : tmp486;
  assign tmp476 = s3 ? tmp477 : tmp482;
  assign tmp492 = ~(l1 ? tmp120 : tmp24);
  assign tmp491 = s0 ? 1 : tmp492;
  assign tmp490 = s1 ? tmp491 : tmp362;
  assign tmp489 = s2 ? tmp490 : tmp364;
  assign tmp488 = s3 ? tmp489 : tmp365;
  assign tmp475 = s4 ? tmp476 : tmp488;
  assign tmp497 = s0 ? tmp485 : 1;
  assign tmp496 = s1 ? tmp497 : 1;
  assign tmp495 = s2 ? tmp496 : tmp443;
  assign tmp494 = s3 ? tmp495 : 1;
  assign tmp498 = s3 ? tmp377 : 1;
  assign tmp493 = s4 ? tmp494 : tmp498;
  assign tmp474 = s5 ? tmp475 : tmp493;
  assign tmp448 = ~(s6 ? tmp449 : tmp474);
  assign tmp447 = s7 ? 1 : tmp448;
  assign tmp446 = s8 ? tmp378 : tmp447;
  assign tmp303 = s9 ? tmp304 : tmp446;
  assign tmp507 = s0 ? tmp336 : tmp312;
  assign tmp508 = s0 ? tmp326 : tmp312;
  assign tmp506 = s1 ? tmp507 : tmp508;
  assign tmp510 = s0 ? tmp326 : tmp173;
  assign tmp512 = l1 ? tmp120 : tmp384;
  assign tmp511 = ~(s0 ? tmp120 : tmp512);
  assign tmp509 = s1 ? tmp510 : tmp511;
  assign tmp505 = s2 ? tmp506 : tmp509;
  assign tmp504 = s3 ? tmp309 : tmp505;
  assign tmp516 = ~(s0 ? tmp512 : tmp120);
  assign tmp515 = s1 ? tmp335 : tmp516;
  assign tmp518 = s0 ? tmp310 : tmp174;
  assign tmp517 = s1 ? tmp518 : tmp33;
  assign tmp514 = s2 ? tmp515 : tmp517;
  assign tmp521 = ~(s0 ? 1 : tmp312);
  assign tmp520 = s1 ? tmp120 : tmp521;
  assign tmp519 = ~(s2 ? tmp342 : tmp520);
  assign tmp513 = s3 ? tmp514 : tmp519;
  assign tmp503 = s4 ? tmp504 : tmp513;
  assign tmp526 = s1 ? tmp328 : tmp336;
  assign tmp528 = ~(s0 ? tmp120 : tmp316);
  assign tmp527 = s1 ? tmp326 : tmp528;
  assign tmp525 = s2 ? tmp526 : tmp527;
  assign tmp530 = s1 ? tmp355 : tmp442;
  assign tmp531 = s1 ? 1 : tmp312;
  assign tmp529 = s2 ? tmp530 : tmp531;
  assign tmp524 = s3 ? tmp525 : tmp529;
  assign tmp533 = s2 ? tmp490 : tmp336;
  assign tmp536 = s0 ? tmp355 : 1;
  assign tmp535 = s1 ? tmp536 : 1;
  assign tmp534 = s2 ? tmp535 : 1;
  assign tmp532 = s3 ? tmp533 : tmp534;
  assign tmp523 = s4 ? tmp524 : tmp532;
  assign tmp537 = s4 ? tmp438 : tmp444;
  assign tmp522 = s5 ? tmp523 : tmp537;
  assign tmp502 = ~(s6 ? tmp503 : tmp522);
  assign tmp501 = s7 ? 1 : tmp502;
  assign tmp500 = s8 ? tmp501 : 1;
  assign tmp540 = s6 ? tmp307 : tmp345;
  assign tmp541 = s6 ? tmp449 : tmp474;
  assign tmp539 = s7 ? tmp540 : tmp541;
  assign tmp542 = ~(s7 ? tmp379 : tmp502);
  assign tmp538 = ~(s8 ? tmp539 : tmp542);
  assign tmp499 = s9 ? tmp500 : tmp538;
  assign tmp302 = s10 ? tmp303 : tmp499;
  assign tmp552 = l1 ? tmp19 : tmp203;
  assign tmp553 = ~(l1 ? tmp311 : tmp322);
  assign tmp551 = ~(s0 ? tmp552 : tmp553);
  assign tmp550 = s1 ? tmp311 : tmp551;
  assign tmp556 = s0 ? tmp322 : tmp311;
  assign tmp558 = l1 ? tmp311 : tmp322;
  assign tmp557 = s0 ? tmp558 : tmp311;
  assign tmp555 = s1 ? tmp556 : tmp557;
  assign tmp561 = ~(l1 ? 1 : tmp203);
  assign tmp560 = s0 ? tmp558 : tmp561;
  assign tmp559 = s1 ? tmp560 : tmp311;
  assign tmp554 = s2 ? tmp555 : tmp559;
  assign tmp549 = s3 ? tmp550 : tmp554;
  assign tmp566 = ~(l1 ? tmp19 : tmp203);
  assign tmp565 = s0 ? tmp322 : tmp566;
  assign tmp564 = s1 ? tmp565 : tmp311;
  assign tmp568 = s0 ? tmp311 : 0;
  assign tmp569 = ~(l1 ? tmp19 : 0);
  assign tmp567 = s1 ? tmp568 : tmp569;
  assign tmp563 = s2 ? tmp564 : tmp567;
  assign tmp571 = s1 ? tmp552 : 0;
  assign tmp573 = s0 ? 1 : tmp311;
  assign tmp572 = ~(s1 ? tmp311 : tmp573);
  assign tmp570 = ~(s2 ? tmp571 : tmp572);
  assign tmp562 = s3 ? tmp563 : tmp570;
  assign tmp548 = s4 ? tmp549 : tmp562;
  assign tmp578 = s1 ? tmp560 : tmp322;
  assign tmp580 = l1 ? tmp311 : 1;
  assign tmp582 = l1 ? 1 : tmp311;
  assign tmp581 = s0 ? tmp582 : tmp31;
  assign tmp579 = s1 ? tmp580 : tmp581;
  assign tmp577 = s2 ? tmp578 : tmp579;
  assign tmp585 = l1 ? 1 : tmp322;
  assign tmp584 = s1 ? tmp585 : 1;
  assign tmp587 = s0 ? tmp580 : 1;
  assign tmp586 = s1 ? 1 : tmp587;
  assign tmp583 = s2 ? tmp584 : tmp586;
  assign tmp576 = s3 ? tmp577 : tmp583;
  assign tmp591 = s0 ? 1 : tmp580;
  assign tmp593 = l1 ? tmp19 : 0;
  assign tmp592 = ~(s0 ? tmp593 : 0);
  assign tmp590 = s1 ? tmp591 : tmp592;
  assign tmp594 = l1 ? tmp322 : 1;
  assign tmp589 = s2 ? tmp590 : tmp594;
  assign tmp588 = s3 ? tmp589 : 1;
  assign tmp575 = s4 ? tmp576 : tmp588;
  assign tmp574 = s5 ? tmp575 : 1;
  assign tmp547 = ~(s6 ? tmp548 : tmp574);
  assign tmp546 = s7 ? 1 : tmp547;
  assign tmp601 = ~(l2 ? 1 : tmp312);
  assign tmp600 = l1 ? tmp330 : tmp601;
  assign tmp603 = l1 ? tmp74 : tmp203;
  assign tmp604 = l1 ? tmp330 : tmp32;
  assign tmp602 = s0 ? tmp603 : tmp604;
  assign tmp599 = s1 ? tmp600 : tmp602;
  assign tmp608 = l1 ? tmp392 : tmp32;
  assign tmp607 = s0 ? tmp608 : tmp600;
  assign tmp609 = s0 ? tmp604 : tmp600;
  assign tmp606 = s1 ? tmp607 : tmp609;
  assign tmp611 = s0 ? tmp604 : tmp375;
  assign tmp610 = s1 ? tmp611 : tmp600;
  assign tmp605 = s2 ? tmp606 : tmp610;
  assign tmp598 = s3 ? tmp599 : tmp605;
  assign tmp615 = s0 ? tmp608 : tmp603;
  assign tmp614 = s1 ? tmp615 : tmp600;
  assign tmp617 = s0 ? tmp600 : 1;
  assign tmp618 = l1 ? tmp74 : 0;
  assign tmp616 = s1 ? tmp617 : tmp618;
  assign tmp613 = s2 ? tmp614 : tmp616;
  assign tmp620 = s1 ? tmp603 : 0;
  assign tmp623 = ~(l1 ? tmp330 : tmp601);
  assign tmp622 = ~(s0 ? 1 : tmp623);
  assign tmp621 = s1 ? tmp600 : tmp622;
  assign tmp619 = s2 ? tmp620 : tmp621;
  assign tmp612 = s3 ? tmp613 : tmp619;
  assign tmp597 = s4 ? tmp598 : tmp612;
  assign tmp628 = s1 ? tmp611 : tmp608;
  assign tmp630 = l1 ? tmp330 : 0;
  assign tmp632 = l1 ? tmp373 : tmp601;
  assign tmp631 = s0 ? tmp632 : tmp375;
  assign tmp629 = s1 ? tmp630 : tmp631;
  assign tmp627 = s2 ? tmp628 : tmp629;
  assign tmp635 = l1 ? tmp373 : tmp32;
  assign tmp634 = s1 ? tmp635 : 0;
  assign tmp638 = l1 ? tmp373 : 0;
  assign tmp637 = ~(s0 ? tmp630 : tmp638);
  assign tmp636 = ~(s1 ? 1 : tmp637);
  assign tmp633 = s2 ? tmp634 : tmp636;
  assign tmp626 = s3 ? tmp627 : tmp633;
  assign tmp643 = ~(l1 ? tmp330 : 0);
  assign tmp642 = s0 ? 1 : tmp643;
  assign tmp644 = ~(s0 ? tmp618 : tmp174);
  assign tmp641 = s1 ? tmp642 : tmp644;
  assign tmp645 = ~(l1 ? tmp392 : 0);
  assign tmp640 = s2 ? tmp641 : tmp645;
  assign tmp648 = s0 ? 1 : tmp436;
  assign tmp647 = s1 ? tmp648 : 1;
  assign tmp646 = s2 ? tmp647 : 1;
  assign tmp639 = ~(s3 ? tmp640 : tmp646);
  assign tmp625 = s4 ? tmp626 : tmp639;
  assign tmp624 = s5 ? tmp625 : 0;
  assign tmp596 = s6 ? tmp597 : tmp624;
  assign tmp595 = s7 ? 1 : tmp596;
  assign tmp545 = s8 ? tmp546 : tmp595;
  assign tmp655 = l1 ? tmp311 : tmp26;
  assign tmp654 = s1 ? tmp655 : tmp551;
  assign tmp659 = l1 ? tmp322 : tmp31;
  assign tmp660 = ~(l1 ? tmp120 : tmp102);
  assign tmp658 = s0 ? tmp659 : tmp660;
  assign tmp662 = l1 ? tmp311 : tmp31;
  assign tmp661 = s0 ? tmp662 : tmp660;
  assign tmp657 = s1 ? tmp658 : tmp661;
  assign tmp664 = s0 ? tmp662 : tmp31;
  assign tmp663 = s1 ? tmp664 : tmp660;
  assign tmp656 = s2 ? tmp657 : tmp663;
  assign tmp653 = s3 ? tmp654 : tmp656;
  assign tmp667 = s1 ? tmp565 : tmp660;
  assign tmp669 = s0 ? tmp655 : tmp174;
  assign tmp668 = s1 ? tmp669 : tmp569;
  assign tmp666 = s2 ? tmp667 : tmp668;
  assign tmp672 = l1 ? tmp120 : tmp102;
  assign tmp673 = ~(s0 ? 1 : tmp660);
  assign tmp671 = s1 ? tmp672 : tmp673;
  assign tmp670 = ~(s2 ? tmp571 : tmp671);
  assign tmp665 = s3 ? tmp666 : tmp670;
  assign tmp652 = s4 ? tmp653 : tmp665;
  assign tmp678 = s1 ? tmp560 : tmp659;
  assign tmp681 = l1 ? 1 : tmp26;
  assign tmp680 = s0 ? tmp681 : tmp131;
  assign tmp679 = s1 ? tmp580 : tmp680;
  assign tmp677 = s2 ? tmp678 : tmp679;
  assign tmp683 = s1 ? tmp131 : 1;
  assign tmp686 = l1 ? tmp120 : 0;
  assign tmp685 = ~(s0 ? tmp686 : 0);
  assign tmp684 = s1 ? 1 : tmp685;
  assign tmp682 = s2 ? tmp683 : tmp684;
  assign tmp676 = s3 ? tmp677 : tmp682;
  assign tmp691 = ~(l1 ? tmp120 : 0);
  assign tmp690 = s0 ? 1 : tmp691;
  assign tmp689 = s1 ? tmp690 : tmp592;
  assign tmp688 = s2 ? tmp689 : tmp594;
  assign tmp687 = s3 ? tmp688 : 1;
  assign tmp675 = s4 ? tmp676 : tmp687;
  assign tmp674 = s5 ? tmp675 : 1;
  assign tmp651 = ~(s6 ? tmp652 : tmp674);
  assign tmp650 = s7 ? 1 : tmp651;
  assign tmp649 = s8 ? tmp595 : tmp650;
  assign tmp544 = s9 ? tmp545 : tmp649;
  assign tmp701 = ~(l1 ? tmp120 : tmp601);
  assign tmp700 = s0 ? tmp322 : tmp701;
  assign tmp702 = s0 ? tmp558 : tmp701;
  assign tmp699 = s1 ? tmp700 : tmp702;
  assign tmp704 = s0 ? tmp558 : tmp31;
  assign tmp703 = s1 ? tmp704 : tmp701;
  assign tmp698 = s2 ? tmp699 : tmp703;
  assign tmp697 = s3 ? tmp550 : tmp698;
  assign tmp707 = s1 ? tmp565 : tmp701;
  assign tmp709 = s0 ? tmp311 : tmp174;
  assign tmp708 = s1 ? tmp709 : tmp569;
  assign tmp706 = s2 ? tmp707 : tmp708;
  assign tmp712 = l1 ? tmp120 : tmp601;
  assign tmp713 = ~(s0 ? 1 : tmp701);
  assign tmp711 = s1 ? tmp712 : tmp713;
  assign tmp710 = ~(s2 ? tmp571 : tmp711);
  assign tmp705 = s3 ? tmp706 : tmp710;
  assign tmp696 = s4 ? tmp697 : tmp705;
  assign tmp719 = s0 ? tmp582 : tmp131;
  assign tmp718 = s1 ? tmp580 : tmp719;
  assign tmp717 = s2 ? tmp578 : tmp718;
  assign tmp720 = s2 ? tmp584 : tmp684;
  assign tmp716 = s3 ? tmp717 : tmp720;
  assign tmp715 = s4 ? tmp716 : tmp687;
  assign tmp714 = s5 ? tmp715 : 1;
  assign tmp695 = ~(s6 ? tmp696 : tmp714);
  assign tmp694 = s7 ? 1 : tmp695;
  assign tmp693 = s8 ? tmp694 : 1;
  assign tmp723 = s6 ? tmp548 : tmp574;
  assign tmp724 = s6 ? tmp652 : tmp674;
  assign tmp722 = s7 ? tmp723 : tmp724;
  assign tmp725 = ~(s7 ? tmp596 : tmp695);
  assign tmp721 = ~(s8 ? tmp722 : tmp725);
  assign tmp692 = s9 ? tmp693 : tmp721;
  assign tmp543 = s10 ? tmp544 : tmp692;
  assign tmp301 = s12 ? tmp302 : tmp543;
  assign tmp5 = s13 ? tmp6 : tmp301;
  assign tmp736 = l1 ? 1 : tmp313;
  assign tmp737 = s0 ? tmp484 : tmp355;
  assign tmp735 = s1 ? tmp736 : tmp737;
  assign tmp741 = l1 ? 1 : tmp323;
  assign tmp742 = l1 ? 1 : tmp324;
  assign tmp740 = s0 ? tmp741 : tmp742;
  assign tmp743 = s0 ? tmp355 : tmp742;
  assign tmp739 = s1 ? tmp740 : tmp743;
  assign tmp745 = s0 ? tmp355 : tmp83;
  assign tmp746 = s0 ? tmp742 : tmp736;
  assign tmp744 = s1 ? tmp745 : tmp746;
  assign tmp738 = s2 ? tmp739 : tmp744;
  assign tmp734 = s3 ? tmp735 : tmp738;
  assign tmp750 = s0 ? tmp736 : tmp742;
  assign tmp749 = s1 ? tmp745 : tmp750;
  assign tmp752 = s0 ? tmp736 : tmp83;
  assign tmp751 = s1 ? tmp752 : tmp355;
  assign tmp748 = s2 ? tmp749 : tmp751;
  assign tmp754 = s1 ? tmp484 : 1;
  assign tmp756 = s0 ? tmp742 : tmp324;
  assign tmp757 = s0 ? 1 : tmp742;
  assign tmp755 = s1 ? tmp756 : tmp757;
  assign tmp753 = s2 ? tmp754 : tmp755;
  assign tmp747 = s3 ? tmp748 : tmp753;
  assign tmp733 = s4 ? tmp734 : tmp747;
  assign tmp762 = s1 ? tmp745 : tmp741;
  assign tmp763 = s1 ? tmp221 : tmp352;
  assign tmp761 = s2 ? tmp762 : tmp763;
  assign tmp767 = l1 ? 1 : tmp356;
  assign tmp766 = s0 ? tmp767 : 1;
  assign tmp765 = s1 ? 1 : tmp766;
  assign tmp764 = s2 ? tmp354 : tmp765;
  assign tmp760 = s3 ? tmp761 : tmp764;
  assign tmp771 = s0 ? 1 : tmp221;
  assign tmp772 = s0 ? tmp83 : 1;
  assign tmp770 = s1 ? tmp771 : tmp772;
  assign tmp769 = s2 ? tmp770 : tmp221;
  assign tmp768 = s3 ? tmp769 : tmp365;
  assign tmp759 = s4 ? tmp760 : tmp768;
  assign tmp758 = s5 ? tmp759 : tmp368;
  assign tmp732 = ~(s6 ? tmp733 : tmp758);
  assign tmp731 = s7 ? 1 : tmp732;
  assign tmp780 = l3 ? 1 : tmp17;
  assign tmp779 = ~(l2 ? tmp780 : tmp120);
  assign tmp778 = l1 ? 1 : tmp779;
  assign tmp783 = ~(l2 ? tmp780 : 1);
  assign tmp782 = l1 ? 1 : tmp783;
  assign tmp785 = ~(l2 ? tmp780 : tmp19);
  assign tmp784 = l1 ? 1 : tmp785;
  assign tmp781 = s0 ? tmp782 : tmp784;
  assign tmp777 = s1 ? tmp778 : tmp781;
  assign tmp788 = s0 ? tmp784 : tmp742;
  assign tmp787 = s1 ? tmp740 : tmp788;
  assign tmp790 = s0 ? tmp784 : tmp83;
  assign tmp791 = s0 ? tmp742 : tmp778;
  assign tmp789 = s1 ? tmp790 : tmp791;
  assign tmp786 = s2 ? tmp787 : tmp789;
  assign tmp776 = s3 ? tmp777 : tmp786;
  assign tmp795 = s0 ? tmp778 : tmp742;
  assign tmp794 = s1 ? tmp790 : tmp795;
  assign tmp797 = s0 ? tmp778 : tmp83;
  assign tmp798 = l1 ? 1 : tmp69;
  assign tmp796 = s1 ? tmp797 : tmp798;
  assign tmp793 = s2 ? tmp794 : tmp796;
  assign tmp800 = s1 ? tmp782 : 1;
  assign tmp803 = ~(l1 ? 1 : tmp324);
  assign tmp802 = ~(s0 ? tmp17 : tmp803);
  assign tmp801 = s1 ? tmp742 : tmp802;
  assign tmp799 = s2 ? tmp800 : tmp801;
  assign tmp792 = s3 ? tmp793 : tmp799;
  assign tmp775 = s4 ? tmp776 : tmp792;
  assign tmp808 = s1 ? tmp790 : tmp741;
  assign tmp811 = ~(l2 ? tmp780 : 0);
  assign tmp810 = l1 ? 1 : tmp811;
  assign tmp812 = s0 ? tmp742 : tmp83;
  assign tmp809 = s1 ? tmp810 : tmp812;
  assign tmp807 = s2 ? tmp808 : tmp809;
  assign tmp814 = s1 ? tmp784 : tmp356;
  assign tmp816 = ~(l1 ? 1 : tmp356);
  assign tmp815 = ~(s1 ? tmp93 : tmp816);
  assign tmp813 = s2 ? tmp814 : tmp815;
  assign tmp806 = s3 ? tmp807 : tmp813;
  assign tmp820 = s0 ? 1 : tmp810;
  assign tmp822 = l1 ? 1 : tmp21;
  assign tmp821 = s0 ? tmp83 : tmp822;
  assign tmp819 = s1 ? tmp820 : tmp821;
  assign tmp818 = s2 ? tmp819 : tmp810;
  assign tmp825 = s0 ? tmp810 : tmp767;
  assign tmp824 = s1 ? tmp825 : 1;
  assign tmp823 = s2 ? tmp824 : 1;
  assign tmp817 = s3 ? tmp818 : tmp823;
  assign tmp805 = s4 ? tmp806 : tmp817;
  assign tmp830 = ~(l1 ? 1 : tmp21);
  assign tmp829 = s1 ? tmp372 : tmp830;
  assign tmp828 = s2 ? tmp829 : tmp374;
  assign tmp827 = s3 ? tmp828 : 0;
  assign tmp832 = s2 ? tmp75 : tmp810;
  assign tmp831 = ~(s3 ? tmp832 : 1);
  assign tmp826 = ~(s4 ? tmp827 : tmp831);
  assign tmp804 = s5 ? tmp805 : tmp826;
  assign tmp774 = ~(s6 ? tmp775 : tmp804);
  assign tmp773 = s7 ? 1 : tmp774;
  assign tmp730 = s8 ? tmp731 : tmp773;
  assign tmp840 = ~(l2 ? tmp780 : tmp17);
  assign tmp839 = l1 ? 1 : tmp840;
  assign tmp841 = s0 ? tmp782 : tmp798;
  assign tmp838 = s1 ? tmp839 : tmp841;
  assign tmp844 = s0 ? tmp782 : tmp822;
  assign tmp843 = s1 ? tmp821 : tmp844;
  assign tmp846 = s0 ? tmp782 : tmp83;
  assign tmp847 = s0 ? tmp822 : tmp839;
  assign tmp845 = s1 ? tmp846 : tmp847;
  assign tmp842 = s2 ? tmp843 : tmp845;
  assign tmp837 = s3 ? tmp838 : tmp842;
  assign tmp851 = s0 ? tmp798 : tmp83;
  assign tmp852 = s0 ? tmp839 : tmp822;
  assign tmp850 = s1 ? tmp851 : tmp852;
  assign tmp854 = s0 ? tmp839 : tmp83;
  assign tmp853 = s1 ? tmp854 : tmp798;
  assign tmp849 = s2 ? tmp850 : tmp853;
  assign tmp857 = ~(s0 ? tmp17 : tmp830);
  assign tmp856 = s1 ? tmp822 : tmp857;
  assign tmp855 = s2 ? tmp800 : tmp856;
  assign tmp848 = s3 ? tmp849 : tmp855;
  assign tmp836 = s4 ? tmp837 : tmp848;
  assign tmp862 = s1 ? tmp851 : tmp83;
  assign tmp864 = s0 ? tmp822 : tmp83;
  assign tmp863 = s1 ? tmp798 : tmp864;
  assign tmp861 = s2 ? tmp862 : tmp863;
  assign tmp866 = s1 ? tmp782 : tmp822;
  assign tmp867 = ~(s1 ? tmp93 : tmp830);
  assign tmp865 = s2 ? tmp866 : tmp867;
  assign tmp860 = s3 ? tmp861 : tmp865;
  assign tmp869 = s2 ? tmp819 : tmp798;
  assign tmp872 = s0 ? tmp798 : tmp767;
  assign tmp871 = s1 ? tmp872 : 1;
  assign tmp870 = s2 ? tmp871 : 1;
  assign tmp868 = s3 ? tmp869 : tmp870;
  assign tmp859 = s4 ? tmp860 : tmp868;
  assign tmp877 = s0 ? tmp822 : 1;
  assign tmp876 = s1 ? tmp877 : tmp822;
  assign tmp878 = s1 ? tmp83 : 1;
  assign tmp875 = s2 ? tmp876 : tmp878;
  assign tmp874 = s3 ? tmp875 : 1;
  assign tmp880 = s2 ? tmp75 : tmp798;
  assign tmp879 = s3 ? tmp880 : 1;
  assign tmp873 = s4 ? tmp874 : tmp879;
  assign tmp858 = s5 ? tmp859 : tmp873;
  assign tmp835 = ~(s6 ? tmp836 : tmp858);
  assign tmp834 = s7 ? 1 : tmp835;
  assign tmp833 = s8 ? tmp773 : tmp834;
  assign tmp729 = s9 ? tmp730 : tmp833;
  assign tmp882 = s8 ? tmp773 : 1;
  assign tmp885 = s6 ? tmp733 : tmp758;
  assign tmp886 = s6 ? tmp836 : tmp858;
  assign tmp884 = s7 ? tmp885 : tmp886;
  assign tmp887 = s6 ? tmp775 : tmp804;
  assign tmp883 = ~(s8 ? tmp884 : tmp887);
  assign tmp881 = s9 ? tmp882 : tmp883;
  assign tmp728 = s10 ? tmp729 : tmp881;
  assign tmp898 = l3 ? 1 : tmp21;
  assign tmp897 = l2 ? tmp19 : tmp898;
  assign tmp896 = l1 ? tmp74 : tmp897;
  assign tmp901 = l2 ? 1 : tmp898;
  assign tmp900 = l1 ? tmp901 : tmp897;
  assign tmp899 = s0 ? tmp19 : tmp900;
  assign tmp895 = s1 ? tmp896 : tmp899;
  assign tmp903 = s0 ? tmp406 : tmp900;
  assign tmp905 = s0 ? tmp406 : 1;
  assign tmp904 = s1 ? tmp905 : tmp900;
  assign tmp902 = s2 ? tmp903 : tmp904;
  assign tmp894 = s3 ? tmp895 : tmp902;
  assign tmp909 = s0 ? tmp896 : tmp363;
  assign tmp908 = s1 ? tmp909 : tmp900;
  assign tmp911 = s0 ? tmp896 : 1;
  assign tmp910 = s1 ? tmp911 : tmp19;
  assign tmp907 = s2 ? tmp908 : tmp910;
  assign tmp913 = s1 ? tmp19 : tmp316;
  assign tmp917 = ~(l2 ? tmp19 : tmp898);
  assign tmp916 = ~(l1 ? tmp17 : tmp917);
  assign tmp915 = s0 ? tmp900 : tmp916;
  assign tmp918 = s0 ? tmp397 : tmp900;
  assign tmp914 = s1 ? tmp915 : tmp918;
  assign tmp912 = s2 ? tmp913 : tmp914;
  assign tmp906 = s3 ? tmp907 : tmp912;
  assign tmp893 = s4 ? tmp894 : tmp906;
  assign tmp924 = s0 ? tmp900 : 1;
  assign tmp923 = s1 ? tmp924 : tmp406;
  assign tmp927 = l2 ? tmp19 : tmp21;
  assign tmp926 = l1 ? tmp901 : tmp927;
  assign tmp929 = l1 ? tmp17 : tmp917;
  assign tmp928 = ~(s0 ? tmp929 : 0);
  assign tmp925 = s1 ? tmp926 : tmp928;
  assign tmp922 = s2 ? tmp923 : tmp925;
  assign tmp933 = ~(l2 ? tmp19 : tmp21);
  assign tmp932 = ~(l1 ? tmp17 : tmp933);
  assign tmp931 = s1 ? tmp406 : tmp932;
  assign tmp935 = s0 ? tmp397 : 1;
  assign tmp936 = s0 ? tmp926 : tmp932;
  assign tmp934 = s1 ? tmp935 : tmp936;
  assign tmp930 = s2 ? tmp931 : tmp934;
  assign tmp921 = s3 ? tmp922 : tmp930;
  assign tmp940 = s0 ? tmp397 : tmp926;
  assign tmp941 = s0 ? tmp363 : 0;
  assign tmp939 = s1 ? tmp940 : tmp941;
  assign tmp942 = l1 ? tmp74 : tmp927;
  assign tmp938 = s2 ? tmp939 : tmp942;
  assign tmp946 = l1 ? tmp31 : tmp927;
  assign tmp948 = ~(l2 ? 1 : tmp17);
  assign tmp947 = l1 ? tmp74 : tmp948;
  assign tmp945 = s0 ? tmp946 : tmp947;
  assign tmp944 = s1 ? tmp945 : tmp932;
  assign tmp949 = s1 ? 1 : tmp316;
  assign tmp943 = s2 ? tmp944 : tmp949;
  assign tmp937 = s3 ? tmp938 : tmp943;
  assign tmp920 = s4 ? tmp921 : tmp937;
  assign tmp955 = l1 ? tmp17 : tmp933;
  assign tmp954 = s0 ? tmp955 : 0;
  assign tmp953 = s1 ? tmp954 : tmp54;
  assign tmp956 = ~(s1 ? tmp31 : tmp174);
  assign tmp952 = s2 ? tmp953 : tmp956;
  assign tmp959 = l1 ? tmp31 : tmp948;
  assign tmp958 = s1 ? tmp375 : tmp959;
  assign tmp957 = ~(s2 ? 1 : tmp958);
  assign tmp951 = s3 ? tmp952 : tmp957;
  assign tmp962 = s1 ? 1 : tmp397;
  assign tmp963 = l1 ? tmp26 : tmp927;
  assign tmp961 = s2 ? tmp962 : tmp963;
  assign tmp966 = l2 ? 1 : tmp17;
  assign tmp965 = ~(l1 ? tmp17 : tmp966);
  assign tmp964 = s1 ? 1 : tmp965;
  assign tmp960 = ~(s3 ? tmp961 : tmp964);
  assign tmp950 = ~(s4 ? tmp951 : tmp960);
  assign tmp919 = s5 ? tmp920 : tmp950;
  assign tmp892 = ~(s6 ? tmp893 : tmp919);
  assign tmp891 = s7 ? 1 : tmp892;
  assign tmp973 = l2 ? tmp17 : tmp898;
  assign tmp972 = l1 ? tmp74 : tmp973;
  assign tmp975 = l1 ? tmp74 : tmp116;
  assign tmp976 = l1 ? tmp901 : tmp973;
  assign tmp974 = s0 ? tmp975 : tmp976;
  assign tmp971 = s1 ? tmp972 : tmp974;
  assign tmp981 = l2 ? tmp780 : tmp898;
  assign tmp980 = l1 ? tmp901 : tmp981;
  assign tmp979 = s0 ? tmp74 : tmp980;
  assign tmp983 = l1 ? tmp74 : tmp392;
  assign tmp982 = s0 ? tmp983 : tmp980;
  assign tmp978 = s1 ? tmp979 : tmp982;
  assign tmp985 = s0 ? tmp983 : 1;
  assign tmp986 = s0 ? tmp980 : tmp976;
  assign tmp984 = s1 ? tmp985 : tmp986;
  assign tmp977 = s2 ? tmp978 : tmp984;
  assign tmp970 = s3 ? tmp971 : tmp977;
  assign tmp990 = s0 ? tmp972 : tmp237;
  assign tmp991 = s0 ? tmp976 : tmp980;
  assign tmp989 = s1 ? tmp990 : tmp991;
  assign tmp993 = s0 ? tmp972 : 1;
  assign tmp994 = l1 ? tmp74 : tmp17;
  assign tmp992 = s1 ? tmp993 : tmp994;
  assign tmp988 = s2 ? tmp989 : tmp992;
  assign tmp996 = s1 ? tmp975 : tmp316;
  assign tmp999 = l1 ? tmp26 : tmp981;
  assign tmp998 = s0 ? tmp980 : tmp999;
  assign tmp1002 = l2 ? tmp780 : 1;
  assign tmp1001 = l1 ? 1 : tmp1002;
  assign tmp1000 = s0 ? tmp1001 : tmp980;
  assign tmp997 = s1 ? tmp998 : tmp1000;
  assign tmp995 = s2 ? tmp996 : tmp997;
  assign tmp987 = s3 ? tmp988 : tmp995;
  assign tmp969 = s4 ? tmp970 : tmp987;
  assign tmp1008 = s0 ? tmp976 : 1;
  assign tmp1007 = s1 ? tmp1008 : tmp74;
  assign tmp1011 = l2 ? tmp17 : tmp21;
  assign tmp1010 = l1 ? tmp901 : tmp1011;
  assign tmp1012 = s0 ? tmp999 : 1;
  assign tmp1009 = s1 ? tmp1010 : tmp1012;
  assign tmp1006 = s2 ? tmp1007 : tmp1009;
  assign tmp1016 = ~(l2 ? tmp780 : tmp21);
  assign tmp1015 = ~(l1 ? tmp17 : tmp1016);
  assign tmp1014 = s1 ? tmp983 : tmp1015;
  assign tmp1018 = s0 ? tmp1001 : 1;
  assign tmp1021 = l2 ? tmp780 : tmp21;
  assign tmp1020 = l1 ? tmp901 : tmp1021;
  assign tmp1022 = l1 ? tmp26 : tmp1021;
  assign tmp1019 = s0 ? tmp1020 : tmp1022;
  assign tmp1017 = s1 ? tmp1018 : tmp1019;
  assign tmp1013 = s2 ? tmp1014 : tmp1017;
  assign tmp1005 = s3 ? tmp1006 : tmp1013;
  assign tmp1026 = s0 ? tmp397 : tmp1010;
  assign tmp1027 = s0 ? tmp237 : tmp373;
  assign tmp1025 = s1 ? tmp1026 : tmp1027;
  assign tmp1028 = l1 ? tmp74 : tmp1011;
  assign tmp1024 = s2 ? tmp1025 : tmp1028;
  assign tmp1032 = l1 ? tmp31 : tmp1011;
  assign tmp1031 = s0 ? tmp1032 : tmp1028;
  assign tmp1030 = s1 ? tmp1031 : tmp932;
  assign tmp1029 = s2 ? tmp1030 : tmp949;
  assign tmp1023 = s3 ? tmp1024 : tmp1029;
  assign tmp1004 = s4 ? tmp1005 : tmp1023;
  assign tmp1038 = l1 ? tmp17 : tmp1016;
  assign tmp1037 = s0 ? tmp1038 : 0;
  assign tmp1039 = ~(l1 ? 1 : tmp17);
  assign tmp1036 = s1 ? tmp1037 : tmp1039;
  assign tmp1035 = s2 ? tmp1036 : tmp956;
  assign tmp1034 = s3 ? tmp1035 : tmp957;
  assign tmp1042 = s1 ? 1 : tmp1001;
  assign tmp1043 = l1 ? tmp26 : tmp1011;
  assign tmp1041 = s2 ? tmp1042 : tmp1043;
  assign tmp1040 = ~(s3 ? tmp1041 : tmp964);
  assign tmp1033 = ~(s4 ? tmp1034 : tmp1040);
  assign tmp1003 = s5 ? tmp1004 : tmp1033;
  assign tmp968 = ~(s6 ? tmp969 : tmp1003);
  assign tmp967 = s7 ? 1 : tmp968;
  assign tmp890 = s8 ? tmp891 : tmp967;
  assign tmp889 = s9 ? tmp890 : tmp967;
  assign tmp1045 = s8 ? tmp967 : 1;
  assign tmp1048 = s6 ? tmp893 : tmp919;
  assign tmp1054 = l1 ? tmp901 : tmp116;
  assign tmp1053 = s0 ? tmp975 : tmp1054;
  assign tmp1052 = s1 ? tmp975 : tmp1053;
  assign tmp1058 = l1 ? tmp901 : tmp1002;
  assign tmp1057 = s0 ? tmp237 : tmp1058;
  assign tmp1059 = s0 ? tmp975 : tmp1058;
  assign tmp1056 = s1 ? tmp1057 : tmp1059;
  assign tmp1061 = s0 ? tmp975 : 1;
  assign tmp1062 = s0 ? tmp1058 : tmp1054;
  assign tmp1060 = s1 ? tmp1061 : tmp1062;
  assign tmp1055 = s2 ? tmp1056 : tmp1060;
  assign tmp1051 = s3 ? tmp1052 : tmp1055;
  assign tmp1066 = s0 ? tmp975 : tmp237;
  assign tmp1067 = s0 ? tmp1054 : tmp1058;
  assign tmp1065 = s1 ? tmp1066 : tmp1067;
  assign tmp1068 = s1 ? tmp1061 : tmp994;
  assign tmp1064 = s2 ? tmp1065 : tmp1068;
  assign tmp1072 = l1 ? tmp26 : tmp1002;
  assign tmp1071 = s0 ? tmp1058 : tmp1072;
  assign tmp1073 = s0 ? tmp1001 : tmp1058;
  assign tmp1070 = s1 ? tmp1071 : tmp1073;
  assign tmp1069 = s2 ? tmp996 : tmp1070;
  assign tmp1063 = s3 ? tmp1064 : tmp1069;
  assign tmp1050 = s4 ? tmp1051 : tmp1063;
  assign tmp1079 = s0 ? tmp1054 : 1;
  assign tmp1078 = s1 ? tmp1079 : tmp237;
  assign tmp1081 = s0 ? tmp1072 : 1;
  assign tmp1080 = s1 ? tmp1054 : tmp1081;
  assign tmp1077 = s2 ? tmp1078 : tmp1080;
  assign tmp1084 = ~(l1 ? tmp17 : tmp783);
  assign tmp1083 = s1 ? tmp975 : tmp1084;
  assign tmp1085 = s1 ? tmp1018 : tmp1071;
  assign tmp1082 = s2 ? tmp1083 : tmp1085;
  assign tmp1076 = s3 ? tmp1077 : tmp1082;
  assign tmp1089 = s0 ? tmp397 : tmp1054;
  assign tmp1088 = s1 ? tmp1089 : tmp1027;
  assign tmp1087 = s2 ? tmp1088 : tmp975;
  assign tmp1093 = l1 ? tmp31 : tmp116;
  assign tmp1092 = s0 ? tmp1093 : tmp975;
  assign tmp1094 = ~(l1 ? tmp17 : tmp173);
  assign tmp1091 = s1 ? tmp1092 : tmp1094;
  assign tmp1090 = s2 ? tmp1091 : tmp949;
  assign tmp1086 = s3 ? tmp1087 : tmp1090;
  assign tmp1075 = s4 ? tmp1076 : tmp1086;
  assign tmp1100 = l1 ? tmp17 : tmp783;
  assign tmp1099 = s0 ? tmp1100 : 0;
  assign tmp1098 = s1 ? tmp1099 : tmp1039;
  assign tmp1101 = ~(s1 ? tmp207 : tmp31);
  assign tmp1097 = s2 ? tmp1098 : tmp1101;
  assign tmp1103 = s1 ? tmp375 : tmp202;
  assign tmp1102 = ~(s2 ? 1 : tmp1103);
  assign tmp1096 = s3 ? tmp1097 : tmp1102;
  assign tmp1106 = l1 ? tmp26 : tmp116;
  assign tmp1105 = s2 ? tmp1042 : tmp1106;
  assign tmp1108 = ~(l1 ? tmp17 : tmp31);
  assign tmp1107 = s1 ? 1 : tmp1108;
  assign tmp1104 = ~(s3 ? tmp1105 : tmp1107);
  assign tmp1095 = ~(s4 ? tmp1096 : tmp1104);
  assign tmp1074 = s5 ? tmp1075 : tmp1095;
  assign tmp1049 = s6 ? tmp1050 : tmp1074;
  assign tmp1047 = s7 ? tmp1048 : tmp1049;
  assign tmp1109 = s6 ? tmp969 : tmp1003;
  assign tmp1046 = ~(s8 ? tmp1047 : tmp1109);
  assign tmp1044 = s9 ? tmp1045 : tmp1046;
  assign tmp888 = s10 ? tmp889 : tmp1044;
  assign tmp727 = s12 ? tmp728 : tmp888;
  assign tmp1119 = l1 ? tmp19 : tmp18;
  assign tmp1121 = l1 ? tmp19 : tmp185;
  assign tmp1123 = l2 ? 1 : tmp20;
  assign tmp1122 = ~(l1 ? tmp1123 : tmp45);
  assign tmp1120 = s0 ? tmp1121 : tmp1122;
  assign tmp1118 = s1 ? tmp1119 : tmp1120;
  assign tmp1128 = ~(l2 ? tmp17 : tmp20);
  assign tmp1127 = ~(l1 ? tmp897 : tmp1128);
  assign tmp1126 = s0 ? tmp322 : tmp1127;
  assign tmp1130 = l1 ? tmp322 : tmp117;
  assign tmp1129 = s0 ? tmp1130 : tmp1127;
  assign tmp1125 = s1 ? tmp1126 : tmp1129;
  assign tmp1132 = s0 ? tmp1130 : tmp31;
  assign tmp1134 = l1 ? tmp897 : tmp1128;
  assign tmp1135 = l1 ? tmp897 : tmp18;
  assign tmp1133 = ~(s0 ? tmp1134 : tmp1135);
  assign tmp1131 = s1 ? tmp1132 : tmp1133;
  assign tmp1124 = ~(s2 ? tmp1125 : tmp1131);
  assign tmp1117 = s3 ? tmp1118 : tmp1124;
  assign tmp1140 = l1 ? tmp322 : tmp45;
  assign tmp1139 = s0 ? tmp1140 : tmp322;
  assign tmp1141 = ~(s0 ? tmp1135 : tmp1134);
  assign tmp1138 = s1 ? tmp1139 : tmp1141;
  assign tmp1143 = s0 ? tmp1119 : 1;
  assign tmp1144 = l1 ? tmp19 : tmp33;
  assign tmp1142 = ~(s1 ? tmp1143 : tmp1144);
  assign tmp1137 = s2 ? tmp1138 : tmp1142;
  assign tmp1146 = s1 ? tmp1121 : 1;
  assign tmp1149 = l1 ? tmp927 : tmp1128;
  assign tmp1148 = s0 ? tmp1134 : tmp1149;
  assign tmp1151 = l1 ? tmp316 : 1;
  assign tmp1150 = s0 ? tmp1151 : tmp1134;
  assign tmp1147 = s1 ? tmp1148 : tmp1150;
  assign tmp1145 = ~(s2 ? tmp1146 : tmp1147);
  assign tmp1136 = ~(s3 ? tmp1137 : tmp1145);
  assign tmp1116 = s4 ? tmp1117 : tmp1136;
  assign tmp1158 = l1 ? tmp1123 : tmp45;
  assign tmp1157 = s0 ? tmp1158 : tmp31;
  assign tmp1156 = s1 ? tmp1157 : tmp322;
  assign tmp1160 = l1 ? tmp1123 : tmp780;
  assign tmp1161 = ~(s0 ? tmp1149 : tmp203);
  assign tmp1159 = s1 ? tmp1160 : tmp1161;
  assign tmp1155 = s2 ? tmp1156 : tmp1159;
  assign tmp1164 = ~(l1 ? tmp927 : tmp21);
  assign tmp1163 = s1 ? tmp1130 : tmp1164;
  assign tmp1166 = s0 ? tmp1151 : 1;
  assign tmp1168 = l1 ? tmp897 : tmp21;
  assign tmp1169 = l1 ? tmp927 : tmp21;
  assign tmp1167 = s0 ? tmp1168 : tmp1169;
  assign tmp1165 = ~(s1 ? tmp1166 : tmp1167);
  assign tmp1162 = s2 ? tmp1163 : tmp1165;
  assign tmp1154 = s3 ? tmp1155 : tmp1162;
  assign tmp1174 = l1 ? tmp897 : tmp164;
  assign tmp1173 = s0 ? 1 : tmp1174;
  assign tmp1175 = s0 ? tmp593 : tmp54;
  assign tmp1172 = s1 ? tmp1173 : tmp1175;
  assign tmp1176 = ~(l1 ? tmp322 : tmp780);
  assign tmp1171 = s2 ? tmp1172 : tmp1176;
  assign tmp1180 = l1 ? 1 : tmp780;
  assign tmp1181 = ~(l1 ? tmp19 : tmp26);
  assign tmp1179 = s0 ? tmp1180 : tmp1181;
  assign tmp1178 = s1 ? tmp1179 : tmp1164;
  assign tmp1177 = ~(s2 ? tmp1178 : 0);
  assign tmp1170 = ~(s3 ? tmp1171 : tmp1177);
  assign tmp1153 = s4 ? tmp1154 : tmp1170;
  assign tmp1186 = s0 ? tmp1169 : 1;
  assign tmp1185 = s1 ? tmp1186 : tmp94;
  assign tmp1184 = s2 ? tmp1185 : 0;
  assign tmp1188 = s1 ? 1 : tmp1039;
  assign tmp1187 = s2 ? 1 : tmp1188;
  assign tmp1183 = s3 ? tmp1184 : tmp1187;
  assign tmp1192 = ~(l1 ? tmp316 : 1);
  assign tmp1191 = s1 ? tmp174 : tmp1192;
  assign tmp1193 = l1 ? tmp966 : tmp780;
  assign tmp1190 = s2 ? tmp1191 : tmp1193;
  assign tmp1195 = ~(l1 ? tmp927 : tmp26);
  assign tmp1194 = s1 ? tmp174 : tmp1195;
  assign tmp1189 = ~(s3 ? tmp1190 : tmp1194);
  assign tmp1182 = ~(s4 ? tmp1183 : tmp1189);
  assign tmp1152 = ~(s5 ? tmp1153 : tmp1182);
  assign tmp1115 = ~(s6 ? tmp1116 : tmp1152);
  assign tmp1114 = s7 ? 1 : tmp1115;
  assign tmp1202 = l2 ? tmp780 : tmp19;
  assign tmp1203 = ~(l2 ? tmp780 : tmp20);
  assign tmp1201 = l1 ? tmp1202 : tmp1203;
  assign tmp1205 = l1 ? tmp74 : tmp811;
  assign tmp1206 = l1 ? tmp973 : tmp1203;
  assign tmp1204 = s0 ? tmp1205 : tmp1206;
  assign tmp1200 = s1 ? tmp1201 : tmp1204;
  assign tmp1210 = l1 ? tmp981 : tmp1128;
  assign tmp1209 = s0 ? tmp608 : tmp1210;
  assign tmp1213 = ~(l2 ? tmp780 : tmp33);
  assign tmp1212 = l1 ? tmp392 : tmp1213;
  assign tmp1211 = s0 ? tmp1212 : tmp1210;
  assign tmp1208 = s1 ? tmp1209 : tmp1211;
  assign tmp1215 = s0 ? tmp1212 : tmp375;
  assign tmp1217 = l1 ? tmp981 : tmp1203;
  assign tmp1216 = s0 ? tmp1210 : tmp1217;
  assign tmp1214 = s1 ? tmp1215 : tmp1216;
  assign tmp1207 = s2 ? tmp1208 : tmp1214;
  assign tmp1199 = s3 ? tmp1200 : tmp1207;
  assign tmp1222 = l1 ? tmp392 : tmp1203;
  assign tmp1221 = s0 ? tmp1222 : tmp603;
  assign tmp1223 = s0 ? tmp1217 : tmp1210;
  assign tmp1220 = s1 ? tmp1221 : tmp1223;
  assign tmp1225 = s0 ? tmp1201 : 1;
  assign tmp1226 = l1 ? tmp74 : tmp69;
  assign tmp1224 = s1 ? tmp1225 : tmp1226;
  assign tmp1219 = s2 ? tmp1220 : tmp1224;
  assign tmp1228 = s1 ? tmp1205 : 1;
  assign tmp1231 = l1 ? tmp1021 : tmp1128;
  assign tmp1230 = s0 ? tmp1210 : tmp1231;
  assign tmp1233 = l1 ? tmp316 : tmp21;
  assign tmp1232 = s0 ? tmp1233 : tmp1210;
  assign tmp1229 = s1 ? tmp1230 : tmp1232;
  assign tmp1227 = s2 ? tmp1228 : tmp1229;
  assign tmp1218 = s3 ? tmp1219 : tmp1227;
  assign tmp1198 = s4 ? tmp1199 : tmp1218;
  assign tmp1239 = s0 ? tmp1206 : tmp203;
  assign tmp1238 = s1 ? tmp1239 : tmp608;
  assign tmp1241 = l1 ? tmp973 : tmp69;
  assign tmp1242 = s0 ? tmp1231 : tmp375;
  assign tmp1240 = s1 ? tmp1241 : tmp1242;
  assign tmp1237 = s2 ? tmp1238 : tmp1240;
  assign tmp1244 = s1 ? tmp1212 : tmp1169;
  assign tmp1246 = s0 ? tmp1233 : 1;
  assign tmp1248 = l1 ? tmp981 : tmp21;
  assign tmp1249 = l1 ? tmp1021 : tmp21;
  assign tmp1247 = s0 ? tmp1248 : tmp1249;
  assign tmp1245 = s1 ? tmp1246 : tmp1247;
  assign tmp1243 = s2 ? tmp1244 : tmp1245;
  assign tmp1236 = s3 ? tmp1237 : tmp1243;
  assign tmp1254 = l1 ? tmp981 : tmp840;
  assign tmp1253 = s0 ? 1 : tmp1254;
  assign tmp1255 = s0 ? tmp618 : tmp97;
  assign tmp1252 = s1 ? tmp1253 : tmp1255;
  assign tmp1256 = l1 ? tmp392 : tmp69;
  assign tmp1251 = s2 ? tmp1252 : tmp1256;
  assign tmp1260 = ~(l1 ? tmp1202 : tmp21);
  assign tmp1259 = s0 ? tmp1180 : tmp1260;
  assign tmp1258 = s1 ? tmp1259 : tmp1164;
  assign tmp1257 = ~(s2 ? tmp1258 : 0);
  assign tmp1250 = s3 ? tmp1251 : tmp1257;
  assign tmp1235 = s4 ? tmp1236 : tmp1250;
  assign tmp1265 = ~(l1 ? tmp31 : tmp17);
  assign tmp1264 = s1 ? tmp1186 : tmp1265;
  assign tmp1263 = s2 ? tmp1264 : 0;
  assign tmp1262 = s3 ? tmp1263 : tmp1187;
  assign tmp1269 = ~(l1 ? tmp316 : tmp21);
  assign tmp1268 = s1 ? tmp174 : tmp1269;
  assign tmp1267 = s2 ? tmp1268 : tmp1193;
  assign tmp1266 = ~(s3 ? tmp1267 : tmp1194);
  assign tmp1261 = s4 ? tmp1262 : tmp1266;
  assign tmp1234 = s5 ? tmp1235 : tmp1261;
  assign tmp1197 = ~(s6 ? tmp1198 : tmp1234);
  assign tmp1196 = s7 ? 1 : tmp1197;
  assign tmp1113 = s8 ? tmp1114 : tmp1196;
  assign tmp1276 = l1 ? tmp1202 : tmp185;
  assign tmp1278 = l1 ? tmp973 : tmp185;
  assign tmp1277 = s0 ? tmp224 : tmp1278;
  assign tmp1275 = s1 ? tmp1276 : tmp1277;
  assign tmp1282 = l2 ? tmp898 : tmp33;
  assign tmp1283 = ~(l1 ? tmp981 : tmp193);
  assign tmp1281 = s0 ? tmp1282 : tmp1283;
  assign tmp1285 = l1 ? tmp392 : tmp185;
  assign tmp1286 = l1 ? tmp981 : tmp193;
  assign tmp1284 = ~(s0 ? tmp1285 : tmp1286);
  assign tmp1280 = s1 ? tmp1281 : tmp1284;
  assign tmp1288 = s0 ? tmp1285 : tmp185;
  assign tmp1290 = l1 ? tmp981 : tmp185;
  assign tmp1289 = s0 ? tmp1286 : tmp1290;
  assign tmp1287 = ~(s1 ? tmp1288 : tmp1289);
  assign tmp1279 = ~(s2 ? tmp1280 : tmp1287);
  assign tmp1274 = s3 ? tmp1275 : tmp1279;
  assign tmp1294 = s0 ? tmp1285 : tmp603;
  assign tmp1295 = s0 ? tmp1290 : tmp1286;
  assign tmp1293 = s1 ? tmp1294 : tmp1295;
  assign tmp1297 = s0 ? tmp1276 : 1;
  assign tmp1298 = l1 ? tmp74 : tmp33;
  assign tmp1296 = s1 ? tmp1297 : tmp1298;
  assign tmp1292 = s2 ? tmp1293 : tmp1296;
  assign tmp1300 = s1 ? tmp224 : 1;
  assign tmp1303 = l1 ? tmp1021 : tmp193;
  assign tmp1302 = s0 ? tmp1286 : tmp1303;
  assign tmp1304 = s0 ? tmp1151 : tmp1286;
  assign tmp1301 = s1 ? tmp1302 : tmp1304;
  assign tmp1299 = s2 ? tmp1300 : tmp1301;
  assign tmp1291 = s3 ? tmp1292 : tmp1299;
  assign tmp1273 = s4 ? tmp1274 : tmp1291;
  assign tmp1310 = s0 ? tmp1278 : tmp203;
  assign tmp1311 = ~(l2 ? tmp898 : tmp33);
  assign tmp1309 = s1 ? tmp1310 : tmp1311;
  assign tmp1313 = s0 ? tmp1303 : tmp221;
  assign tmp1312 = s1 ? tmp1278 : tmp1313;
  assign tmp1308 = s2 ? tmp1309 : tmp1312;
  assign tmp1316 = l1 ? tmp927 : tmp193;
  assign tmp1315 = s1 ? tmp1285 : tmp1316;
  assign tmp1319 = l1 ? tmp1021 : 1;
  assign tmp1318 = s0 ? tmp1286 : tmp1319;
  assign tmp1317 = s1 ? tmp1166 : tmp1318;
  assign tmp1314 = s2 ? tmp1315 : tmp1317;
  assign tmp1307 = s3 ? tmp1308 : tmp1314;
  assign tmp1323 = s0 ? 1 : tmp1290;
  assign tmp1324 = s0 ? tmp618 : tmp207;
  assign tmp1322 = s1 ? tmp1323 : tmp1324;
  assign tmp1321 = s2 ? tmp1322 : tmp1285;
  assign tmp1328 = ~(l1 ? tmp1202 : 1);
  assign tmp1327 = s0 ? tmp23 : tmp1328;
  assign tmp1329 = ~(l1 ? tmp927 : 1);
  assign tmp1326 = s1 ? tmp1327 : tmp1329;
  assign tmp1325 = ~(s2 ? tmp1326 : 0);
  assign tmp1320 = s3 ? tmp1321 : tmp1325;
  assign tmp1306 = s4 ? tmp1307 : tmp1320;
  assign tmp1334 = s0 ? tmp1316 : 1;
  assign tmp1333 = s1 ? tmp1334 : tmp94;
  assign tmp1335 = ~(s1 ? tmp135 : 1);
  assign tmp1332 = s2 ? tmp1333 : tmp1335;
  assign tmp1337 = s1 ? 1 : tmp54;
  assign tmp1336 = s2 ? 1 : tmp1337;
  assign tmp1331 = s3 ? tmp1332 : tmp1336;
  assign tmp1340 = l1 ? tmp966 : tmp24;
  assign tmp1339 = s2 ? tmp1191 : tmp1340;
  assign tmp1341 = s1 ? tmp174 : tmp1329;
  assign tmp1338 = ~(s3 ? tmp1339 : tmp1341);
  assign tmp1330 = s4 ? tmp1331 : tmp1338;
  assign tmp1305 = s5 ? tmp1306 : tmp1330;
  assign tmp1272 = ~(s6 ? tmp1273 : tmp1305);
  assign tmp1271 = s7 ? 1 : tmp1272;
  assign tmp1270 = s8 ? tmp1196 : tmp1271;
  assign tmp1112 = s9 ? tmp1113 : tmp1270;
  assign tmp1349 = l1 ? tmp1202 : tmp18;
  assign tmp1351 = l1 ? tmp973 : tmp18;
  assign tmp1350 = s0 ? tmp224 : tmp1351;
  assign tmp1348 = s1 ? tmp1349 : tmp1350;
  assign tmp1355 = ~(l1 ? tmp981 : tmp264);
  assign tmp1354 = s0 ? tmp1282 : tmp1355;
  assign tmp1357 = l1 ? tmp392 : tmp38;
  assign tmp1358 = l1 ? tmp981 : tmp264;
  assign tmp1356 = ~(s0 ? tmp1357 : tmp1358);
  assign tmp1353 = s1 ? tmp1354 : tmp1356;
  assign tmp1360 = s0 ? tmp1357 : tmp185;
  assign tmp1362 = l1 ? tmp981 : tmp18;
  assign tmp1361 = s0 ? tmp1358 : tmp1362;
  assign tmp1359 = ~(s1 ? tmp1360 : tmp1361);
  assign tmp1352 = ~(s2 ? tmp1353 : tmp1359);
  assign tmp1347 = s3 ? tmp1348 : tmp1352;
  assign tmp1367 = l1 ? tmp392 : tmp18;
  assign tmp1366 = s0 ? tmp1367 : tmp603;
  assign tmp1368 = s0 ? tmp1362 : tmp1358;
  assign tmp1365 = s1 ? tmp1366 : tmp1368;
  assign tmp1370 = s0 ? tmp1349 : 1;
  assign tmp1369 = s1 ? tmp1370 : tmp1298;
  assign tmp1364 = s2 ? tmp1365 : tmp1369;
  assign tmp1374 = l1 ? tmp1021 : tmp264;
  assign tmp1373 = s0 ? tmp1358 : tmp1374;
  assign tmp1375 = s0 ? tmp1151 : tmp1358;
  assign tmp1372 = s1 ? tmp1373 : tmp1375;
  assign tmp1371 = s2 ? tmp1300 : tmp1372;
  assign tmp1363 = s3 ? tmp1364 : tmp1371;
  assign tmp1346 = s4 ? tmp1347 : tmp1363;
  assign tmp1381 = s0 ? tmp1351 : tmp203;
  assign tmp1380 = s1 ? tmp1381 : tmp1311;
  assign tmp1383 = l1 ? tmp973 : tmp164;
  assign tmp1384 = s0 ? tmp1374 : tmp221;
  assign tmp1382 = s1 ? tmp1383 : tmp1384;
  assign tmp1379 = s2 ? tmp1380 : tmp1382;
  assign tmp1387 = l1 ? tmp927 : tmp228;
  assign tmp1386 = s1 ? tmp1357 : tmp1387;
  assign tmp1390 = l1 ? tmp981 : tmp228;
  assign tmp1391 = l1 ? tmp1021 : tmp26;
  assign tmp1389 = s0 ? tmp1390 : tmp1391;
  assign tmp1388 = s1 ? tmp1166 : tmp1389;
  assign tmp1385 = s2 ? tmp1386 : tmp1388;
  assign tmp1378 = s3 ? tmp1379 : tmp1385;
  assign tmp1396 = l1 ? tmp981 : tmp164;
  assign tmp1395 = s0 ? 1 : tmp1396;
  assign tmp1394 = s1 ? tmp1395 : tmp1324;
  assign tmp1397 = l1 ? tmp392 : tmp164;
  assign tmp1393 = s2 ? tmp1394 : tmp1397;
  assign tmp1401 = l1 ? 1 : tmp81;
  assign tmp1402 = ~(l1 ? tmp1202 : tmp26);
  assign tmp1400 = s0 ? tmp1401 : tmp1402;
  assign tmp1399 = s1 ? tmp1400 : tmp1164;
  assign tmp1398 = ~(s2 ? tmp1399 : 0);
  assign tmp1392 = s3 ? tmp1393 : tmp1398;
  assign tmp1377 = s4 ? tmp1378 : tmp1392;
  assign tmp1407 = s0 ? tmp1387 : 1;
  assign tmp1406 = s1 ? tmp1407 : tmp94;
  assign tmp1408 = ~(s1 ? tmp397 : 1);
  assign tmp1405 = s2 ? tmp1406 : tmp1408;
  assign tmp1404 = s3 ? tmp1405 : tmp1187;
  assign tmp1411 = l1 ? tmp966 : tmp81;
  assign tmp1410 = s2 ? tmp1191 : tmp1411;
  assign tmp1409 = ~(s3 ? tmp1410 : tmp1194);
  assign tmp1403 = s4 ? tmp1404 : tmp1409;
  assign tmp1376 = s5 ? tmp1377 : tmp1403;
  assign tmp1345 = ~(s6 ? tmp1346 : tmp1376);
  assign tmp1344 = s7 ? 1 : tmp1345;
  assign tmp1343 = s8 ? tmp1344 : 1;
  assign tmp1414 = s6 ? tmp1116 : tmp1152;
  assign tmp1415 = s6 ? tmp1273 : tmp1305;
  assign tmp1413 = s7 ? tmp1414 : tmp1415;
  assign tmp1417 = s6 ? tmp1198 : tmp1234;
  assign tmp1418 = s6 ? tmp1346 : tmp1376;
  assign tmp1416 = s7 ? tmp1417 : tmp1418;
  assign tmp1412 = ~(s8 ? tmp1413 : tmp1416);
  assign tmp1342 = s9 ? tmp1343 : tmp1412;
  assign tmp1111 = s10 ? tmp1112 : tmp1342;
  assign tmp1427 = l1 ? tmp19 : tmp901;
  assign tmp1429 = ~(l1 ? tmp1123 : tmp20);
  assign tmp1428 = s0 ? tmp363 : tmp1429;
  assign tmp1426 = s1 ? tmp1427 : tmp1428;
  assign tmp1433 = ~(l1 ? tmp897 : tmp898);
  assign tmp1432 = s0 ? tmp336 : tmp1433;
  assign tmp1434 = s0 ? tmp321 : tmp1433;
  assign tmp1431 = s1 ? tmp1432 : tmp1434;
  assign tmp1436 = s0 ? tmp321 : 0;
  assign tmp1438 = l1 ? tmp897 : tmp898;
  assign tmp1439 = l1 ? tmp897 : tmp901;
  assign tmp1437 = ~(s0 ? tmp1438 : tmp1439);
  assign tmp1435 = s1 ? tmp1436 : tmp1437;
  assign tmp1430 = ~(s2 ? tmp1431 : tmp1435);
  assign tmp1425 = s3 ? tmp1426 : tmp1430;
  assign tmp1444 = l1 ? tmp322 : tmp20;
  assign tmp1443 = s0 ? tmp1444 : tmp337;
  assign tmp1445 = ~(s0 ? tmp1439 : tmp1438);
  assign tmp1442 = s1 ? tmp1443 : tmp1445;
  assign tmp1447 = s0 ? tmp1427 : 1;
  assign tmp1446 = ~(s1 ? tmp1447 : tmp363);
  assign tmp1441 = s2 ? tmp1442 : tmp1446;
  assign tmp1449 = s1 ? tmp363 : 1;
  assign tmp1452 = l1 ? tmp927 : tmp898;
  assign tmp1451 = s0 ? tmp1438 : tmp1452;
  assign tmp1453 = s0 ? tmp1151 : tmp1438;
  assign tmp1450 = s1 ? tmp1451 : tmp1453;
  assign tmp1448 = ~(s2 ? tmp1449 : tmp1450);
  assign tmp1440 = ~(s3 ? tmp1441 : tmp1448);
  assign tmp1424 = s4 ? tmp1425 : tmp1440;
  assign tmp1460 = l1 ? tmp1123 : tmp20;
  assign tmp1459 = s0 ? tmp1460 : 0;
  assign tmp1458 = s1 ? tmp1459 : tmp336;
  assign tmp1462 = l1 ? tmp1123 : tmp102;
  assign tmp1463 = ~(s0 ? tmp1452 : 1);
  assign tmp1461 = s1 ? tmp1462 : tmp1463;
  assign tmp1457 = s2 ? tmp1458 : tmp1461;
  assign tmp1465 = s1 ? tmp321 : tmp1195;
  assign tmp1468 = l1 ? tmp897 : tmp26;
  assign tmp1467 = s0 ? tmp1468 : tmp1169;
  assign tmp1466 = ~(s1 ? tmp1166 : tmp1467);
  assign tmp1464 = s2 ? tmp1465 : tmp1466;
  assign tmp1456 = s3 ? tmp1457 : tmp1464;
  assign tmp1472 = s0 ? 1 : tmp1468;
  assign tmp1473 = s0 ? tmp363 : tmp54;
  assign tmp1471 = s1 ? tmp1472 : tmp1473;
  assign tmp1474 = ~(l1 ? tmp322 : tmp102);
  assign tmp1470 = s2 ? tmp1471 : tmp1474;
  assign tmp1478 = l1 ? 1 : tmp102;
  assign tmp1477 = s0 ? tmp1478 : tmp1181;
  assign tmp1476 = s1 ? tmp1477 : tmp1164;
  assign tmp1475 = ~(s2 ? tmp1476 : 0);
  assign tmp1469 = ~(s3 ? tmp1470 : tmp1475);
  assign tmp1455 = s4 ? tmp1456 : tmp1469;
  assign tmp1484 = l1 ? tmp927 : tmp26;
  assign tmp1483 = s0 ? tmp1484 : 1;
  assign tmp1482 = s1 ? tmp1483 : tmp94;
  assign tmp1481 = s2 ? tmp1482 : tmp374;
  assign tmp1480 = s3 ? tmp1481 : tmp1187;
  assign tmp1487 = l1 ? tmp966 : tmp102;
  assign tmp1486 = s2 ? tmp1191 : tmp1487;
  assign tmp1485 = ~(s3 ? tmp1486 : tmp1194);
  assign tmp1479 = ~(s4 ? tmp1480 : tmp1485);
  assign tmp1454 = ~(s5 ? tmp1455 : tmp1479);
  assign tmp1423 = ~(s6 ? tmp1424 : tmp1454);
  assign tmp1422 = s7 ? 1 : tmp1423;
  assign tmp1493 = l1 ? tmp1202 : tmp898;
  assign tmp1496 = l2 ? tmp898 : 1;
  assign tmp1495 = l1 ? tmp74 : tmp1496;
  assign tmp1497 = l1 ? tmp973 : tmp898;
  assign tmp1494 = s0 ? tmp1495 : tmp1497;
  assign tmp1492 = s1 ? tmp1493 : tmp1494;
  assign tmp1501 = l1 ? tmp981 : tmp898;
  assign tmp1500 = s0 ? tmp391 : tmp1501;
  assign tmp1504 = l2 ? tmp898 : tmp19;
  assign tmp1503 = l1 ? tmp392 : tmp1504;
  assign tmp1502 = s0 ? tmp1503 : tmp1501;
  assign tmp1499 = s1 ? tmp1500 : tmp1502;
  assign tmp1506 = s0 ? tmp1503 : tmp135;
  assign tmp1505 = s1 ? tmp1506 : tmp1501;
  assign tmp1498 = s2 ? tmp1499 : tmp1505;
  assign tmp1491 = s3 ? tmp1492 : tmp1498;
  assign tmp1511 = l1 ? tmp392 : tmp898;
  assign tmp1510 = s0 ? tmp1511 : tmp237;
  assign tmp1509 = s1 ? tmp1510 : tmp1501;
  assign tmp1513 = s0 ? tmp1493 : 1;
  assign tmp1514 = l1 ? tmp74 : tmp898;
  assign tmp1512 = s1 ? tmp1513 : tmp1514;
  assign tmp1508 = s2 ? tmp1509 : tmp1512;
  assign tmp1516 = s1 ? tmp1495 : 1;
  assign tmp1519 = l1 ? tmp1021 : tmp898;
  assign tmp1518 = s0 ? tmp1501 : tmp1519;
  assign tmp1520 = s0 ? tmp1233 : tmp1501;
  assign tmp1517 = s1 ? tmp1518 : tmp1520;
  assign tmp1515 = s2 ? tmp1516 : tmp1517;
  assign tmp1507 = s3 ? tmp1508 : tmp1515;
  assign tmp1490 = s4 ? tmp1491 : tmp1507;
  assign tmp1526 = s0 ? tmp1497 : 1;
  assign tmp1525 = s1 ? tmp1526 : tmp391;
  assign tmp1529 = l2 ? tmp898 : tmp21;
  assign tmp1528 = l1 ? tmp973 : tmp1529;
  assign tmp1530 = s0 ? tmp1519 : tmp135;
  assign tmp1527 = s1 ? tmp1528 : tmp1530;
  assign tmp1524 = s2 ? tmp1525 : tmp1527;
  assign tmp1533 = l1 ? tmp927 : tmp1529;
  assign tmp1532 = s1 ? tmp1503 : tmp1533;
  assign tmp1536 = l1 ? tmp981 : tmp1529;
  assign tmp1535 = s0 ? tmp1536 : tmp1249;
  assign tmp1534 = s1 ? tmp1246 : tmp1535;
  assign tmp1531 = s2 ? tmp1532 : tmp1534;
  assign tmp1523 = s3 ? tmp1524 : tmp1531;
  assign tmp1540 = s0 ? 1 : tmp1536;
  assign tmp1541 = s0 ? tmp237 : tmp97;
  assign tmp1539 = s1 ? tmp1540 : tmp1541;
  assign tmp1542 = l1 ? tmp392 : tmp1529;
  assign tmp1538 = s2 ? tmp1539 : tmp1542;
  assign tmp1547 = ~(l2 ? tmp898 : tmp21);
  assign tmp1546 = l1 ? 1 : tmp1547;
  assign tmp1545 = s0 ? tmp1546 : tmp1260;
  assign tmp1544 = s1 ? tmp1545 : tmp1164;
  assign tmp1543 = ~(s2 ? tmp1544 : 0);
  assign tmp1537 = s3 ? tmp1538 : tmp1543;
  assign tmp1522 = s4 ? tmp1523 : tmp1537;
  assign tmp1552 = s0 ? tmp1533 : 1;
  assign tmp1551 = s1 ? tmp1552 : tmp1265;
  assign tmp1553 = ~(s1 ? tmp221 : 1);
  assign tmp1550 = s2 ? tmp1551 : tmp1553;
  assign tmp1549 = s3 ? tmp1550 : tmp1187;
  assign tmp1556 = l1 ? tmp966 : tmp1547;
  assign tmp1555 = s2 ? tmp1268 : tmp1556;
  assign tmp1554 = ~(s3 ? tmp1555 : tmp1194);
  assign tmp1548 = s4 ? tmp1549 : tmp1554;
  assign tmp1521 = s5 ? tmp1522 : tmp1548;
  assign tmp1489 = ~(s6 ? tmp1490 : tmp1521);
  assign tmp1488 = s7 ? 1 : tmp1489;
  assign tmp1421 = s8 ? tmp1422 : tmp1488;
  assign tmp1563 = l1 ? tmp1202 : 1;
  assign tmp1565 = l1 ? tmp973 : 1;
  assign tmp1564 = s0 ? tmp237 : tmp1565;
  assign tmp1562 = s1 ? tmp1563 : tmp1564;
  assign tmp1568 = l1 ? tmp392 : 1;
  assign tmp1569 = l1 ? tmp981 : 1;
  assign tmp1567 = s0 ? tmp1568 : tmp1569;
  assign tmp1571 = s0 ? tmp1568 : 1;
  assign tmp1570 = s1 ? tmp1571 : tmp1569;
  assign tmp1566 = s2 ? tmp1567 : tmp1570;
  assign tmp1561 = s3 ? tmp1562 : tmp1566;
  assign tmp1575 = s0 ? tmp1568 : tmp237;
  assign tmp1574 = s1 ? tmp1575 : tmp1569;
  assign tmp1577 = s0 ? tmp1563 : 1;
  assign tmp1576 = s1 ? tmp1577 : tmp237;
  assign tmp1573 = s2 ? tmp1574 : tmp1576;
  assign tmp1579 = s1 ? tmp237 : 1;
  assign tmp1581 = s0 ? tmp1569 : tmp1319;
  assign tmp1582 = s0 ? tmp1151 : tmp1569;
  assign tmp1580 = s1 ? tmp1581 : tmp1582;
  assign tmp1578 = s2 ? tmp1579 : tmp1580;
  assign tmp1572 = s3 ? tmp1573 : tmp1578;
  assign tmp1560 = s4 ? tmp1561 : tmp1572;
  assign tmp1588 = s0 ? tmp1565 : 1;
  assign tmp1587 = s1 ? tmp1588 : tmp1568;
  assign tmp1590 = s0 ? tmp1319 : 1;
  assign tmp1589 = s1 ? tmp1565 : tmp1590;
  assign tmp1586 = s2 ? tmp1587 : tmp1589;
  assign tmp1593 = l1 ? tmp927 : 1;
  assign tmp1592 = s1 ? tmp1568 : tmp1593;
  assign tmp1594 = s1 ? tmp1166 : tmp1581;
  assign tmp1591 = s2 ? tmp1592 : tmp1594;
  assign tmp1585 = s3 ? tmp1586 : tmp1591;
  assign tmp1598 = s0 ? 1 : tmp1569;
  assign tmp1599 = s0 ? tmp237 : tmp207;
  assign tmp1597 = s1 ? tmp1598 : tmp1599;
  assign tmp1596 = s2 ? tmp1597 : tmp1568;
  assign tmp1602 = s0 ? tmp83 : tmp1328;
  assign tmp1601 = s1 ? tmp1602 : tmp1329;
  assign tmp1600 = ~(s2 ? tmp1601 : 0);
  assign tmp1595 = s3 ? tmp1596 : tmp1600;
  assign tmp1584 = s4 ? tmp1585 : tmp1595;
  assign tmp1607 = s0 ? tmp1593 : 1;
  assign tmp1606 = s1 ? tmp1607 : tmp94;
  assign tmp1608 = ~(s1 ? tmp83 : 1);
  assign tmp1605 = s2 ? tmp1606 : tmp1608;
  assign tmp1604 = s3 ? tmp1605 : tmp1336;
  assign tmp1611 = l1 ? tmp966 : 0;
  assign tmp1610 = s2 ? tmp1191 : tmp1611;
  assign tmp1609 = ~(s3 ? tmp1610 : tmp1341);
  assign tmp1603 = s4 ? tmp1604 : tmp1609;
  assign tmp1583 = s5 ? tmp1584 : tmp1603;
  assign tmp1559 = ~(s6 ? tmp1560 : tmp1583);
  assign tmp1558 = s7 ? 1 : tmp1559;
  assign tmp1557 = s8 ? tmp1488 : tmp1558;
  assign tmp1420 = s9 ? tmp1421 : tmp1557;
  assign tmp1619 = l1 ? tmp1202 : tmp901;
  assign tmp1621 = l1 ? tmp973 : tmp901;
  assign tmp1620 = s0 ? tmp237 : tmp1621;
  assign tmp1618 = s1 ? tmp1619 : tmp1620;
  assign tmp1624 = l1 ? tmp392 : tmp74;
  assign tmp1625 = l1 ? tmp981 : tmp901;
  assign tmp1623 = s0 ? tmp1624 : tmp1625;
  assign tmp1627 = s0 ? tmp1624 : 1;
  assign tmp1626 = s1 ? tmp1627 : tmp1625;
  assign tmp1622 = s2 ? tmp1623 : tmp1626;
  assign tmp1617 = s3 ? tmp1618 : tmp1622;
  assign tmp1632 = l1 ? tmp392 : tmp901;
  assign tmp1631 = s0 ? tmp1632 : tmp237;
  assign tmp1630 = s1 ? tmp1631 : tmp1625;
  assign tmp1634 = s0 ? tmp1619 : 1;
  assign tmp1633 = s1 ? tmp1634 : tmp237;
  assign tmp1629 = s2 ? tmp1630 : tmp1633;
  assign tmp1638 = l1 ? tmp1021 : tmp901;
  assign tmp1637 = s0 ? tmp1625 : tmp1638;
  assign tmp1639 = s0 ? tmp1151 : tmp1625;
  assign tmp1636 = s1 ? tmp1637 : tmp1639;
  assign tmp1635 = s2 ? tmp1579 : tmp1636;
  assign tmp1628 = s3 ? tmp1629 : tmp1635;
  assign tmp1616 = s4 ? tmp1617 : tmp1628;
  assign tmp1645 = s0 ? tmp1621 : 1;
  assign tmp1644 = s1 ? tmp1645 : tmp1624;
  assign tmp1647 = l1 ? tmp973 : tmp26;
  assign tmp1648 = s0 ? tmp1638 : 1;
  assign tmp1646 = s1 ? tmp1647 : tmp1648;
  assign tmp1643 = s2 ? tmp1644 : tmp1646;
  assign tmp1650 = s1 ? tmp1624 : tmp1484;
  assign tmp1653 = l1 ? tmp981 : tmp26;
  assign tmp1652 = s0 ? tmp1653 : tmp1391;
  assign tmp1651 = s1 ? tmp1166 : tmp1652;
  assign tmp1649 = s2 ? tmp1650 : tmp1651;
  assign tmp1642 = s3 ? tmp1643 : tmp1649;
  assign tmp1657 = s0 ? 1 : tmp1653;
  assign tmp1656 = s1 ? tmp1657 : tmp1599;
  assign tmp1658 = l1 ? tmp392 : tmp26;
  assign tmp1655 = s2 ? tmp1656 : tmp1658;
  assign tmp1661 = s0 ? tmp1478 : tmp1402;
  assign tmp1660 = s1 ? tmp1661 : tmp1164;
  assign tmp1659 = ~(s2 ? tmp1660 : 0);
  assign tmp1654 = s3 ? tmp1655 : tmp1659;
  assign tmp1641 = s4 ? tmp1642 : tmp1654;
  assign tmp1662 = s4 ? tmp1480 : tmp1485;
  assign tmp1640 = s5 ? tmp1641 : tmp1662;
  assign tmp1615 = ~(s6 ? tmp1616 : tmp1640);
  assign tmp1614 = s7 ? 1 : tmp1615;
  assign tmp1613 = s8 ? tmp1614 : 1;
  assign tmp1665 = s6 ? tmp1424 : tmp1454;
  assign tmp1666 = s6 ? tmp1560 : tmp1583;
  assign tmp1664 = s7 ? tmp1665 : tmp1666;
  assign tmp1668 = s6 ? tmp1490 : tmp1521;
  assign tmp1669 = s6 ? tmp1616 : tmp1640;
  assign tmp1667 = s7 ? tmp1668 : tmp1669;
  assign tmp1663 = ~(s8 ? tmp1664 : tmp1667);
  assign tmp1612 = s9 ? tmp1613 : tmp1663;
  assign tmp1419 = s10 ? tmp1420 : tmp1612;
  assign tmp1110 = s12 ? tmp1111 : tmp1419;
  assign tmp726 = s13 ? tmp727 : tmp1110;
  assign tmp4 = s14 ? tmp5 : tmp726;
  assign tmp1681 = l1 ? tmp927 : 0;
  assign tmp1684 = l2 ? 1 : tmp110;
  assign tmp1683 = l1 ? tmp1684 : 1;
  assign tmp1682 = ~(s0 ? 1 : tmp1683);
  assign tmp1680 = s1 ? tmp1681 : tmp1682;
  assign tmp1689 = l2 ? tmp19 : tmp16;
  assign tmp1690 = ~(l2 ? tmp110 : 1);
  assign tmp1688 = ~(l1 ? tmp1689 : tmp1690);
  assign tmp1687 = s0 ? 1 : tmp1688;
  assign tmp1692 = l1 ? tmp966 : 1;
  assign tmp1691 = s0 ? tmp1692 : tmp1688;
  assign tmp1686 = s1 ? tmp1687 : tmp1691;
  assign tmp1694 = s0 ? tmp1692 : 1;
  assign tmp1693 = s1 ? tmp1694 : tmp1688;
  assign tmp1685 = ~(s2 ? tmp1686 : tmp1693);
  assign tmp1679 = s3 ? tmp1680 : tmp1685;
  assign tmp1697 = s1 ? 1 : tmp1688;
  assign tmp1699 = s0 ? tmp1681 : 0;
  assign tmp1698 = ~(s1 ? tmp1699 : 0);
  assign tmp1696 = s2 ? tmp1697 : tmp1698;
  assign tmp1702 = ~(l1 ? tmp74 : tmp24);
  assign tmp1701 = s1 ? 1 : tmp1702;
  assign tmp1705 = l1 ? tmp1689 : tmp1690;
  assign tmp1706 = l1 ? tmp19 : tmp1690;
  assign tmp1704 = s0 ? tmp1705 : tmp1706;
  assign tmp1708 = l1 ? tmp19 : tmp24;
  assign tmp1707 = s0 ? tmp1708 : tmp1705;
  assign tmp1703 = ~(s1 ? tmp1704 : tmp1707);
  assign tmp1700 = s2 ? tmp1701 : tmp1703;
  assign tmp1695 = ~(s3 ? tmp1696 : tmp1700);
  assign tmp1678 = s4 ? tmp1679 : tmp1695;
  assign tmp1714 = s0 ? tmp1683 : 1;
  assign tmp1713 = s1 ? tmp1714 : 1;
  assign tmp1716 = ~(s0 ? tmp1706 : 0);
  assign tmp1715 = s1 ? tmp1683 : tmp1716;
  assign tmp1712 = s2 ? tmp1713 : tmp1715;
  assign tmp1719 = ~(l1 ? tmp19 : tmp1690);
  assign tmp1718 = s1 ? tmp594 : tmp1719;
  assign tmp1722 = l1 ? tmp74 : tmp31;
  assign tmp1721 = s0 ? tmp1708 : tmp1722;
  assign tmp1723 = s0 ? tmp1705 : tmp1708;
  assign tmp1720 = ~(s1 ? tmp1721 : tmp1723);
  assign tmp1717 = s2 ? tmp1718 : tmp1720;
  assign tmp1711 = s3 ? tmp1712 : tmp1717;
  assign tmp1728 = l1 ? tmp1689 : 0;
  assign tmp1727 = s0 ? tmp23 : tmp1728;
  assign tmp1726 = s1 ? tmp1727 : 0;
  assign tmp1725 = s2 ? tmp1726 : 0;
  assign tmp1731 = s0 ? 1 : tmp569;
  assign tmp1732 = ~(l1 ? tmp19 : tmp24);
  assign tmp1730 = s1 ? tmp1731 : tmp1732;
  assign tmp1734 = l1 ? tmp74 : tmp24;
  assign tmp1733 = ~(s1 ? tmp131 : tmp1734);
  assign tmp1729 = ~(s2 ? tmp1730 : tmp1733);
  assign tmp1724 = ~(s3 ? tmp1725 : tmp1729);
  assign tmp1710 = s4 ? tmp1711 : tmp1724;
  assign tmp1739 = s0 ? tmp1706 : 1;
  assign tmp1738 = s1 ? tmp1739 : tmp203;
  assign tmp1737 = s2 ? tmp1738 : 0;
  assign tmp1742 = ~(l1 ? tmp19 : tmp31);
  assign tmp1741 = s1 ? 1 : tmp1742;
  assign tmp1743 = ~(s1 ? tmp83 : 0);
  assign tmp1740 = ~(s2 ? tmp1741 : tmp1743);
  assign tmp1736 = s3 ? tmp1737 : tmp1740;
  assign tmp1746 = s1 ? tmp593 : tmp1708;
  assign tmp1747 = ~(l1 ? tmp322 : 1);
  assign tmp1745 = s2 ? tmp1746 : tmp1747;
  assign tmp1749 = l1 ? tmp19 : tmp31;
  assign tmp1748 = s1 ? tmp1749 : tmp593;
  assign tmp1744 = s3 ? tmp1745 : tmp1748;
  assign tmp1735 = ~(s4 ? tmp1736 : tmp1744);
  assign tmp1709 = ~(s5 ? tmp1710 : tmp1735);
  assign tmp1677 = s6 ? tmp1678 : tmp1709;
  assign tmp1676 = s7 ? 1 : tmp1677;
  assign tmp1757 = ~(l1 ? tmp31 : 1);
  assign tmp1756 = s1 ? tmp1739 : tmp1757;
  assign tmp1755 = s2 ? tmp1756 : 0;
  assign tmp1754 = s3 ? tmp1755 : tmp1740;
  assign tmp1753 = ~(s4 ? tmp1754 : tmp1744);
  assign tmp1752 = ~(s5 ? tmp1710 : tmp1753);
  assign tmp1751 = s6 ? tmp1678 : tmp1752;
  assign tmp1750 = s7 ? 1 : tmp1751;
  assign tmp1675 = s8 ? tmp1676 : tmp1750;
  assign tmp1674 = s9 ? tmp1675 : tmp1750;
  assign tmp1759 = s8 ? tmp1750 : 1;
  assign tmp1761 = s7 ? tmp1677 : tmp1751;
  assign tmp1760 = s8 ? tmp1761 : tmp1751;
  assign tmp1758 = s9 ? tmp1759 : tmp1760;
  assign tmp1673 = s10 ? tmp1674 : tmp1758;
  assign tmp1771 = ~(l2 ? 1 : tmp110);
  assign tmp1770 = l1 ? tmp24 : tmp1771;
  assign tmp1769 = s1 ? tmp1770 : 0;
  assign tmp1774 = ~(l1 ? tmp24 : tmp16);
  assign tmp1773 = s0 ? 1 : tmp1774;
  assign tmp1775 = s1 ? 1 : tmp1774;
  assign tmp1772 = ~(s2 ? tmp1773 : tmp1775);
  assign tmp1768 = s3 ? tmp1769 : tmp1772;
  assign tmp1779 = s0 ? tmp1770 : 0;
  assign tmp1778 = ~(s1 ? tmp1779 : 0);
  assign tmp1777 = s2 ? tmp1775 : tmp1778;
  assign tmp1782 = ~(l1 ? tmp31 : tmp19);
  assign tmp1781 = s1 ? 1 : tmp1782;
  assign tmp1784 = l1 ? tmp24 : tmp16;
  assign tmp1786 = l1 ? tmp24 : tmp19;
  assign tmp1785 = s0 ? tmp1786 : tmp1784;
  assign tmp1783 = ~(s1 ? tmp1784 : tmp1785);
  assign tmp1780 = s2 ? tmp1781 : tmp1783;
  assign tmp1776 = ~(s3 ? tmp1777 : tmp1780);
  assign tmp1767 = s4 ? tmp1768 : tmp1776;
  assign tmp1792 = ~(s0 ? tmp1784 : 0);
  assign tmp1791 = s1 ? 1 : tmp1792;
  assign tmp1790 = s2 ? 1 : tmp1791;
  assign tmp1796 = ~(l2 ? tmp110 : tmp33);
  assign tmp1795 = ~(l1 ? tmp24 : tmp1796);
  assign tmp1794 = s1 ? 1 : tmp1795;
  assign tmp1798 = s0 ? tmp1786 : tmp207;
  assign tmp1800 = l1 ? tmp24 : tmp1796;
  assign tmp1799 = s0 ? tmp1800 : tmp1786;
  assign tmp1797 = ~(s1 ? tmp1798 : tmp1799);
  assign tmp1793 = s2 ? tmp1794 : tmp1797;
  assign tmp1789 = s3 ? tmp1790 : tmp1793;
  assign tmp1805 = l1 ? tmp31 : tmp19;
  assign tmp1806 = l1 ? tmp24 : tmp32;
  assign tmp1804 = s0 ? tmp1805 : tmp1806;
  assign tmp1803 = s1 ? tmp1804 : 0;
  assign tmp1802 = s2 ? tmp1803 : 0;
  assign tmp1810 = ~(l1 ? tmp24 : tmp32);
  assign tmp1809 = s0 ? 1 : tmp1810;
  assign tmp1811 = ~(l1 ? tmp24 : tmp19);
  assign tmp1808 = s1 ? tmp1809 : tmp1811;
  assign tmp1812 = ~(s1 ? 1 : tmp1805);
  assign tmp1807 = ~(s2 ? tmp1808 : tmp1812);
  assign tmp1801 = ~(s3 ? tmp1802 : tmp1807);
  assign tmp1788 = s4 ? tmp1789 : tmp1801;
  assign tmp1817 = s0 ? tmp1800 : tmp207;
  assign tmp1816 = s1 ? tmp1817 : 0;
  assign tmp1815 = s2 ? tmp1816 : 0;
  assign tmp1819 = s1 ? tmp19 : tmp54;
  assign tmp1820 = s1 ? tmp1805 : 0;
  assign tmp1818 = s2 ? tmp1819 : tmp1820;
  assign tmp1814 = s3 ? tmp1815 : tmp1818;
  assign tmp1823 = s1 ? 1 : tmp1811;
  assign tmp1822 = s2 ? tmp1823 : 1;
  assign tmp1824 = s1 ? tmp741 : tmp1810;
  assign tmp1821 = ~(s3 ? tmp1822 : tmp1824);
  assign tmp1813 = ~(s4 ? tmp1814 : tmp1821);
  assign tmp1787 = ~(s5 ? tmp1788 : tmp1813);
  assign tmp1766 = s6 ? tmp1767 : tmp1787;
  assign tmp1765 = s7 ? 1 : tmp1766;
  assign tmp1829 = s1 ? tmp1784 : 0;
  assign tmp1828 = s3 ? tmp1829 : tmp1772;
  assign tmp1833 = s0 ? tmp1784 : 0;
  assign tmp1832 = ~(s1 ? tmp1833 : 0);
  assign tmp1831 = s2 ? tmp1775 : tmp1832;
  assign tmp1830 = ~(s3 ? tmp1831 : tmp1780);
  assign tmp1827 = s4 ? tmp1828 : tmp1830;
  assign tmp1839 = s0 ? 1 : tmp1811;
  assign tmp1838 = s1 ? tmp1839 : tmp1811;
  assign tmp1837 = ~(s2 ? tmp1838 : tmp1812);
  assign tmp1836 = ~(s3 ? tmp1802 : tmp1837);
  assign tmp1835 = s4 ? tmp1789 : tmp1836;
  assign tmp1834 = ~(s5 ? tmp1835 : tmp1813);
  assign tmp1826 = s6 ? tmp1827 : tmp1834;
  assign tmp1825 = s7 ? 1 : tmp1826;
  assign tmp1764 = s8 ? tmp1765 : tmp1825;
  assign tmp1846 = s1 ? tmp741 : tmp1811;
  assign tmp1845 = ~(s3 ? tmp1822 : tmp1846);
  assign tmp1844 = ~(s4 ? tmp1814 : tmp1845);
  assign tmp1843 = ~(s5 ? tmp1788 : tmp1844);
  assign tmp1842 = s6 ? tmp1767 : tmp1843;
  assign tmp1841 = s7 ? 1 : tmp1842;
  assign tmp1840 = s8 ? tmp1825 : tmp1841;
  assign tmp1763 = s9 ? tmp1764 : tmp1840;
  assign tmp1848 = s8 ? tmp1825 : 1;
  assign tmp1850 = s7 ? tmp1766 : tmp1842;
  assign tmp1849 = s8 ? tmp1850 : tmp1826;
  assign tmp1847 = s9 ? tmp1848 : tmp1849;
  assign tmp1762 = s10 ? tmp1763 : tmp1847;
  assign tmp1672 = s12 ? tmp1673 : tmp1762;
  assign tmp1860 = l1 ? tmp927 : tmp164;
  assign tmp1862 = l1 ? tmp1684 : tmp81;
  assign tmp1861 = ~(s0 ? tmp135 : tmp1862);
  assign tmp1859 = s1 ? tmp1860 : tmp1861;
  assign tmp1865 = l1 ? tmp966 : tmp316;
  assign tmp1866 = ~(l1 ? tmp1689 : tmp164);
  assign tmp1864 = s0 ? tmp1865 : tmp1866;
  assign tmp1868 = s0 ? tmp1865 : 1;
  assign tmp1867 = s1 ? tmp1868 : tmp1866;
  assign tmp1863 = ~(s2 ? tmp1864 : tmp1867);
  assign tmp1858 = s3 ? tmp1859 : tmp1863;
  assign tmp1872 = s0 ? tmp1401 : 1;
  assign tmp1871 = s1 ? tmp1872 : tmp1866;
  assign tmp1874 = s0 ? tmp1860 : 0;
  assign tmp1873 = ~(s1 ? tmp1874 : tmp55);
  assign tmp1870 = s2 ? tmp1871 : tmp1873;
  assign tmp1877 = ~(l1 ? tmp74 : tmp185);
  assign tmp1876 = s1 ? tmp135 : tmp1877;
  assign tmp1880 = l1 ? tmp1689 : tmp164;
  assign tmp1881 = l1 ? tmp19 : tmp164;
  assign tmp1879 = s0 ? tmp1880 : tmp1881;
  assign tmp1882 = s0 ? tmp1121 : tmp1880;
  assign tmp1878 = ~(s1 ? tmp1879 : tmp1882);
  assign tmp1875 = s2 ? tmp1876 : tmp1878;
  assign tmp1869 = ~(s3 ? tmp1870 : tmp1875);
  assign tmp1857 = s4 ? tmp1858 : tmp1869;
  assign tmp1888 = s0 ? tmp1862 : 1;
  assign tmp1887 = s1 ? tmp1888 : 1;
  assign tmp1890 = ~(s0 ? tmp1881 : 0);
  assign tmp1889 = s1 ? tmp1862 : tmp1890;
  assign tmp1886 = s2 ? tmp1887 : tmp1889;
  assign tmp1893 = l1 ? tmp322 : tmp316;
  assign tmp1894 = ~(l1 ? tmp19 : tmp18);
  assign tmp1892 = s1 ? tmp1893 : tmp1894;
  assign tmp1896 = s0 ? tmp1121 : tmp603;
  assign tmp1898 = l1 ? tmp1689 : tmp18;
  assign tmp1897 = s0 ? tmp1898 : tmp1119;
  assign tmp1895 = ~(s1 ? tmp1896 : tmp1897);
  assign tmp1891 = s2 ? tmp1892 : tmp1895;
  assign tmp1885 = s3 ? tmp1886 : tmp1891;
  assign tmp1902 = s0 ? tmp221 : tmp1898;
  assign tmp1901 = s1 ? tmp1902 : tmp82;
  assign tmp1903 = ~(l1 ? 1 : tmp81);
  assign tmp1900 = s2 ? tmp1901 : tmp1903;
  assign tmp1907 = ~(l1 ? tmp19 : tmp901);
  assign tmp1906 = s0 ? tmp1401 : tmp1907;
  assign tmp1905 = s1 ? tmp1906 : tmp1894;
  assign tmp1908 = ~(s1 ? tmp375 : tmp224);
  assign tmp1904 = ~(s2 ? tmp1905 : tmp1908);
  assign tmp1899 = ~(s3 ? tmp1900 : tmp1904);
  assign tmp1884 = s4 ? tmp1885 : tmp1899;
  assign tmp1913 = s0 ? tmp1119 : tmp83;
  assign tmp1912 = s1 ? tmp1913 : tmp94;
  assign tmp1911 = s2 ? tmp1912 : 0;
  assign tmp1915 = s1 ? tmp83 : tmp566;
  assign tmp1917 = ~(l1 ? 1 : tmp102);
  assign tmp1916 = ~(s1 ? 1 : tmp1917);
  assign tmp1914 = ~(s2 ? tmp1915 : tmp1916);
  assign tmp1910 = s3 ? tmp1911 : tmp1914;
  assign tmp1920 = s1 ? tmp363 : tmp1121;
  assign tmp1921 = ~(l1 ? tmp322 : tmp81);
  assign tmp1919 = s2 ? tmp1920 : tmp1921;
  assign tmp1922 = s1 ? tmp552 : tmp1427;
  assign tmp1918 = s3 ? tmp1919 : tmp1922;
  assign tmp1909 = ~(s4 ? tmp1910 : tmp1918);
  assign tmp1883 = ~(s5 ? tmp1884 : tmp1909);
  assign tmp1856 = s6 ? tmp1857 : tmp1883;
  assign tmp1855 = s7 ? 1 : tmp1856;
  assign tmp1929 = l1 ? 1 : tmp116;
  assign tmp1930 = l1 ? tmp1684 : tmp17;
  assign tmp1928 = ~(s0 ? tmp1929 : tmp1930);
  assign tmp1927 = s1 ? tmp1169 : tmp1928;
  assign tmp1933 = l1 ? tmp966 : tmp17;
  assign tmp1934 = ~(l1 ? tmp1689 : tmp840);
  assign tmp1932 = s0 ? tmp1933 : tmp1934;
  assign tmp1936 = s0 ? tmp1933 : 1;
  assign tmp1938 = l1 ? tmp1689 : tmp840;
  assign tmp1939 = l1 ? tmp1689 : tmp21;
  assign tmp1937 = ~(s0 ? tmp1938 : tmp1939);
  assign tmp1935 = s1 ? tmp1936 : tmp1937;
  assign tmp1931 = ~(s2 ? tmp1932 : tmp1935);
  assign tmp1926 = s3 ? tmp1927 : tmp1931;
  assign tmp1944 = l1 ? 1 : tmp17;
  assign tmp1943 = s0 ? tmp1944 : 1;
  assign tmp1945 = ~(s0 ? tmp1939 : tmp1938);
  assign tmp1942 = s1 ? tmp1943 : tmp1945;
  assign tmp1947 = s0 ? tmp1169 : 0;
  assign tmp1946 = ~(s1 ? tmp1947 : tmp1039);
  assign tmp1941 = s2 ? tmp1942 : tmp1946;
  assign tmp1949 = s1 ? tmp1929 : tmp1877;
  assign tmp1952 = l1 ? tmp19 : tmp840;
  assign tmp1951 = s0 ? tmp1938 : tmp1952;
  assign tmp1954 = l1 ? tmp19 : tmp811;
  assign tmp1953 = s0 ? tmp1954 : tmp1938;
  assign tmp1950 = ~(s1 ? tmp1951 : tmp1953);
  assign tmp1948 = s2 ? tmp1949 : tmp1950;
  assign tmp1940 = ~(s3 ? tmp1941 : tmp1948);
  assign tmp1925 = s4 ? tmp1926 : tmp1940;
  assign tmp1960 = s0 ? tmp1930 : 1;
  assign tmp1959 = s1 ? tmp1960 : 1;
  assign tmp1962 = ~(s0 ? tmp1952 : 0);
  assign tmp1961 = s1 ? tmp1930 : tmp1962;
  assign tmp1958 = s2 ? tmp1959 : tmp1961;
  assign tmp1965 = l1 ? tmp322 : tmp17;
  assign tmp1966 = ~(l1 ? tmp19 : tmp1203);
  assign tmp1964 = s1 ? tmp1965 : tmp1966;
  assign tmp1968 = s0 ? tmp1954 : tmp603;
  assign tmp1970 = l1 ? tmp1689 : tmp1203;
  assign tmp1971 = l1 ? tmp19 : tmp1203;
  assign tmp1969 = s0 ? tmp1970 : tmp1971;
  assign tmp1967 = ~(s1 ? tmp1968 : tmp1969);
  assign tmp1963 = s2 ? tmp1964 : tmp1967;
  assign tmp1957 = s3 ? tmp1958 : tmp1963;
  assign tmp1976 = l1 ? tmp1689 : tmp1128;
  assign tmp1975 = s0 ? tmp221 : tmp1976;
  assign tmp1977 = ~(s0 ? 1 : tmp1944);
  assign tmp1974 = s1 ? tmp1975 : tmp1977;
  assign tmp1973 = s2 ? tmp1974 : tmp1039;
  assign tmp1981 = ~(l1 ? tmp19 : tmp898);
  assign tmp1980 = s0 ? tmp1944 : tmp1981;
  assign tmp1979 = s1 ? tmp1980 : tmp1894;
  assign tmp1978 = ~(s2 ? tmp1979 : tmp1908);
  assign tmp1972 = ~(s3 ? tmp1973 : tmp1978);
  assign tmp1956 = s4 ? tmp1957 : tmp1972;
  assign tmp1986 = s0 ? tmp1971 : tmp83;
  assign tmp1985 = s1 ? tmp1986 : tmp1265;
  assign tmp1984 = s2 ? tmp1985 : 0;
  assign tmp1983 = s3 ? tmp1984 : tmp1914;
  assign tmp1989 = s1 ? tmp363 : tmp1954;
  assign tmp1990 = ~(l1 ? tmp322 : tmp17);
  assign tmp1988 = s2 ? tmp1989 : tmp1990;
  assign tmp1987 = s3 ? tmp1988 : tmp1922;
  assign tmp1982 = ~(s4 ? tmp1983 : tmp1987);
  assign tmp1955 = ~(s5 ? tmp1956 : tmp1982);
  assign tmp1924 = s6 ? tmp1925 : tmp1955;
  assign tmp1923 = s7 ? 1 : tmp1924;
  assign tmp1854 = s8 ? tmp1855 : tmp1923;
  assign tmp1997 = l1 ? tmp927 : tmp324;
  assign tmp1999 = l1 ? tmp1684 : tmp392;
  assign tmp1998 = ~(s0 ? tmp1929 : tmp1999);
  assign tmp1996 = s1 ? tmp1997 : tmp1998;
  assign tmp2002 = l1 ? tmp966 : tmp116;
  assign tmp2003 = ~(l1 ? tmp1689 : tmp779);
  assign tmp2001 = s0 ? tmp2002 : tmp2003;
  assign tmp2005 = s0 ? tmp2002 : 1;
  assign tmp2007 = l1 ? tmp1689 : tmp779;
  assign tmp2008 = l1 ? tmp1689 : tmp324;
  assign tmp2006 = ~(s0 ? tmp2007 : tmp2008);
  assign tmp2004 = s1 ? tmp2005 : tmp2006;
  assign tmp2000 = ~(s2 ? tmp2001 : tmp2004);
  assign tmp1995 = s3 ? tmp1996 : tmp2000;
  assign tmp2013 = l1 ? 1 : tmp392;
  assign tmp2012 = s0 ? tmp2013 : 1;
  assign tmp2014 = ~(s0 ? tmp2008 : tmp2007);
  assign tmp2011 = s1 ? tmp2012 : tmp2014;
  assign tmp2016 = s0 ? tmp1997 : 0;
  assign tmp2015 = ~(s1 ? tmp2016 : tmp1039);
  assign tmp2010 = s2 ? tmp2011 : tmp2015;
  assign tmp2020 = l1 ? tmp19 : tmp779;
  assign tmp2019 = s0 ? tmp2007 : tmp2020;
  assign tmp2021 = s0 ? tmp1954 : tmp2007;
  assign tmp2018 = ~(s1 ? tmp2019 : tmp2021);
  assign tmp2017 = s2 ? tmp1949 : tmp2018;
  assign tmp2009 = ~(s3 ? tmp2010 : tmp2017);
  assign tmp1994 = s4 ? tmp1995 : tmp2009;
  assign tmp2027 = s0 ? tmp1999 : 1;
  assign tmp2026 = s1 ? tmp2027 : 1;
  assign tmp2029 = l1 ? tmp1684 : tmp373;
  assign tmp2030 = ~(s0 ? tmp2020 : 0);
  assign tmp2028 = s1 ? tmp2029 : tmp2030;
  assign tmp2025 = s2 ? tmp2026 : tmp2028;
  assign tmp2033 = l1 ? tmp322 : tmp116;
  assign tmp2034 = ~(l1 ? tmp19 : tmp811);
  assign tmp2032 = s1 ? tmp2033 : tmp2034;
  assign tmp2037 = l1 ? tmp1689 : tmp811;
  assign tmp2036 = s0 ? tmp2037 : tmp1954;
  assign tmp2035 = ~(s1 ? tmp1968 : tmp2036);
  assign tmp2031 = s2 ? tmp2032 : tmp2035;
  assign tmp2024 = s3 ? tmp2025 : tmp2031;
  assign tmp2042 = l1 ? tmp1689 : tmp356;
  assign tmp2041 = s0 ? tmp221 : tmp2042;
  assign tmp2040 = s1 ? tmp2041 : tmp1977;
  assign tmp2043 = ~(l1 ? 1 : tmp373);
  assign tmp2039 = s2 ? tmp2040 : tmp2043;
  assign tmp2047 = l1 ? 1 : tmp373;
  assign tmp2048 = ~(l1 ? tmp19 : tmp356);
  assign tmp2046 = s0 ? tmp2047 : tmp2048;
  assign tmp2049 = ~(l1 ? tmp19 : tmp185);
  assign tmp2045 = s1 ? tmp2046 : tmp2049;
  assign tmp2044 = ~(s2 ? tmp2045 : tmp1908);
  assign tmp2038 = ~(s3 ? tmp2039 : tmp2044);
  assign tmp2023 = s4 ? tmp2024 : tmp2038;
  assign tmp2054 = s0 ? tmp1954 : tmp83;
  assign tmp2053 = s1 ? tmp2054 : tmp1265;
  assign tmp2052 = s2 ? tmp2053 : 0;
  assign tmp2056 = ~(s1 ? 1 : tmp54);
  assign tmp2055 = ~(s2 ? tmp1915 : tmp2056);
  assign tmp2051 = s3 ? tmp2052 : tmp2055;
  assign tmp2059 = ~(l1 ? tmp322 : tmp373);
  assign tmp2058 = s2 ? tmp1989 : tmp2059;
  assign tmp2060 = s1 ? tmp552 : tmp363;
  assign tmp2057 = s3 ? tmp2058 : tmp2060;
  assign tmp2050 = ~(s4 ? tmp2051 : tmp2057);
  assign tmp2022 = ~(s5 ? tmp2023 : tmp2050);
  assign tmp1993 = s6 ? tmp1994 : tmp2022;
  assign tmp1992 = s7 ? 1 : tmp1993;
  assign tmp1991 = s8 ? tmp1923 : tmp1992;
  assign tmp1853 = s9 ? tmp1854 : tmp1991;
  assign tmp2062 = s8 ? tmp1923 : 1;
  assign tmp2064 = s7 ? tmp1856 : tmp1993;
  assign tmp2063 = s8 ? tmp2064 : tmp1924;
  assign tmp2061 = s9 ? tmp2062 : tmp2063;
  assign tmp1852 = s10 ? tmp1853 : tmp2061;
  assign tmp2073 = l1 ? tmp966 : tmp1684;
  assign tmp2074 = s0 ? 1 : tmp1692;
  assign tmp2072 = s1 ? tmp2073 : tmp2074;
  assign tmp2078 = l1 ? tmp966 : tmp110;
  assign tmp2077 = s0 ? 1 : tmp2078;
  assign tmp2079 = s0 ? tmp1692 : tmp2078;
  assign tmp2076 = s1 ? tmp2077 : tmp2079;
  assign tmp2080 = s1 ? tmp1694 : tmp2078;
  assign tmp2075 = s2 ? tmp2076 : tmp2080;
  assign tmp2071 = s3 ? tmp2072 : tmp2075;
  assign tmp2083 = s1 ? 1 : tmp2078;
  assign tmp2085 = s0 ? tmp2073 : 1;
  assign tmp2084 = s1 ? tmp2085 : 1;
  assign tmp2082 = s2 ? tmp2083 : tmp2084;
  assign tmp2087 = s1 ? 1 : tmp208;
  assign tmp2090 = l1 ? tmp1123 : tmp110;
  assign tmp2089 = s0 ? tmp2078 : tmp2090;
  assign tmp2091 = s0 ? tmp208 : tmp2078;
  assign tmp2088 = s1 ? tmp2089 : tmp2091;
  assign tmp2086 = s2 ? tmp2087 : tmp2088;
  assign tmp2081 = s3 ? tmp2082 : tmp2086;
  assign tmp2070 = s4 ? tmp2071 : tmp2081;
  assign tmp2096 = s1 ? tmp1694 : 1;
  assign tmp2098 = s0 ? tmp2090 : 1;
  assign tmp2097 = s1 ? tmp1692 : tmp2098;
  assign tmp2095 = s2 ? tmp2096 : tmp2097;
  assign tmp2102 = l2 ? tmp110 : tmp33;
  assign tmp2101 = l1 ? tmp1123 : tmp2102;
  assign tmp2100 = s1 ? tmp594 : tmp2101;
  assign tmp2104 = s0 ? tmp208 : tmp174;
  assign tmp2106 = l1 ? tmp966 : tmp2102;
  assign tmp2107 = l1 ? tmp1123 : tmp33;
  assign tmp2105 = s0 ? tmp2106 : tmp2107;
  assign tmp2103 = s1 ? tmp2104 : tmp2105;
  assign tmp2099 = s2 ? tmp2100 : tmp2103;
  assign tmp2094 = s3 ? tmp2095 : tmp2099;
  assign tmp2112 = l1 ? tmp966 : tmp322;
  assign tmp2111 = s0 ? tmp208 : tmp2112;
  assign tmp2110 = s1 ? tmp2111 : 1;
  assign tmp2109 = s2 ? tmp2110 : 1;
  assign tmp2115 = s0 ? 1 : tmp322;
  assign tmp2114 = s1 ? tmp2115 : tmp2107;
  assign tmp2116 = s1 ? tmp83 : tmp208;
  assign tmp2113 = s2 ? tmp2114 : tmp2116;
  assign tmp2108 = s3 ? tmp2109 : tmp2113;
  assign tmp2093 = s4 ? tmp2094 : tmp2108;
  assign tmp2121 = s0 ? tmp2101 : tmp174;
  assign tmp2120 = s1 ? tmp2121 : tmp31;
  assign tmp2119 = s2 ? tmp2120 : 1;
  assign tmp2123 = s1 ? tmp135 : 1;
  assign tmp2124 = ~(s1 ? tmp208 : 1);
  assign tmp2122 = ~(s2 ? tmp2123 : tmp2124);
  assign tmp2118 = s3 ? tmp2119 : tmp2122;
  assign tmp2127 = s1 ? tmp207 : tmp208;
  assign tmp2128 = l1 ? tmp1123 : 1;
  assign tmp2126 = s2 ? tmp2127 : tmp2128;
  assign tmp2130 = l1 ? tmp31 : tmp323;
  assign tmp2131 = l1 ? tmp1123 : tmp322;
  assign tmp2129 = s1 ? tmp2130 : tmp2131;
  assign tmp2125 = s3 ? tmp2126 : tmp2129;
  assign tmp2117 = s4 ? tmp2118 : tmp2125;
  assign tmp2092 = s5 ? tmp2093 : tmp2117;
  assign tmp2069 = ~(s6 ? tmp2070 : tmp2092);
  assign tmp2068 = s7 ? 1 : tmp2069;
  assign tmp2136 = s1 ? tmp2078 : tmp2074;
  assign tmp2135 = s3 ? tmp2136 : tmp2075;
  assign tmp2140 = s0 ? tmp2078 : 1;
  assign tmp2139 = s1 ? tmp2140 : 1;
  assign tmp2138 = s2 ? tmp2083 : tmp2139;
  assign tmp2137 = s3 ? tmp2138 : tmp2086;
  assign tmp2134 = s4 ? tmp2135 : tmp2137;
  assign tmp2146 = s0 ? 1 : tmp336;
  assign tmp2145 = s1 ? tmp2146 : tmp2107;
  assign tmp2144 = s2 ? tmp2145 : tmp2116;
  assign tmp2143 = s3 ? tmp2109 : tmp2144;
  assign tmp2142 = s4 ? tmp2094 : tmp2143;
  assign tmp2150 = s1 ? tmp2121 : tmp207;
  assign tmp2149 = s2 ? tmp2150 : 1;
  assign tmp2148 = s3 ? tmp2149 : tmp2122;
  assign tmp2147 = s4 ? tmp2148 : tmp2125;
  assign tmp2141 = s5 ? tmp2142 : tmp2147;
  assign tmp2133 = ~(s6 ? tmp2134 : tmp2141);
  assign tmp2132 = s7 ? 1 : tmp2133;
  assign tmp2067 = s8 ? tmp2068 : tmp2132;
  assign tmp2157 = s1 ? tmp2130 : tmp2107;
  assign tmp2156 = s3 ? tmp2126 : tmp2157;
  assign tmp2155 = s4 ? tmp2148 : tmp2156;
  assign tmp2154 = s5 ? tmp2093 : tmp2155;
  assign tmp2153 = ~(s6 ? tmp2070 : tmp2154);
  assign tmp2152 = s7 ? 1 : tmp2153;
  assign tmp2151 = s8 ? tmp2132 : tmp2152;
  assign tmp2066 = s9 ? tmp2067 : tmp2151;
  assign tmp2159 = s8 ? tmp2132 : 1;
  assign tmp2162 = s6 ? tmp2070 : tmp2092;
  assign tmp2163 = s6 ? tmp2070 : tmp2154;
  assign tmp2161 = s7 ? tmp2162 : tmp2163;
  assign tmp2164 = s6 ? tmp2134 : tmp2141;
  assign tmp2160 = ~(s8 ? tmp2161 : tmp2164);
  assign tmp2158 = s9 ? tmp2159 : tmp2160;
  assign tmp2065 = s10 ? tmp2066 : tmp2158;
  assign tmp1851 = s12 ? tmp1852 : tmp2065;
  assign tmp1671 = s13 ? tmp1672 : tmp1851;
  assign tmp2176 = ~(l1 ? tmp1123 : tmp33);
  assign tmp2175 = s0 ? tmp19 : tmp2176;
  assign tmp2174 = s1 ? tmp19 : tmp2175;
  assign tmp2179 = ~(l1 ? tmp897 : tmp19);
  assign tmp2178 = s0 ? tmp336 : tmp2179;
  assign tmp2181 = s0 ? tmp336 : 0;
  assign tmp2180 = s1 ? tmp2181 : tmp2179;
  assign tmp2177 = ~(s2 ? tmp2178 : tmp2180);
  assign tmp2173 = s3 ? tmp2174 : tmp2177;
  assign tmp2184 = s1 ? tmp336 : tmp2179;
  assign tmp2186 = s0 ? tmp19 : 1;
  assign tmp2185 = ~(s1 ? tmp2186 : tmp19);
  assign tmp2183 = s2 ? tmp2184 : tmp2185;
  assign tmp2188 = s1 ? tmp19 : tmp135;
  assign tmp2191 = l1 ? tmp897 : tmp19;
  assign tmp2192 = l1 ? tmp927 : tmp19;
  assign tmp2190 = s0 ? tmp2191 : tmp2192;
  assign tmp2194 = l1 ? tmp316 : tmp19;
  assign tmp2193 = s0 ? tmp2194 : tmp2191;
  assign tmp2189 = s1 ? tmp2190 : tmp2193;
  assign tmp2187 = ~(s2 ? tmp2188 : tmp2189);
  assign tmp2182 = ~(s3 ? tmp2183 : tmp2187);
  assign tmp2172 = s4 ? tmp2173 : tmp2182;
  assign tmp2200 = s0 ? tmp2107 : 0;
  assign tmp2199 = s1 ? tmp2200 : tmp336;
  assign tmp2202 = l1 ? tmp1123 : tmp185;
  assign tmp2203 = ~(s0 ? tmp2192 : 1);
  assign tmp2201 = s1 ? tmp2202 : tmp2203;
  assign tmp2198 = s2 ? tmp2199 : tmp2201;
  assign tmp2206 = ~(l1 ? tmp927 : tmp19);
  assign tmp2205 = s1 ? tmp336 : tmp2206;
  assign tmp2207 = ~(s1 ? tmp2194 : tmp2190);
  assign tmp2204 = s2 ? tmp2205 : tmp2207;
  assign tmp2197 = s3 ? tmp2198 : tmp2204;
  assign tmp2211 = s0 ? tmp19 : tmp2191;
  assign tmp2210 = s1 ? tmp2211 : tmp941;
  assign tmp2212 = ~(l1 ? tmp322 : tmp185);
  assign tmp2209 = s2 ? tmp2210 : tmp2212;
  assign tmp2216 = ~(l1 ? tmp19 : tmp32);
  assign tmp2215 = s0 ? tmp221 : tmp2216;
  assign tmp2214 = s1 ? tmp2215 : tmp2206;
  assign tmp2217 = ~(s1 ? 1 : tmp135);
  assign tmp2213 = ~(s2 ? tmp2214 : tmp2217);
  assign tmp2208 = ~(s3 ? tmp2209 : tmp2213);
  assign tmp2196 = s4 ? tmp2197 : tmp2208;
  assign tmp2222 = s0 ? tmp2192 : 1;
  assign tmp2221 = s1 ? tmp2222 : tmp1757;
  assign tmp2220 = s2 ? tmp2221 : tmp374;
  assign tmp2225 = l1 ? 1 : tmp32;
  assign tmp2224 = s1 ? tmp2225 : 0;
  assign tmp2223 = s2 ? tmp2123 : tmp2224;
  assign tmp2219 = s3 ? tmp2220 : tmp2223;
  assign tmp2229 = ~(l1 ? tmp316 : tmp19);
  assign tmp2228 = s1 ? tmp207 : tmp2229;
  assign tmp2230 = l1 ? tmp966 : tmp185;
  assign tmp2227 = s2 ? tmp2228 : tmp2230;
  assign tmp2232 = ~(l1 ? tmp927 : tmp32);
  assign tmp2231 = s1 ? tmp208 : tmp2232;
  assign tmp2226 = ~(s3 ? tmp2227 : tmp2231);
  assign tmp2218 = ~(s4 ? tmp2219 : tmp2226);
  assign tmp2195 = ~(s5 ? tmp2196 : tmp2218);
  assign tmp2171 = ~(s6 ? tmp2172 : tmp2195);
  assign tmp2170 = s7 ? 1 : tmp2171;
  assign tmp2238 = l1 ? tmp1202 : tmp19;
  assign tmp2240 = l1 ? tmp973 : tmp19;
  assign tmp2239 = s0 ? tmp406 : tmp2240;
  assign tmp2237 = s1 ? tmp2238 : tmp2239;
  assign tmp2243 = l1 ? tmp981 : tmp19;
  assign tmp2242 = s0 ? tmp391 : tmp2243;
  assign tmp2245 = s0 ? tmp391 : tmp135;
  assign tmp2244 = s1 ? tmp2245 : tmp2243;
  assign tmp2241 = s2 ? tmp2242 : tmp2244;
  assign tmp2236 = s3 ? tmp2237 : tmp2241;
  assign tmp2248 = s1 ? tmp391 : tmp2243;
  assign tmp2250 = s0 ? tmp2238 : 1;
  assign tmp2249 = s1 ? tmp2250 : tmp406;
  assign tmp2247 = s2 ? tmp2248 : tmp2249;
  assign tmp2252 = s1 ? tmp406 : tmp135;
  assign tmp2255 = l1 ? tmp1021 : tmp19;
  assign tmp2254 = s0 ? tmp2243 : tmp2255;
  assign tmp2256 = s0 ? tmp2194 : tmp2243;
  assign tmp2253 = s1 ? tmp2254 : tmp2256;
  assign tmp2251 = s2 ? tmp2252 : tmp2253;
  assign tmp2246 = s3 ? tmp2247 : tmp2251;
  assign tmp2235 = s4 ? tmp2236 : tmp2246;
  assign tmp2262 = s0 ? tmp2240 : 1;
  assign tmp2261 = s1 ? tmp2262 : tmp391;
  assign tmp2264 = l1 ? tmp973 : tmp24;
  assign tmp2265 = s0 ? tmp2255 : tmp135;
  assign tmp2263 = s1 ? tmp2264 : tmp2265;
  assign tmp2260 = s2 ? tmp2261 : tmp2263;
  assign tmp2267 = s1 ? tmp391 : tmp2192;
  assign tmp2268 = s1 ? tmp2194 : tmp2254;
  assign tmp2266 = s2 ? tmp2267 : tmp2268;
  assign tmp2259 = s3 ? tmp2260 : tmp2266;
  assign tmp2272 = s0 ? tmp19 : tmp2243;
  assign tmp2273 = s0 ? tmp237 : tmp174;
  assign tmp2271 = s1 ? tmp2272 : tmp2273;
  assign tmp2274 = l1 ? tmp392 : tmp24;
  assign tmp2270 = s2 ? tmp2271 : tmp2274;
  assign tmp2278 = ~(l1 ? tmp1202 : tmp32);
  assign tmp2277 = s0 ? tmp221 : tmp2278;
  assign tmp2276 = s1 ? tmp2277 : tmp2206;
  assign tmp2275 = ~(s2 ? tmp2276 : tmp2217);
  assign tmp2269 = s3 ? tmp2270 : tmp2275;
  assign tmp2258 = s4 ? tmp2259 : tmp2269;
  assign tmp2281 = s2 ? tmp2221 : tmp1553;
  assign tmp2280 = s3 ? tmp2281 : tmp2223;
  assign tmp2279 = s4 ? tmp2280 : tmp2226;
  assign tmp2257 = s5 ? tmp2258 : tmp2279;
  assign tmp2234 = ~(s6 ? tmp2235 : tmp2257);
  assign tmp2233 = s7 ? 1 : tmp2234;
  assign tmp2169 = s8 ? tmp2170 : tmp2233;
  assign tmp2288 = l1 ? tmp1202 : tmp392;
  assign tmp2290 = l1 ? tmp973 : tmp392;
  assign tmp2289 = s0 ? tmp975 : tmp2290;
  assign tmp2287 = s1 ? tmp2288 : tmp2289;
  assign tmp2294 = l1 ? tmp981 : tmp1202;
  assign tmp2293 = s0 ? tmp1568 : tmp2294;
  assign tmp2296 = l1 ? tmp392 : tmp116;
  assign tmp2295 = s0 ? tmp2296 : tmp2294;
  assign tmp2292 = s1 ? tmp2293 : tmp2295;
  assign tmp2298 = s0 ? tmp2296 : 1;
  assign tmp2300 = l1 ? tmp981 : tmp392;
  assign tmp2299 = s0 ? tmp2294 : tmp2300;
  assign tmp2297 = s1 ? tmp2298 : tmp2299;
  assign tmp2291 = s2 ? tmp2292 : tmp2297;
  assign tmp2286 = s3 ? tmp2287 : tmp2291;
  assign tmp2304 = s0 ? tmp392 : tmp237;
  assign tmp2305 = s0 ? tmp2300 : tmp2294;
  assign tmp2303 = s1 ? tmp2304 : tmp2305;
  assign tmp2307 = s0 ? tmp2288 : 1;
  assign tmp2306 = s1 ? tmp2307 : tmp994;
  assign tmp2302 = s2 ? tmp2303 : tmp2306;
  assign tmp2309 = s1 ? tmp975 : tmp135;
  assign tmp2312 = l1 ? tmp1021 : tmp1202;
  assign tmp2311 = s0 ? tmp2294 : tmp2312;
  assign tmp2314 = l1 ? tmp316 : tmp1202;
  assign tmp2313 = s0 ? tmp2314 : tmp2294;
  assign tmp2310 = s1 ? tmp2311 : tmp2313;
  assign tmp2308 = s2 ? tmp2309 : tmp2310;
  assign tmp2301 = s3 ? tmp2302 : tmp2308;
  assign tmp2285 = s4 ? tmp2286 : tmp2301;
  assign tmp2320 = s0 ? tmp2290 : 1;
  assign tmp2319 = s1 ? tmp2320 : tmp1568;
  assign tmp2322 = l1 ? tmp973 : tmp373;
  assign tmp2323 = s0 ? tmp2312 : 1;
  assign tmp2321 = s1 ? tmp2322 : tmp2323;
  assign tmp2318 = s2 ? tmp2319 : tmp2321;
  assign tmp2326 = l1 ? tmp927 : tmp1202;
  assign tmp2325 = s1 ? tmp2296 : tmp2326;
  assign tmp2328 = s0 ? tmp2314 : 1;
  assign tmp2327 = s1 ? tmp2328 : tmp2311;
  assign tmp2324 = s2 ? tmp2325 : tmp2327;
  assign tmp2317 = s3 ? tmp2318 : tmp2324;
  assign tmp2332 = s0 ? tmp19 : tmp2300;
  assign tmp2331 = s1 ? tmp2332 : tmp1027;
  assign tmp2333 = l1 ? tmp392 : tmp373;
  assign tmp2330 = s2 ? tmp2331 : tmp2333;
  assign tmp2337 = ~(l1 ? tmp1202 : tmp392);
  assign tmp2336 = s0 ? tmp767 : tmp2337;
  assign tmp2335 = s1 ? tmp2336 : tmp2206;
  assign tmp2334 = ~(s2 ? tmp2335 : tmp2217);
  assign tmp2329 = s3 ? tmp2330 : tmp2334;
  assign tmp2316 = s4 ? tmp2317 : tmp2329;
  assign tmp2342 = s0 ? tmp2326 : 1;
  assign tmp2343 = ~(l1 ? tmp31 : tmp21);
  assign tmp2341 = s1 ? tmp2342 : tmp2343;
  assign tmp2340 = s2 ? tmp2341 : tmp1608;
  assign tmp2339 = s3 ? tmp2340 : tmp2223;
  assign tmp2347 = ~(l1 ? tmp316 : tmp1202);
  assign tmp2346 = s1 ? tmp207 : tmp2347;
  assign tmp2348 = l1 ? tmp966 : tmp356;
  assign tmp2345 = s2 ? tmp2346 : tmp2348;
  assign tmp2344 = ~(s3 ? tmp2345 : tmp2231);
  assign tmp2338 = s4 ? tmp2339 : tmp2344;
  assign tmp2315 = s5 ? tmp2316 : tmp2338;
  assign tmp2284 = ~(s6 ? tmp2285 : tmp2315);
  assign tmp2283 = s7 ? 1 : tmp2284;
  assign tmp2282 = s8 ? tmp2233 : tmp2283;
  assign tmp2168 = s9 ? tmp2169 : tmp2282;
  assign tmp2357 = s0 ? tmp1624 : tmp2294;
  assign tmp2358 = s0 ? tmp392 : tmp2294;
  assign tmp2356 = s1 ? tmp2357 : tmp2358;
  assign tmp2360 = s0 ? tmp392 : 1;
  assign tmp2359 = s1 ? tmp2360 : tmp2299;
  assign tmp2355 = s2 ? tmp2356 : tmp2359;
  assign tmp2354 = s3 ? tmp2287 : tmp2355;
  assign tmp2353 = s4 ? tmp2354 : tmp2301;
  assign tmp2365 = s1 ? tmp2320 : tmp1624;
  assign tmp2364 = s2 ? tmp2365 : tmp2321;
  assign tmp2367 = s1 ? tmp392 : tmp2326;
  assign tmp2366 = s2 ? tmp2367 : tmp2327;
  assign tmp2363 = s3 ? tmp2364 : tmp2366;
  assign tmp2362 = s4 ? tmp2363 : tmp2329;
  assign tmp2370 = s2 ? tmp2341 : tmp374;
  assign tmp2369 = s3 ? tmp2370 : tmp2223;
  assign tmp2368 = s4 ? tmp2369 : tmp2344;
  assign tmp2361 = s5 ? tmp2362 : tmp2368;
  assign tmp2352 = ~(s6 ? tmp2353 : tmp2361);
  assign tmp2351 = s7 ? 1 : tmp2352;
  assign tmp2350 = s8 ? tmp2351 : 1;
  assign tmp2373 = s6 ? tmp2172 : tmp2195;
  assign tmp2374 = s6 ? tmp2285 : tmp2315;
  assign tmp2372 = s7 ? tmp2373 : tmp2374;
  assign tmp2376 = s6 ? tmp2235 : tmp2257;
  assign tmp2377 = s6 ? tmp2353 : tmp2361;
  assign tmp2375 = s7 ? tmp2376 : tmp2377;
  assign tmp2371 = ~(s8 ? tmp2372 : tmp2375);
  assign tmp2349 = s9 ? tmp2350 : tmp2371;
  assign tmp2167 = s10 ? tmp2168 : tmp2349;
  assign tmp2386 = l1 ? tmp81 : tmp897;
  assign tmp2388 = ~(l1 ? tmp15 : tmp917);
  assign tmp2387 = s0 ? tmp135 : tmp2388;
  assign tmp2385 = s1 ? tmp2386 : tmp2387;
  assign tmp2391 = l1 ? tmp26 : tmp33;
  assign tmp2393 = l2 ? tmp19 : tmp110;
  assign tmp2392 = ~(l1 ? tmp2393 : tmp897);
  assign tmp2390 = s0 ? tmp2391 : tmp2392;
  assign tmp2395 = s0 ? tmp2391 : 0;
  assign tmp2394 = s1 ? tmp2395 : tmp2392;
  assign tmp2389 = ~(s2 ? tmp2390 : tmp2394);
  assign tmp2384 = s3 ? tmp2385 : tmp2389;
  assign tmp2400 = l1 ? tmp31 : tmp917;
  assign tmp2399 = s0 ? tmp2400 : 0;
  assign tmp2398 = s1 ? tmp2399 : tmp2392;
  assign tmp2402 = s0 ? tmp2386 : 1;
  assign tmp2401 = ~(s1 ? tmp2402 : tmp135);
  assign tmp2397 = s2 ? tmp2398 : tmp2401;
  assign tmp2404 = s1 ? tmp135 : tmp1893;
  assign tmp2407 = l1 ? tmp2393 : tmp897;
  assign tmp2408 = l1 ? tmp117 : tmp897;
  assign tmp2406 = s0 ? tmp2407 : tmp2408;
  assign tmp2410 = l1 ? tmp117 : tmp316;
  assign tmp2409 = s0 ? tmp2410 : tmp2407;
  assign tmp2405 = s1 ? tmp2406 : tmp2409;
  assign tmp2403 = ~(s2 ? tmp2404 : tmp2405);
  assign tmp2396 = ~(s3 ? tmp2397 : tmp2403);
  assign tmp2383 = s4 ? tmp2384 : tmp2396;
  assign tmp2417 = l1 ? tmp15 : tmp917;
  assign tmp2416 = s0 ? tmp2417 : 0;
  assign tmp2415 = s1 ? tmp2416 : tmp208;
  assign tmp2419 = l1 ? tmp15 : tmp933;
  assign tmp2420 = ~(s0 ? tmp2408 : 1);
  assign tmp2418 = s1 ? tmp2419 : tmp2420;
  assign tmp2414 = s2 ? tmp2415 : tmp2418;
  assign tmp2423 = ~(l1 ? tmp117 : tmp927);
  assign tmp2422 = s1 ? tmp1298 : tmp2423;
  assign tmp2425 = s0 ? tmp2410 : tmp594;
  assign tmp2427 = l1 ? tmp2393 : tmp927;
  assign tmp2428 = l1 ? tmp117 : tmp927;
  assign tmp2426 = s0 ? tmp2427 : tmp2428;
  assign tmp2424 = ~(s1 ? tmp2425 : tmp2426);
  assign tmp2421 = s2 ? tmp2422 : tmp2424;
  assign tmp2413 = s3 ? tmp2414 : tmp2421;
  assign tmp2433 = l1 ? tmp31 : tmp316;
  assign tmp2432 = s0 ? tmp2433 : tmp2427;
  assign tmp2434 = s0 ? 1 : tmp83;
  assign tmp2431 = s1 ? tmp2432 : tmp2434;
  assign tmp2435 = ~(l1 ? tmp31 : tmp933);
  assign tmp2430 = s2 ? tmp2431 : tmp2435;
  assign tmp2439 = l1 ? tmp31 : tmp933;
  assign tmp2440 = ~(l1 ? tmp117 : tmp948);
  assign tmp2438 = s0 ? tmp2439 : tmp2440;
  assign tmp2437 = s1 ? tmp2438 : tmp2423;
  assign tmp2441 = ~(s1 ? 1 : tmp1893);
  assign tmp2436 = ~(s2 ? tmp2437 : tmp2441);
  assign tmp2429 = ~(s3 ? tmp2430 : tmp2436);
  assign tmp2412 = s4 ? tmp2413 : tmp2429;
  assign tmp2446 = s0 ? tmp2428 : tmp31;
  assign tmp2445 = s1 ? tmp2446 : 0;
  assign tmp2447 = ~(s1 ? tmp202 : tmp207);
  assign tmp2444 = s2 ? tmp2445 : tmp2447;
  assign tmp2449 = s1 ? 1 : tmp569;
  assign tmp2451 = ~(l1 ? tmp31 : tmp966);
  assign tmp2450 = s1 ? tmp202 : tmp2451;
  assign tmp2448 = s2 ? tmp2449 : tmp2450;
  assign tmp2443 = s3 ? tmp2444 : tmp2448;
  assign tmp2455 = ~(l1 ? tmp117 : tmp316);
  assign tmp2454 = s1 ? tmp74 : tmp2455;
  assign tmp2456 = l1 ? tmp74 : tmp933;
  assign tmp2453 = s2 ? tmp2454 : tmp2456;
  assign tmp2457 = s1 ? tmp618 : tmp2440;
  assign tmp2452 = ~(s3 ? tmp2453 : tmp2457);
  assign tmp2442 = ~(s4 ? tmp2443 : tmp2452);
  assign tmp2411 = ~(s5 ? tmp2412 : tmp2442);
  assign tmp2382 = ~(s6 ? tmp2383 : tmp2411);
  assign tmp2381 = s7 ? 1 : tmp2382;
  assign tmp2464 = l2 ? tmp780 : tmp17;
  assign tmp2463 = l1 ? tmp2464 : tmp897;
  assign tmp2466 = l1 ? tmp109 : tmp897;
  assign tmp2465 = s0 ? tmp135 : tmp2466;
  assign tmp2462 = s1 ? tmp2463 : tmp2465;
  assign tmp2469 = l1 ? tmp17 : tmp19;
  assign tmp2471 = l2 ? tmp780 : tmp110;
  assign tmp2470 = l1 ? tmp2471 : tmp897;
  assign tmp2468 = s0 ? tmp2469 : tmp2470;
  assign tmp2473 = s0 ? tmp2469 : tmp135;
  assign tmp2472 = s1 ? tmp2473 : tmp2470;
  assign tmp2467 = s2 ? tmp2468 : tmp2472;
  assign tmp2461 = s3 ? tmp2462 : tmp2467;
  assign tmp2478 = l1 ? tmp116 : tmp897;
  assign tmp2477 = s0 ? tmp2478 : 1;
  assign tmp2476 = s1 ? tmp2477 : tmp2470;
  assign tmp2480 = s0 ? tmp2463 : 1;
  assign tmp2479 = s1 ? tmp2480 : tmp135;
  assign tmp2475 = s2 ? tmp2476 : tmp2479;
  assign tmp2485 = l2 ? tmp780 : tmp33;
  assign tmp2484 = l1 ? tmp2485 : tmp897;
  assign tmp2483 = s0 ? tmp2470 : tmp2484;
  assign tmp2486 = s0 ? tmp2410 : tmp2470;
  assign tmp2482 = s1 ? tmp2483 : tmp2486;
  assign tmp2481 = s2 ? tmp2404 : tmp2482;
  assign tmp2474 = s3 ? tmp2475 : tmp2481;
  assign tmp2460 = s4 ? tmp2461 : tmp2474;
  assign tmp2492 = s0 ? tmp2466 : 1;
  assign tmp2493 = l1 ? tmp116 : tmp19;
  assign tmp2491 = s1 ? tmp2492 : tmp2493;
  assign tmp2495 = l1 ? tmp109 : tmp927;
  assign tmp2496 = s0 ? tmp2484 : tmp135;
  assign tmp2494 = s1 ? tmp2495 : tmp2496;
  assign tmp2490 = s2 ? tmp2491 : tmp2494;
  assign tmp2499 = l1 ? tmp898 : tmp33;
  assign tmp2498 = s1 ? tmp2499 : tmp2423;
  assign tmp2502 = l1 ? tmp2471 : tmp927;
  assign tmp2503 = l1 ? tmp2485 : tmp927;
  assign tmp2501 = s0 ? tmp2502 : tmp2503;
  assign tmp2500 = ~(s1 ? tmp2425 : tmp2501);
  assign tmp2497 = ~(s2 ? tmp2498 : tmp2500);
  assign tmp2489 = s3 ? tmp2490 : tmp2497;
  assign tmp2507 = s0 ? tmp2433 : tmp2502;
  assign tmp2506 = s1 ? tmp2507 : tmp2434;
  assign tmp2508 = l1 ? tmp116 : tmp927;
  assign tmp2505 = s2 ? tmp2506 : tmp2508;
  assign tmp2512 = ~(l1 ? tmp2485 : tmp948);
  assign tmp2511 = s0 ? tmp2439 : tmp2512;
  assign tmp2510 = s1 ? tmp2511 : tmp2423;
  assign tmp2509 = ~(s2 ? tmp2510 : tmp2441);
  assign tmp2504 = s3 ? tmp2505 : tmp2509;
  assign tmp2488 = s4 ? tmp2489 : tmp2504;
  assign tmp2516 = ~(s1 ? tmp187 : tmp207);
  assign tmp2515 = s2 ? tmp2445 : tmp2516;
  assign tmp2514 = s3 ? tmp2515 : tmp2448;
  assign tmp2513 = s4 ? tmp2514 : tmp2452;
  assign tmp2487 = s5 ? tmp2488 : tmp2513;
  assign tmp2459 = ~(s6 ? tmp2460 : tmp2487);
  assign tmp2458 = s7 ? 1 : tmp2459;
  assign tmp2380 = s8 ? tmp2381 : tmp2458;
  assign tmp2523 = l1 ? tmp2464 : tmp116;
  assign tmp2525 = l1 ? tmp109 : tmp116;
  assign tmp2524 = s0 ? tmp1929 : tmp2525;
  assign tmp2522 = s1 ? tmp2523 : tmp2524;
  assign tmp2528 = l1 ? tmp17 : tmp116;
  assign tmp2529 = l1 ? tmp2471 : tmp1002;
  assign tmp2527 = s0 ? tmp2528 : tmp2529;
  assign tmp2531 = s0 ? tmp2528 : 1;
  assign tmp2533 = l1 ? tmp2471 : tmp116;
  assign tmp2532 = s0 ? tmp2529 : tmp2533;
  assign tmp2530 = s1 ? tmp2531 : tmp2532;
  assign tmp2526 = s2 ? tmp2527 : tmp2530;
  assign tmp2521 = s3 ? tmp2522 : tmp2526;
  assign tmp2537 = s0 ? tmp116 : 1;
  assign tmp2538 = s0 ? tmp2533 : tmp2529;
  assign tmp2536 = s1 ? tmp2537 : tmp2538;
  assign tmp2540 = s0 ? tmp2523 : 1;
  assign tmp2539 = s1 ? tmp2540 : tmp1944;
  assign tmp2535 = s2 ? tmp2536 : tmp2539;
  assign tmp2542 = s1 ? tmp1929 : tmp1893;
  assign tmp2545 = l1 ? tmp2485 : tmp1002;
  assign tmp2544 = s0 ? tmp2529 : tmp2545;
  assign tmp2547 = l1 ? tmp117 : tmp1002;
  assign tmp2546 = s0 ? tmp2547 : tmp2529;
  assign tmp2543 = s1 ? tmp2544 : tmp2546;
  assign tmp2541 = s2 ? tmp2542 : tmp2543;
  assign tmp2534 = s3 ? tmp2535 : tmp2541;
  assign tmp2520 = s4 ? tmp2521 : tmp2534;
  assign tmp2553 = s0 ? tmp2525 : 1;
  assign tmp2554 = l1 ? tmp116 : 1;
  assign tmp2552 = s1 ? tmp2553 : tmp2554;
  assign tmp2556 = s0 ? tmp2545 : 1;
  assign tmp2555 = s1 ? tmp2525 : tmp2556;
  assign tmp2551 = s2 ? tmp2552 : tmp2555;
  assign tmp2560 = ~(l2 ? tmp17 : 1);
  assign tmp2559 = l1 ? tmp898 : tmp2560;
  assign tmp2561 = ~(l1 ? tmp117 : tmp1002);
  assign tmp2558 = s1 ? tmp2559 : tmp2561;
  assign tmp2563 = s0 ? tmp2547 : tmp594;
  assign tmp2562 = ~(s1 ? tmp2563 : tmp2544);
  assign tmp2557 = ~(s2 ? tmp2558 : tmp2562);
  assign tmp2550 = s3 ? tmp2551 : tmp2557;
  assign tmp2567 = s0 ? tmp2433 : tmp2533;
  assign tmp2568 = s0 ? 1 : tmp1944;
  assign tmp2566 = s1 ? tmp2567 : tmp2568;
  assign tmp2565 = s2 ? tmp2566 : tmp116;
  assign tmp2572 = l1 ? tmp31 : tmp2560;
  assign tmp2573 = ~(l1 ? tmp2485 : tmp116);
  assign tmp2571 = s0 ? tmp2572 : tmp2573;
  assign tmp2570 = s1 ? tmp2571 : tmp2455;
  assign tmp2569 = ~(s2 ? tmp2570 : tmp2441);
  assign tmp2564 = s3 ? tmp2565 : tmp2569;
  assign tmp2549 = s4 ? tmp2550 : tmp2564;
  assign tmp2578 = s0 ? tmp2547 : tmp31;
  assign tmp2577 = s1 ? tmp2578 : tmp830;
  assign tmp2579 = ~(s1 ? tmp174 : tmp31);
  assign tmp2576 = s2 ? tmp2577 : tmp2579;
  assign tmp2581 = s1 ? tmp202 : tmp203;
  assign tmp2580 = s2 ? tmp2449 : tmp2581;
  assign tmp2575 = s3 ? tmp2576 : tmp2580;
  assign tmp2584 = s1 ? tmp74 : tmp2561;
  assign tmp2585 = l1 ? tmp74 : tmp2560;
  assign tmp2583 = s2 ? tmp2584 : tmp2585;
  assign tmp2587 = ~(l1 ? tmp117 : tmp203);
  assign tmp2586 = s1 ? tmp618 : tmp2587;
  assign tmp2582 = ~(s3 ? tmp2583 : tmp2586);
  assign tmp2574 = s4 ? tmp2575 : tmp2582;
  assign tmp2548 = s5 ? tmp2549 : tmp2574;
  assign tmp2519 = ~(s6 ? tmp2520 : tmp2548);
  assign tmp2518 = s7 ? 1 : tmp2519;
  assign tmp2517 = s8 ? tmp2458 : tmp2518;
  assign tmp2379 = s9 ? tmp2380 : tmp2517;
  assign tmp2595 = l1 ? tmp2464 : tmp973;
  assign tmp2597 = l1 ? tmp109 : tmp973;
  assign tmp2596 = s0 ? tmp1929 : tmp2597;
  assign tmp2594 = s1 ? tmp2595 : tmp2596;
  assign tmp2600 = l1 ? tmp17 : tmp392;
  assign tmp2601 = l1 ? tmp2471 : tmp981;
  assign tmp2599 = s0 ? tmp2600 : tmp2601;
  assign tmp2603 = s0 ? tmp2600 : 1;
  assign tmp2605 = l1 ? tmp2471 : tmp973;
  assign tmp2604 = s0 ? tmp2601 : tmp2605;
  assign tmp2602 = s1 ? tmp2603 : tmp2604;
  assign tmp2598 = s2 ? tmp2599 : tmp2602;
  assign tmp2593 = s3 ? tmp2594 : tmp2598;
  assign tmp2610 = l1 ? tmp116 : tmp973;
  assign tmp2609 = s0 ? tmp2610 : 1;
  assign tmp2611 = s0 ? tmp2605 : tmp2601;
  assign tmp2608 = s1 ? tmp2609 : tmp2611;
  assign tmp2613 = s0 ? tmp2595 : 1;
  assign tmp2612 = s1 ? tmp2613 : tmp1944;
  assign tmp2607 = s2 ? tmp2608 : tmp2612;
  assign tmp2617 = l1 ? tmp2485 : tmp981;
  assign tmp2616 = s0 ? tmp2601 : tmp2617;
  assign tmp2618 = s0 ? tmp2547 : tmp2601;
  assign tmp2615 = s1 ? tmp2616 : tmp2618;
  assign tmp2614 = s2 ? tmp2542 : tmp2615;
  assign tmp2606 = s3 ? tmp2607 : tmp2614;
  assign tmp2592 = s4 ? tmp2593 : tmp2606;
  assign tmp2624 = s0 ? tmp2597 : 1;
  assign tmp2625 = l1 ? tmp116 : tmp74;
  assign tmp2623 = s1 ? tmp2624 : tmp2625;
  assign tmp2627 = l1 ? tmp109 : tmp1011;
  assign tmp2628 = s0 ? tmp2617 : 1;
  assign tmp2626 = s1 ? tmp2627 : tmp2628;
  assign tmp2622 = s2 ? tmp2623 : tmp2626;
  assign tmp2632 = ~(l2 ? tmp17 : tmp19);
  assign tmp2631 = l1 ? tmp898 : tmp2632;
  assign tmp2633 = ~(l1 ? tmp117 : tmp1021);
  assign tmp2630 = s1 ? tmp2631 : tmp2633;
  assign tmp2636 = l1 ? tmp2471 : tmp1021;
  assign tmp2637 = l1 ? tmp2485 : tmp1021;
  assign tmp2635 = s0 ? tmp2636 : tmp2637;
  assign tmp2634 = ~(s1 ? tmp2563 : tmp2635);
  assign tmp2629 = ~(s2 ? tmp2630 : tmp2634);
  assign tmp2621 = s3 ? tmp2622 : tmp2629;
  assign tmp2642 = l1 ? tmp2471 : tmp1011;
  assign tmp2641 = s0 ? tmp2433 : tmp2642;
  assign tmp2640 = s1 ? tmp2641 : tmp2568;
  assign tmp2643 = l1 ? tmp116 : tmp1011;
  assign tmp2639 = s2 ? tmp2640 : tmp2643;
  assign tmp2648 = ~(l2 ? tmp17 : tmp21);
  assign tmp2647 = l1 ? tmp31 : tmp2648;
  assign tmp2649 = ~(l1 ? tmp2485 : tmp1011);
  assign tmp2646 = s0 ? tmp2647 : tmp2649;
  assign tmp2645 = s1 ? tmp2646 : tmp2423;
  assign tmp2644 = ~(s2 ? tmp2645 : tmp2441);
  assign tmp2638 = s3 ? tmp2639 : tmp2644;
  assign tmp2620 = s4 ? tmp2621 : tmp2638;
  assign tmp2655 = l1 ? tmp117 : tmp1021;
  assign tmp2654 = s0 ? tmp2655 : tmp31;
  assign tmp2653 = s1 ? tmp2654 : tmp830;
  assign tmp2652 = s2 ? tmp2653 : tmp2447;
  assign tmp2651 = s3 ? tmp2652 : tmp2448;
  assign tmp2658 = l1 ? tmp74 : tmp2648;
  assign tmp2657 = s2 ? tmp2584 : tmp2658;
  assign tmp2656 = ~(s3 ? tmp2657 : tmp2457);
  assign tmp2650 = s4 ? tmp2651 : tmp2656;
  assign tmp2619 = s5 ? tmp2620 : tmp2650;
  assign tmp2591 = ~(s6 ? tmp2592 : tmp2619);
  assign tmp2590 = s7 ? 1 : tmp2591;
  assign tmp2589 = s8 ? tmp2590 : 1;
  assign tmp2661 = s6 ? tmp2383 : tmp2411;
  assign tmp2662 = s6 ? tmp2520 : tmp2548;
  assign tmp2660 = s7 ? tmp2661 : tmp2662;
  assign tmp2664 = s6 ? tmp2460 : tmp2487;
  assign tmp2665 = s6 ? tmp2592 : tmp2619;
  assign tmp2663 = s7 ? tmp2664 : tmp2665;
  assign tmp2659 = ~(s8 ? tmp2660 : tmp2663);
  assign tmp2588 = s9 ? tmp2589 : tmp2659;
  assign tmp2378 = s10 ? tmp2379 : tmp2588;
  assign tmp2166 = s12 ? tmp2167 : tmp2378;
  assign tmp2674 = l1 ? 1 : tmp966;
  assign tmp2677 = l2 ? 1 : tmp780;
  assign tmp2676 = l1 ? tmp2677 : tmp966;
  assign tmp2675 = s0 ? 1 : tmp2676;
  assign tmp2673 = s1 ? tmp2674 : tmp2675;
  assign tmp2679 = s1 ? 1 : tmp2676;
  assign tmp2678 = s2 ? tmp2675 : tmp2679;
  assign tmp2672 = s3 ? tmp2673 : tmp2678;
  assign tmp2683 = s0 ? tmp2674 : 1;
  assign tmp2682 = s1 ? tmp2683 : tmp2676;
  assign tmp2684 = s1 ? tmp2683 : 1;
  assign tmp2681 = s2 ? tmp2682 : tmp2684;
  assign tmp2686 = s1 ? 1 : tmp1749;
  assign tmp2688 = s0 ? tmp1722 : tmp2676;
  assign tmp2687 = s1 ? tmp2676 : tmp2688;
  assign tmp2685 = s2 ? tmp2686 : tmp2687;
  assign tmp2680 = s3 ? tmp2681 : tmp2685;
  assign tmp2671 = s4 ? tmp2672 : tmp2680;
  assign tmp2694 = s0 ? tmp2676 : 1;
  assign tmp2693 = s1 ? tmp2694 : 1;
  assign tmp2695 = s1 ? tmp2676 : tmp2694;
  assign tmp2692 = s2 ? tmp2693 : tmp2695;
  assign tmp2698 = l1 ? tmp2677 : tmp1123;
  assign tmp2697 = s1 ? 1 : tmp2698;
  assign tmp2700 = s0 ? tmp1722 : tmp1749;
  assign tmp2699 = s1 ? tmp2700 : tmp2698;
  assign tmp2696 = s2 ? tmp2697 : tmp2699;
  assign tmp2691 = s3 ? tmp2692 : tmp2696;
  assign tmp2704 = s0 ? tmp131 : tmp2698;
  assign tmp2703 = s1 ? tmp2704 : 1;
  assign tmp2702 = s2 ? tmp2703 : tmp2674;
  assign tmp2708 = l1 ? 1 : tmp1123;
  assign tmp2707 = s0 ? tmp2674 : tmp2708;
  assign tmp2706 = s1 ? tmp2707 : tmp2698;
  assign tmp2709 = s1 ? tmp31 : tmp1749;
  assign tmp2705 = s2 ? tmp2706 : tmp2709;
  assign tmp2701 = s3 ? tmp2702 : tmp2705;
  assign tmp2690 = s4 ? tmp2691 : tmp2701;
  assign tmp2714 = s0 ? tmp2698 : 1;
  assign tmp2713 = s1 ? tmp2714 : 1;
  assign tmp2712 = s2 ? tmp2713 : 1;
  assign tmp2716 = ~(s1 ? tmp131 : tmp966);
  assign tmp2715 = ~(s2 ? tmp1741 : tmp2716);
  assign tmp2711 = s3 ? tmp2712 : tmp2715;
  assign tmp2719 = s1 ? tmp618 : tmp1722;
  assign tmp2718 = s2 ? tmp2719 : tmp2676;
  assign tmp2720 = s1 ? tmp1722 : tmp2698;
  assign tmp2717 = s3 ? tmp2718 : tmp2720;
  assign tmp2710 = s4 ? tmp2711 : tmp2717;
  assign tmp2689 = s5 ? tmp2690 : tmp2710;
  assign tmp2670 = ~(s6 ? tmp2671 : tmp2689);
  assign tmp2669 = s7 ? 1 : tmp2670;
  assign tmp2728 = l2 ? 1 : tmp120;
  assign tmp2727 = l1 ? 1 : tmp2728;
  assign tmp2730 = l1 ? tmp2677 : tmp74;
  assign tmp2729 = s0 ? 1 : tmp2730;
  assign tmp2726 = s1 ? tmp2727 : tmp2729;
  assign tmp2733 = l1 ? tmp2677 : tmp2728;
  assign tmp2732 = s0 ? 1 : tmp2733;
  assign tmp2734 = s1 ? 1 : tmp2733;
  assign tmp2731 = s2 ? tmp2732 : tmp2734;
  assign tmp2725 = s3 ? tmp2726 : tmp2731;
  assign tmp2739 = l1 ? 1 : tmp74;
  assign tmp2738 = s0 ? tmp2739 : 1;
  assign tmp2737 = s1 ? tmp2738 : tmp2733;
  assign tmp2741 = s0 ? tmp2727 : 1;
  assign tmp2740 = s1 ? tmp2741 : 1;
  assign tmp2736 = s2 ? tmp2737 : tmp2740;
  assign tmp2744 = s0 ? tmp1722 : tmp2733;
  assign tmp2743 = s1 ? tmp2733 : tmp2744;
  assign tmp2742 = s2 ? tmp2686 : tmp2743;
  assign tmp2735 = s3 ? tmp2736 : tmp2742;
  assign tmp2724 = s4 ? tmp2725 : tmp2735;
  assign tmp2750 = s0 ? tmp2730 : 1;
  assign tmp2749 = s1 ? tmp2750 : 1;
  assign tmp2752 = l1 ? tmp2677 : tmp31;
  assign tmp2753 = s0 ? tmp2733 : 1;
  assign tmp2751 = s1 ? tmp2752 : tmp2753;
  assign tmp2748 = s2 ? tmp2749 : tmp2751;
  assign tmp2755 = s1 ? 1 : tmp2752;
  assign tmp2756 = s1 ? tmp2700 : tmp2752;
  assign tmp2754 = s2 ? tmp2755 : tmp2756;
  assign tmp2747 = s3 ? tmp2748 : tmp2754;
  assign tmp2760 = s0 ? tmp131 : tmp2752;
  assign tmp2759 = s1 ? tmp2760 : 1;
  assign tmp2758 = s2 ? tmp2759 : tmp131;
  assign tmp2762 = s1 ? tmp131 : tmp2752;
  assign tmp2761 = s2 ? tmp2762 : tmp2709;
  assign tmp2757 = s3 ? tmp2758 : tmp2761;
  assign tmp2746 = s4 ? tmp2747 : tmp2757;
  assign tmp2767 = s0 ? tmp2752 : 1;
  assign tmp2766 = s1 ? tmp2767 : 1;
  assign tmp2765 = s2 ? tmp2766 : 1;
  assign tmp2768 = ~(s2 ? tmp1741 : tmp41);
  assign tmp2764 = s3 ? tmp2765 : tmp2768;
  assign tmp2770 = s2 ? tmp2719 : tmp2752;
  assign tmp2771 = s1 ? tmp1722 : tmp2752;
  assign tmp2769 = s3 ? tmp2770 : tmp2771;
  assign tmp2763 = s4 ? tmp2764 : tmp2769;
  assign tmp2745 = s5 ? tmp2746 : tmp2763;
  assign tmp2723 = ~(s6 ? tmp2724 : tmp2745);
  assign tmp2722 = s7 ? 1 : tmp2723;
  assign tmp2721 = s8 ? tmp2669 : tmp2722;
  assign tmp2668 = s9 ? tmp2669 : tmp2721;
  assign tmp2773 = s8 ? tmp2669 : 1;
  assign tmp2776 = s6 ? tmp2671 : tmp2689;
  assign tmp2777 = s6 ? tmp2724 : tmp2745;
  assign tmp2775 = s7 ? tmp2776 : tmp2777;
  assign tmp2774 = ~(s8 ? tmp2775 : tmp2776);
  assign tmp2772 = s9 ? tmp2773 : tmp2774;
  assign tmp2667 = s10 ? tmp2668 : tmp2772;
  assign tmp2786 = l1 ? tmp81 : tmp74;
  assign tmp2787 = ~(l1 ? tmp26 : tmp323);
  assign tmp2785 = s1 ? tmp2786 : tmp2787;
  assign tmp2791 = ~(l1 ? tmp81 : tmp74);
  assign tmp2790 = s0 ? tmp208 : tmp2791;
  assign tmp2793 = l1 ? tmp26 : tmp323;
  assign tmp2792 = s0 ? tmp2793 : tmp2791;
  assign tmp2789 = s1 ? tmp2790 : tmp2792;
  assign tmp2795 = s0 ? tmp2793 : 0;
  assign tmp2794 = s1 ? tmp2795 : tmp2791;
  assign tmp2788 = ~(s2 ? tmp2789 : tmp2794);
  assign tmp2784 = s3 ? tmp2785 : tmp2788;
  assign tmp2799 = s0 ? tmp2130 : 0;
  assign tmp2798 = s1 ? tmp2799 : tmp2791;
  assign tmp2801 = s0 ? tmp2786 : 1;
  assign tmp2800 = ~(s1 ? tmp2801 : 1);
  assign tmp2797 = s2 ? tmp2798 : tmp2800;
  assign tmp2804 = l1 ? tmp31 : tmp74;
  assign tmp2803 = s1 ? 1 : tmp2804;
  assign tmp2807 = l1 ? tmp45 : tmp74;
  assign tmp2806 = s0 ? tmp2786 : tmp2807;
  assign tmp2809 = l1 ? tmp24 : tmp74;
  assign tmp2808 = s0 ? tmp2809 : tmp2786;
  assign tmp2805 = s1 ? tmp2806 : tmp2808;
  assign tmp2802 = ~(s2 ? tmp2803 : tmp2805);
  assign tmp2796 = ~(s3 ? tmp2797 : tmp2802);
  assign tmp2783 = s4 ? tmp2784 : tmp2796;
  assign tmp2814 = s1 ? tmp2795 : tmp208;
  assign tmp2816 = l1 ? tmp26 : tmp203;
  assign tmp2817 = ~(s0 ? tmp2807 : 1);
  assign tmp2815 = s1 ? tmp2816 : tmp2817;
  assign tmp2813 = s2 ? tmp2814 : tmp2815;
  assign tmp2820 = l1 ? tmp74 : tmp323;
  assign tmp2821 = ~(l1 ? tmp45 : tmp74);
  assign tmp2819 = s1 ? tmp2820 : tmp2821;
  assign tmp2823 = s0 ? tmp2809 : tmp207;
  assign tmp2822 = ~(s1 ? tmp2823 : tmp2806);
  assign tmp2818 = s2 ? tmp2819 : tmp2822;
  assign tmp2812 = s3 ? tmp2813 : tmp2818;
  assign tmp2827 = s0 ? tmp2804 : tmp2786;
  assign tmp2826 = s1 ? tmp2827 : 1;
  assign tmp2828 = ~(l1 ? tmp31 : tmp203);
  assign tmp2825 = s2 ? tmp2826 : tmp2828;
  assign tmp2832 = ~(l1 ? tmp117 : tmp74);
  assign tmp2831 = s0 ? tmp202 : tmp2832;
  assign tmp2830 = s1 ? tmp2831 : tmp2821;
  assign tmp2833 = ~(s1 ? 1 : tmp2804);
  assign tmp2829 = ~(s2 ? tmp2830 : tmp2833);
  assign tmp2824 = ~(s3 ? tmp2825 : tmp2829);
  assign tmp2811 = s4 ? tmp2812 : tmp2824;
  assign tmp2838 = s0 ? tmp2807 : tmp31;
  assign tmp2837 = s1 ? tmp2838 : tmp54;
  assign tmp2836 = s2 ? tmp2837 : tmp2447;
  assign tmp2840 = s1 ? tmp355 : tmp83;
  assign tmp2841 = ~(s1 ? tmp2804 : tmp2828);
  assign tmp2839 = ~(s2 ? tmp2840 : tmp2841);
  assign tmp2835 = s3 ? tmp2836 : tmp2839;
  assign tmp2845 = ~(l1 ? tmp24 : tmp74);
  assign tmp2844 = s1 ? 1 : tmp2845;
  assign tmp2846 = l1 ? tmp901 : tmp203;
  assign tmp2843 = s2 ? tmp2844 : tmp2846;
  assign tmp2847 = s1 ? tmp355 : tmp2821;
  assign tmp2842 = ~(s3 ? tmp2843 : tmp2847);
  assign tmp2834 = ~(s4 ? tmp2835 : tmp2842);
  assign tmp2810 = ~(s5 ? tmp2811 : tmp2834);
  assign tmp2782 = ~(s6 ? tmp2783 : tmp2810);
  assign tmp2781 = s7 ? 1 : tmp2782;
  assign tmp2853 = l1 ? tmp2464 : tmp1504;
  assign tmp2854 = l1 ? tmp17 : tmp1504;
  assign tmp2852 = s1 ? tmp2853 : tmp2854;
  assign tmp2857 = s0 ? tmp2493 : tmp2853;
  assign tmp2858 = s0 ? tmp2854 : tmp2853;
  assign tmp2856 = s1 ? tmp2857 : tmp2858;
  assign tmp2860 = s0 ? tmp2854 : tmp135;
  assign tmp2859 = s1 ? tmp2860 : tmp2853;
  assign tmp2855 = s2 ? tmp2856 : tmp2859;
  assign tmp2851 = s3 ? tmp2852 : tmp2855;
  assign tmp2865 = l1 ? tmp116 : tmp1504;
  assign tmp2864 = s0 ? tmp2865 : 1;
  assign tmp2863 = s1 ? tmp2864 : tmp2853;
  assign tmp2867 = s0 ? tmp2853 : 1;
  assign tmp2868 = l1 ? 1 : tmp898;
  assign tmp2866 = s1 ? tmp2867 : tmp2868;
  assign tmp2862 = s2 ? tmp2863 : tmp2866;
  assign tmp2871 = l1 ? 1 : tmp1496;
  assign tmp2870 = s1 ? tmp2871 : tmp2804;
  assign tmp2875 = l2 ? tmp780 : tmp20;
  assign tmp2874 = l1 ? tmp2875 : tmp1504;
  assign tmp2873 = s0 ? tmp2853 : tmp2874;
  assign tmp2878 = ~(l2 ? tmp17 : tmp33);
  assign tmp2877 = l1 ? tmp24 : tmp2878;
  assign tmp2876 = s0 ? tmp2877 : tmp2853;
  assign tmp2872 = s1 ? tmp2873 : tmp2876;
  assign tmp2869 = s2 ? tmp2870 : tmp2872;
  assign tmp2861 = s3 ? tmp2862 : tmp2869;
  assign tmp2850 = s4 ? tmp2851 : tmp2861;
  assign tmp2884 = s0 ? tmp2854 : 1;
  assign tmp2883 = s1 ? tmp2884 : tmp2493;
  assign tmp2887 = l2 ? tmp898 : 0;
  assign tmp2886 = l1 ? tmp17 : tmp2887;
  assign tmp2888 = s0 ? tmp2874 : tmp135;
  assign tmp2885 = s1 ? tmp2886 : tmp2888;
  assign tmp2882 = s2 ? tmp2883 : tmp2885;
  assign tmp2892 = ~(l2 ? tmp898 : tmp19);
  assign tmp2891 = l1 ? tmp898 : tmp2892;
  assign tmp2893 = ~(l1 ? tmp45 : tmp1504);
  assign tmp2890 = s1 ? tmp2891 : tmp2893;
  assign tmp2895 = s0 ? tmp2877 : tmp207;
  assign tmp2897 = l1 ? tmp2875 : tmp2878;
  assign tmp2896 = s0 ? tmp2853 : tmp2897;
  assign tmp2894 = ~(s1 ? tmp2895 : tmp2896);
  assign tmp2889 = ~(s2 ? tmp2890 : tmp2894);
  assign tmp2881 = s3 ? tmp2882 : tmp2889;
  assign tmp2901 = s0 ? tmp2804 : tmp2853;
  assign tmp2902 = s0 ? 1 : tmp822;
  assign tmp2900 = s1 ? tmp2901 : tmp2902;
  assign tmp2903 = l1 ? tmp116 : tmp2887;
  assign tmp2899 = s2 ? tmp2900 : tmp2903;
  assign tmp2908 = ~(l2 ? tmp898 : 0);
  assign tmp2907 = l1 ? tmp31 : tmp2908;
  assign tmp2909 = ~(l1 ? tmp2485 : tmp2878);
  assign tmp2906 = s0 ? tmp2907 : tmp2909;
  assign tmp2905 = s1 ? tmp2906 : tmp2821;
  assign tmp2904 = ~(s2 ? tmp2905 : tmp2833);
  assign tmp2898 = s3 ? tmp2899 : tmp2904;
  assign tmp2880 = s4 ? tmp2881 : tmp2898;
  assign tmp2915 = l1 ? tmp45 : tmp1504;
  assign tmp2914 = s0 ? tmp2915 : tmp31;
  assign tmp2913 = s1 ? tmp2914 : tmp1039;
  assign tmp2912 = s2 ? tmp2913 : tmp2516;
  assign tmp2911 = s3 ? tmp2912 : tmp2839;
  assign tmp2919 = ~(l1 ? tmp24 : tmp2878);
  assign tmp2918 = s1 ? 1 : tmp2919;
  assign tmp2920 = l1 ? tmp901 : tmp2908;
  assign tmp2917 = s2 ? tmp2918 : tmp2920;
  assign tmp2916 = ~(s3 ? tmp2917 : tmp2847);
  assign tmp2910 = s4 ? tmp2911 : tmp2916;
  assign tmp2879 = s5 ? tmp2880 : tmp2910;
  assign tmp2849 = ~(s6 ? tmp2850 : tmp2879);
  assign tmp2848 = s7 ? 1 : tmp2849;
  assign tmp2780 = s8 ? tmp2781 : tmp2848;
  assign tmp2927 = l1 ? tmp2464 : tmp74;
  assign tmp2928 = l1 ? tmp17 : tmp74;
  assign tmp2926 = s1 ? tmp2927 : tmp2928;
  assign tmp2931 = s0 ? tmp2554 : tmp2927;
  assign tmp2933 = l1 ? tmp17 : 1;
  assign tmp2932 = s0 ? tmp2933 : tmp2927;
  assign tmp2930 = s1 ? tmp2931 : tmp2932;
  assign tmp2935 = s0 ? tmp2933 : 1;
  assign tmp2934 = s1 ? tmp2935 : tmp2927;
  assign tmp2929 = s2 ? tmp2930 : tmp2934;
  assign tmp2925 = s3 ? tmp2926 : tmp2929;
  assign tmp2939 = s0 ? tmp2625 : 1;
  assign tmp2938 = s1 ? tmp2939 : tmp2927;
  assign tmp2941 = s0 ? tmp2927 : 1;
  assign tmp2940 = s1 ? tmp2941 : 1;
  assign tmp2937 = s2 ? tmp2938 : tmp2940;
  assign tmp2945 = l1 ? tmp2875 : tmp74;
  assign tmp2944 = s0 ? tmp2927 : tmp2945;
  assign tmp2946 = s0 ? tmp2809 : tmp2927;
  assign tmp2943 = s1 ? tmp2944 : tmp2946;
  assign tmp2942 = s2 ? tmp2803 : tmp2943;
  assign tmp2936 = s3 ? tmp2937 : tmp2942;
  assign tmp2924 = s4 ? tmp2925 : tmp2936;
  assign tmp2952 = s0 ? tmp2928 : 1;
  assign tmp2951 = s1 ? tmp2952 : tmp2554;
  assign tmp2954 = l1 ? tmp17 : tmp31;
  assign tmp2955 = s0 ? tmp2945 : 1;
  assign tmp2953 = s1 ? tmp2954 : tmp2955;
  assign tmp2950 = s2 ? tmp2951 : tmp2953;
  assign tmp2958 = l1 ? tmp898 : 0;
  assign tmp2957 = s1 ? tmp2958 : tmp2821;
  assign tmp2959 = ~(s1 ? tmp2823 : tmp2944);
  assign tmp2956 = ~(s2 ? tmp2957 : tmp2959);
  assign tmp2949 = s3 ? tmp2950 : tmp2956;
  assign tmp2963 = s0 ? tmp2804 : tmp2927;
  assign tmp2962 = s1 ? tmp2963 : 1;
  assign tmp2964 = l1 ? tmp116 : tmp31;
  assign tmp2961 = s2 ? tmp2962 : tmp2964;
  assign tmp2968 = ~(l1 ? tmp2485 : tmp74);
  assign tmp2967 = s0 ? tmp202 : tmp2968;
  assign tmp2966 = s1 ? tmp2967 : tmp2821;
  assign tmp2965 = ~(s2 ? tmp2966 : tmp2833);
  assign tmp2960 = s3 ? tmp2961 : tmp2965;
  assign tmp2948 = s4 ? tmp2949 : tmp2960;
  assign tmp2971 = s2 ? tmp2837 : tmp2579;
  assign tmp2970 = s3 ? tmp2971 : tmp2839;
  assign tmp2969 = s4 ? tmp2970 : tmp2842;
  assign tmp2947 = s5 ? tmp2948 : tmp2969;
  assign tmp2923 = ~(s6 ? tmp2924 : tmp2947);
  assign tmp2922 = s7 ? 1 : tmp2923;
  assign tmp2921 = s8 ? tmp2848 : tmp2922;
  assign tmp2779 = s9 ? tmp2780 : tmp2921;
  assign tmp2980 = s0 ? tmp2625 : tmp2927;
  assign tmp2981 = s0 ? tmp2928 : tmp2927;
  assign tmp2979 = s1 ? tmp2980 : tmp2981;
  assign tmp2982 = s1 ? tmp2952 : tmp2927;
  assign tmp2978 = s2 ? tmp2979 : tmp2982;
  assign tmp2977 = s3 ? tmp2926 : tmp2978;
  assign tmp2976 = s4 ? tmp2977 : tmp2936;
  assign tmp2987 = s1 ? tmp2952 : tmp2625;
  assign tmp2986 = s2 ? tmp2987 : tmp2953;
  assign tmp2990 = l1 ? tmp898 : tmp323;
  assign tmp2989 = s1 ? tmp2990 : tmp2821;
  assign tmp2988 = ~(s2 ? tmp2989 : tmp2959);
  assign tmp2985 = s3 ? tmp2986 : tmp2988;
  assign tmp2984 = s4 ? tmp2985 : tmp2960;
  assign tmp2991 = s4 ? tmp2835 : tmp2842;
  assign tmp2983 = s5 ? tmp2984 : tmp2991;
  assign tmp2975 = ~(s6 ? tmp2976 : tmp2983);
  assign tmp2974 = s7 ? 1 : tmp2975;
  assign tmp2973 = s8 ? tmp2974 : 1;
  assign tmp2994 = s6 ? tmp2783 : tmp2810;
  assign tmp2995 = s6 ? tmp2924 : tmp2947;
  assign tmp2993 = s7 ? tmp2994 : tmp2995;
  assign tmp2997 = s6 ? tmp2850 : tmp2879;
  assign tmp2998 = s6 ? tmp2976 : tmp2983;
  assign tmp2996 = s7 ? tmp2997 : tmp2998;
  assign tmp2992 = ~(s8 ? tmp2993 : tmp2996);
  assign tmp2972 = s9 ? tmp2973 : tmp2992;
  assign tmp2778 = s10 ? tmp2779 : tmp2972;
  assign tmp2666 = s12 ? tmp2667 : tmp2778;
  assign tmp2165 = s13 ? tmp2166 : tmp2666;
  assign tmp1670 = s14 ? tmp1671 : tmp2165;
  assign tmp3 = s15 ? tmp4 : tmp1670;
  assign tmp3003 = s9 ? tmp8 : tmp103;
  assign tmp3005 = s8 ? tmp103 : 1;
  assign tmp3012 = l1 ? tmp109 : tmp24;
  assign tmp3014 = l1 ? tmp17 : tmp24;
  assign tmp3013 = s0 ? tmp23 : tmp3014;
  assign tmp3011 = s1 ? tmp3012 : tmp3013;
  assign tmp3018 = l1 ? tmp116 : tmp24;
  assign tmp3017 = s0 ? tmp3018 : tmp243;
  assign tmp3019 = s0 ? tmp3012 : tmp243;
  assign tmp3016 = s1 ? tmp3017 : tmp3019;
  assign tmp3021 = s0 ? tmp3012 : tmp23;
  assign tmp3022 = s0 ? tmp243 : tmp3014;
  assign tmp3020 = s1 ? tmp3021 : tmp3022;
  assign tmp3015 = s2 ? tmp3016 : tmp3020;
  assign tmp3010 = s3 ? tmp3011 : tmp3015;
  assign tmp3026 = s0 ? tmp3018 : tmp131;
  assign tmp3027 = s0 ? tmp3014 : tmp243;
  assign tmp3025 = s1 ? tmp3026 : tmp3027;
  assign tmp3029 = s0 ? tmp3012 : tmp83;
  assign tmp3028 = s1 ? tmp3029 : tmp135;
  assign tmp3024 = s2 ? tmp3025 : tmp3028;
  assign tmp3032 = ~(s0 ? 1 : tmp225);
  assign tmp3031 = s1 ? tmp243 : tmp3032;
  assign tmp3030 = s2 ? tmp57 : tmp3031;
  assign tmp3023 = s3 ? tmp3024 : tmp3030;
  assign tmp3009 = s4 ? tmp3010 : tmp3023;
  assign tmp3038 = s0 ? tmp3014 : tmp131;
  assign tmp3037 = s1 ? tmp3038 : tmp3018;
  assign tmp3040 = s0 ? tmp243 : tmp23;
  assign tmp3039 = s1 ? tmp3014 : tmp3040;
  assign tmp3036 = s2 ? tmp3037 : tmp3039;
  assign tmp3043 = l1 ? tmp152 : tmp24;
  assign tmp3042 = s1 ? tmp3043 : tmp243;
  assign tmp3044 = ~(s1 ? 1 : tmp225);
  assign tmp3041 = s2 ? tmp3042 : tmp3044;
  assign tmp3035 = s3 ? tmp3036 : tmp3041;
  assign tmp3049 = ~(l1 ? tmp17 : tmp24);
  assign tmp3048 = s0 ? 1 : tmp3049;
  assign tmp3047 = s1 ? tmp3048 : tmp82;
  assign tmp3050 = ~(l1 ? tmp116 : tmp24);
  assign tmp3046 = s2 ? tmp3047 : tmp3050;
  assign tmp3054 = ~(l1 ? tmp152 : 0);
  assign tmp3053 = s0 ? tmp187 : tmp3054;
  assign tmp3052 = s1 ? tmp3053 : tmp21;
  assign tmp3051 = s2 ? tmp3052 : 1;
  assign tmp3045 = ~(s3 ? tmp3046 : tmp3051);
  assign tmp3034 = s4 ? tmp3035 : tmp3045;
  assign tmp3055 = s4 ? tmp239 : tmp247;
  assign tmp3033 = s5 ? tmp3034 : tmp3055;
  assign tmp3008 = ~(s6 ? tmp3009 : tmp3033);
  assign tmp3007 = s7 ? tmp298 : tmp3008;
  assign tmp3056 = ~(s6 ? tmp105 : tmp140);
  assign tmp3006 = ~(s8 ? tmp3007 : tmp3056);
  assign tmp3004 = s9 ? tmp3005 : tmp3006;
  assign tmp3002 = s10 ? tmp3003 : tmp3004;
  assign tmp3066 = l1 ? tmp330 : tmp102;
  assign tmp3065 = s1 ? tmp3066 : tmp602;
  assign tmp3070 = l1 ? tmp392 : tmp203;
  assign tmp3069 = s0 ? tmp3070 : tmp3066;
  assign tmp3072 = l1 ? tmp330 : tmp203;
  assign tmp3071 = s0 ? tmp3072 : tmp3066;
  assign tmp3068 = s1 ? tmp3069 : tmp3071;
  assign tmp3074 = s0 ? tmp3072 : tmp375;
  assign tmp3073 = s1 ? tmp3074 : tmp3066;
  assign tmp3067 = s2 ? tmp3068 : tmp3073;
  assign tmp3064 = s3 ? tmp3065 : tmp3067;
  assign tmp3077 = s1 ? tmp615 : tmp3066;
  assign tmp3079 = s0 ? tmp3066 : 1;
  assign tmp3078 = s1 ? tmp3079 : tmp618;
  assign tmp3076 = s2 ? tmp3077 : tmp3078;
  assign tmp3083 = ~(l1 ? tmp330 : tmp102);
  assign tmp3082 = ~(s0 ? 1 : tmp3083);
  assign tmp3081 = s1 ? tmp3066 : tmp3082;
  assign tmp3080 = s2 ? tmp620 : tmp3081;
  assign tmp3075 = s3 ? tmp3076 : tmp3080;
  assign tmp3063 = s4 ? tmp3064 : tmp3075;
  assign tmp3088 = s1 ? tmp611 : tmp3070;
  assign tmp3091 = l1 ? tmp373 : tmp102;
  assign tmp3090 = s0 ? tmp3091 : tmp375;
  assign tmp3089 = s1 ? tmp630 : tmp3090;
  assign tmp3087 = s2 ? tmp3088 : tmp3089;
  assign tmp3094 = l1 ? tmp373 : tmp203;
  assign tmp3093 = s1 ? tmp3094 : 0;
  assign tmp3092 = s2 ? tmp3093 : tmp636;
  assign tmp3086 = s3 ? tmp3087 : tmp3092;
  assign tmp3085 = s4 ? tmp3086 : tmp639;
  assign tmp3084 = s5 ? tmp3085 : 0;
  assign tmp3062 = s6 ? tmp3063 : tmp3084;
  assign tmp3061 = s7 ? 1 : tmp3062;
  assign tmp3060 = s8 ? tmp595 : tmp3061;
  assign tmp3059 = s9 ? tmp545 : tmp3060;
  assign tmp3096 = s8 ? tmp595 : 1;
  assign tmp3099 = ~(s6 ? tmp3063 : tmp3084);
  assign tmp3098 = s7 ? tmp723 : tmp3099;
  assign tmp3100 = ~(s6 ? tmp597 : tmp624);
  assign tmp3097 = ~(s8 ? tmp3098 : tmp3100);
  assign tmp3095 = s9 ? tmp3096 : tmp3097;
  assign tmp3058 = s10 ? tmp3059 : tmp3095;
  assign tmp3057 = s12 ? tmp302 : tmp3058;
  assign tmp3001 = s13 ? tmp3002 : tmp3057;
  assign tmp3111 = l2 ? tmp780 : tmp120;
  assign tmp3110 = l1 ? tmp373 : tmp3111;
  assign tmp3113 = l1 ? tmp31 : tmp1002;
  assign tmp3114 = l1 ? tmp373 : tmp1202;
  assign tmp3112 = s0 ? tmp3113 : tmp3114;
  assign tmp3109 = s1 ? tmp3110 : tmp3112;
  assign tmp3118 = l1 ? tmp373 : tmp74;
  assign tmp3119 = l1 ? tmp373 : tmp330;
  assign tmp3117 = s0 ? tmp3118 : tmp3119;
  assign tmp3120 = s0 ? tmp3114 : tmp3119;
  assign tmp3116 = s1 ? tmp3117 : tmp3120;
  assign tmp3122 = s0 ? tmp3114 : tmp207;
  assign tmp3123 = s0 ? tmp3119 : tmp3110;
  assign tmp3121 = s1 ? tmp3122 : tmp3123;
  assign tmp3115 = s2 ? tmp3116 : tmp3121;
  assign tmp3108 = s3 ? tmp3109 : tmp3115;
  assign tmp3127 = s0 ? tmp3110 : tmp3119;
  assign tmp3126 = s1 ? tmp3122 : tmp3127;
  assign tmp3129 = s0 ? tmp3110 : tmp207;
  assign tmp3130 = l1 ? tmp31 : tmp780;
  assign tmp3128 = s1 ? tmp3129 : tmp3130;
  assign tmp3125 = s2 ? tmp3126 : tmp3128;
  assign tmp3132 = s1 ? tmp3113 : 0;
  assign tmp3134 = s0 ? tmp3119 : tmp330;
  assign tmp3135 = s0 ? tmp17 : tmp3119;
  assign tmp3133 = s1 ? tmp3134 : tmp3135;
  assign tmp3131 = s2 ? tmp3132 : tmp3133;
  assign tmp3124 = s3 ? tmp3125 : tmp3131;
  assign tmp3107 = s4 ? tmp3108 : tmp3124;
  assign tmp3141 = s0 ? tmp3114 : tmp54;
  assign tmp3140 = s1 ? tmp3141 : tmp3118;
  assign tmp3144 = l2 ? tmp780 : 0;
  assign tmp3143 = l1 ? tmp373 : tmp3144;
  assign tmp3145 = s0 ? tmp330 : 1;
  assign tmp3142 = s1 ? tmp3143 : tmp3145;
  assign tmp3139 = s2 ? tmp3140 : tmp3142;
  assign tmp3147 = s1 ? tmp3114 : tmp373;
  assign tmp3148 = s1 ? tmp93 : tmp373;
  assign tmp3146 = s2 ? tmp3147 : tmp3148;
  assign tmp3138 = s3 ? tmp3139 : tmp3146;
  assign tmp3153 = ~(l1 ? tmp373 : tmp3144);
  assign tmp3152 = s0 ? 1 : tmp3153;
  assign tmp3155 = l1 ? tmp31 : tmp17;
  assign tmp3154 = ~(s0 ? tmp207 : tmp3155);
  assign tmp3151 = s1 ? tmp3152 : tmp3154;
  assign tmp3150 = s2 ? tmp3151 : tmp3153;
  assign tmp3158 = s0 ? tmp810 : tmp356;
  assign tmp3157 = s1 ? tmp3158 : 1;
  assign tmp3156 = s2 ? tmp3157 : 1;
  assign tmp3149 = ~(s3 ? tmp3150 : tmp3156);
  assign tmp3137 = s4 ? tmp3138 : tmp3149;
  assign tmp3159 = s4 ? tmp827 : tmp831;
  assign tmp3136 = s5 ? tmp3137 : tmp3159;
  assign tmp3106 = s6 ? tmp3107 : tmp3136;
  assign tmp3105 = s7 ? 1 : tmp3106;
  assign tmp3166 = l1 ? tmp373 : tmp2464;
  assign tmp3168 = l1 ? tmp373 : tmp780;
  assign tmp3167 = s0 ? tmp3113 : tmp3168;
  assign tmp3165 = s1 ? tmp3166 : tmp3167;
  assign tmp3172 = l1 ? tmp373 : 1;
  assign tmp3173 = l1 ? tmp373 : tmp17;
  assign tmp3171 = s0 ? tmp3172 : tmp3173;
  assign tmp3175 = l1 ? tmp373 : tmp1002;
  assign tmp3174 = s0 ? tmp3175 : tmp3173;
  assign tmp3170 = s1 ? tmp3171 : tmp3174;
  assign tmp3177 = s0 ? tmp3175 : tmp207;
  assign tmp3178 = s0 ? tmp3173 : tmp3166;
  assign tmp3176 = s1 ? tmp3177 : tmp3178;
  assign tmp3169 = s2 ? tmp3170 : tmp3176;
  assign tmp3164 = s3 ? tmp3165 : tmp3169;
  assign tmp3182 = s0 ? tmp3168 : tmp207;
  assign tmp3183 = s0 ? tmp3166 : tmp3173;
  assign tmp3181 = s1 ? tmp3182 : tmp3183;
  assign tmp3185 = s0 ? tmp3166 : tmp207;
  assign tmp3184 = s1 ? tmp3185 : tmp3130;
  assign tmp3180 = s2 ? tmp3181 : tmp3184;
  assign tmp3188 = s0 ? tmp17 : tmp3173;
  assign tmp3187 = s1 ? tmp3173 : tmp3188;
  assign tmp3186 = s2 ? tmp3132 : tmp3187;
  assign tmp3179 = s3 ? tmp3180 : tmp3186;
  assign tmp3163 = s4 ? tmp3164 : tmp3179;
  assign tmp3194 = s0 ? tmp3168 : tmp54;
  assign tmp3193 = s1 ? tmp3194 : tmp3172;
  assign tmp3196 = s0 ? tmp3173 : 1;
  assign tmp3195 = s1 ? tmp3168 : tmp3196;
  assign tmp3192 = s2 ? tmp3193 : tmp3195;
  assign tmp3198 = s1 ? tmp3175 : tmp830;
  assign tmp3199 = s1 ? tmp93 : tmp3173;
  assign tmp3197 = s2 ? tmp3198 : tmp3199;
  assign tmp3191 = s3 ? tmp3192 : tmp3197;
  assign tmp3202 = ~(l1 ? tmp373 : tmp780);
  assign tmp3201 = s2 ? tmp3151 : tmp3202;
  assign tmp3205 = s0 ? tmp798 : tmp356;
  assign tmp3204 = s1 ? tmp3205 : 1;
  assign tmp3203 = s2 ? tmp3204 : 1;
  assign tmp3200 = ~(s3 ? tmp3201 : tmp3203);
  assign tmp3190 = s4 ? tmp3191 : tmp3200;
  assign tmp3206 = ~(s4 ? tmp874 : tmp879);
  assign tmp3189 = s5 ? tmp3190 : tmp3206;
  assign tmp3162 = s6 ? tmp3163 : tmp3189;
  assign tmp3161 = s7 ? 1 : tmp3162;
  assign tmp3160 = s8 ? tmp3105 : tmp3161;
  assign tmp3104 = s9 ? tmp3105 : tmp3160;
  assign tmp3208 = s8 ? tmp3105 : 1;
  assign tmp3211 = ~(s6 ? tmp3163 : tmp3189);
  assign tmp3210 = s7 ? tmp885 : tmp3211;
  assign tmp3212 = ~(s6 ? tmp3107 : tmp3136);
  assign tmp3209 = ~(s8 ? tmp3210 : tmp3212);
  assign tmp3207 = s9 ? tmp3208 : tmp3209;
  assign tmp3103 = s10 ? tmp3104 : tmp3207;
  assign tmp3219 = l1 ? tmp152 : tmp917;
  assign tmp3221 = l1 ? tmp35 : tmp917;
  assign tmp3220 = s0 ? tmp336 : tmp3221;
  assign tmp3218 = s1 ? tmp3219 : tmp3220;
  assign tmp3224 = l1 ? tmp152 : tmp33;
  assign tmp3223 = s0 ? tmp3224 : tmp3221;
  assign tmp3226 = s0 ? tmp3224 : tmp208;
  assign tmp3225 = s1 ? tmp3226 : tmp3221;
  assign tmp3222 = s2 ? tmp3223 : tmp3225;
  assign tmp3217 = s3 ? tmp3218 : tmp3222;
  assign tmp3231 = l1 ? tmp322 : 0;
  assign tmp3230 = s0 ? tmp3219 : tmp3231;
  assign tmp3229 = s1 ? tmp3230 : tmp3221;
  assign tmp3233 = s0 ? tmp3219 : tmp31;
  assign tmp3232 = s1 ? tmp3233 : tmp336;
  assign tmp3228 = s2 ? tmp3229 : tmp3232;
  assign tmp3235 = s1 ? tmp336 : tmp173;
  assign tmp3237 = s0 ? tmp3221 : tmp929;
  assign tmp3239 = ~(l1 ? tmp35 : tmp917);
  assign tmp3238 = ~(s0 ? tmp397 : tmp3239);
  assign tmp3236 = s1 ? tmp3237 : tmp3238;
  assign tmp3234 = s2 ? tmp3235 : tmp3236;
  assign tmp3227 = s3 ? tmp3228 : tmp3234;
  assign tmp3216 = s4 ? tmp3217 : tmp3227;
  assign tmp3245 = s0 ? tmp3221 : 0;
  assign tmp3244 = s1 ? tmp3245 : tmp3224;
  assign tmp3247 = l1 ? tmp35 : tmp933;
  assign tmp3248 = s0 ? tmp929 : tmp355;
  assign tmp3246 = s1 ? tmp3247 : tmp3248;
  assign tmp3243 = s2 ? tmp3244 : tmp3246;
  assign tmp3250 = s1 ? tmp3224 : tmp955;
  assign tmp3252 = ~(s0 ? tmp3247 : tmp955);
  assign tmp3251 = ~(s1 ? tmp935 : tmp3252);
  assign tmp3249 = s2 ? tmp3250 : tmp3251;
  assign tmp3242 = s3 ? tmp3243 : tmp3249;
  assign tmp3257 = ~(l1 ? tmp35 : tmp933);
  assign tmp3256 = s0 ? tmp397 : tmp3257;
  assign tmp3258 = ~(s0 ? tmp3231 : 1);
  assign tmp3255 = s1 ? tmp3256 : tmp3258;
  assign tmp3259 = ~(l1 ? tmp152 : tmp933);
  assign tmp3254 = s2 ? tmp3255 : tmp3259;
  assign tmp3263 = ~(l1 ? tmp152 : tmp966);
  assign tmp3262 = s0 ? tmp946 : tmp3263;
  assign tmp3261 = s1 ? tmp3262 : tmp932;
  assign tmp3260 = s2 ? tmp3261 : tmp949;
  assign tmp3253 = ~(s3 ? tmp3254 : tmp3260);
  assign tmp3241 = s4 ? tmp3242 : tmp3253;
  assign tmp3268 = l1 ? tmp31 : tmp24;
  assign tmp3267 = ~(s1 ? tmp3268 : tmp174);
  assign tmp3266 = s2 ? tmp953 : tmp3267;
  assign tmp3265 = s3 ? tmp3266 : tmp957;
  assign tmp3264 = s4 ? tmp3265 : tmp960;
  assign tmp3240 = s5 ? tmp3241 : tmp3264;
  assign tmp3215 = s6 ? tmp3216 : tmp3240;
  assign tmp3214 = s7 ? 1 : tmp3215;
  assign tmp3270 = s8 ? tmp3214 : 1;
  assign tmp3269 = s9 ? tmp3270 : tmp3215;
  assign tmp3213 = s10 ? tmp3214 : tmp3269;
  assign tmp3102 = s12 ? tmp3103 : tmp3213;
  assign tmp3273 = s9 ? tmp1113 : tmp1196;
  assign tmp3275 = s8 ? tmp1196 : 1;
  assign tmp3282 = l1 ? tmp1202 : tmp811;
  assign tmp3284 = l1 ? tmp973 : tmp811;
  assign tmp3283 = s0 ? tmp1205 : tmp3284;
  assign tmp3281 = s1 ? tmp3282 : tmp3283;
  assign tmp3288 = l1 ? tmp981 : tmp356;
  assign tmp3287 = s0 ? tmp3070 : tmp3288;
  assign tmp3290 = l1 ? tmp392 : tmp811;
  assign tmp3289 = s0 ? tmp3290 : tmp3288;
  assign tmp3286 = s1 ? tmp3287 : tmp3289;
  assign tmp3292 = s0 ? tmp3290 : tmp375;
  assign tmp3294 = l1 ? tmp981 : tmp811;
  assign tmp3293 = s0 ? tmp3288 : tmp3294;
  assign tmp3291 = s1 ? tmp3292 : tmp3293;
  assign tmp3285 = s2 ? tmp3286 : tmp3291;
  assign tmp3280 = s3 ? tmp3281 : tmp3285;
  assign tmp3298 = s0 ? tmp3290 : tmp603;
  assign tmp3299 = s0 ? tmp3294 : tmp3288;
  assign tmp3297 = s1 ? tmp3298 : tmp3299;
  assign tmp3301 = s0 ? tmp3282 : 1;
  assign tmp3300 = s1 ? tmp3301 : tmp1226;
  assign tmp3296 = s2 ? tmp3297 : tmp3300;
  assign tmp3305 = l1 ? tmp1021 : tmp356;
  assign tmp3304 = s0 ? tmp3288 : tmp3305;
  assign tmp3306 = s0 ? tmp1233 : tmp3288;
  assign tmp3303 = s1 ? tmp3304 : tmp3306;
  assign tmp3302 = s2 ? tmp1228 : tmp3303;
  assign tmp3295 = s3 ? tmp3296 : tmp3302;
  assign tmp3279 = s4 ? tmp3280 : tmp3295;
  assign tmp3312 = s0 ? tmp3284 : tmp203;
  assign tmp3311 = s1 ? tmp3312 : tmp3070;
  assign tmp3314 = s0 ? tmp3305 : tmp375;
  assign tmp3313 = s1 ? tmp1241 : tmp3314;
  assign tmp3310 = s2 ? tmp3311 : tmp3313;
  assign tmp3316 = s1 ? tmp3290 : tmp1169;
  assign tmp3315 = s2 ? tmp3316 : tmp1245;
  assign tmp3309 = s3 ? tmp3310 : tmp3315;
  assign tmp3320 = s0 ? 1 : tmp3294;
  assign tmp3319 = s1 ? tmp3320 : tmp1255;
  assign tmp3318 = s2 ? tmp3319 : tmp1256;
  assign tmp3324 = ~(l1 ? tmp1202 : tmp356);
  assign tmp3323 = s0 ? tmp1180 : tmp3324;
  assign tmp3322 = s1 ? tmp3323 : tmp1329;
  assign tmp3321 = ~(s2 ? tmp3322 : 0);
  assign tmp3317 = s3 ? tmp3318 : tmp3321;
  assign tmp3308 = s4 ? tmp3309 : tmp3317;
  assign tmp3326 = s3 ? tmp1263 : tmp1336;
  assign tmp3327 = ~(s3 ? tmp1267 : tmp1341);
  assign tmp3325 = s4 ? tmp3326 : tmp3327;
  assign tmp3307 = s5 ? tmp3308 : tmp3325;
  assign tmp3278 = s6 ? tmp3279 : tmp3307;
  assign tmp3277 = s7 ? tmp1414 : tmp3278;
  assign tmp3276 = ~(s8 ? tmp3277 : tmp1417);
  assign tmp3274 = s9 ? tmp3275 : tmp3276;
  assign tmp3272 = s10 ? tmp3273 : tmp3274;
  assign tmp3271 = s12 ? tmp3272 : tmp1419;
  assign tmp3101 = s13 ? tmp3102 : tmp3271;
  assign tmp3000 = s14 ? tmp3001 : tmp3101;
  assign tmp3332 = s9 ? tmp2380 : tmp2458;
  assign tmp3334 = s8 ? tmp2458 : 1;
  assign tmp3341 = l1 ? tmp2464 : tmp316;
  assign tmp3343 = l1 ? tmp109 : tmp316;
  assign tmp3342 = s0 ? tmp135 : tmp3343;
  assign tmp3340 = s1 ? tmp3341 : tmp3342;
  assign tmp3346 = l1 ? tmp2471 : tmp316;
  assign tmp3345 = s0 ? tmp2469 : tmp3346;
  assign tmp3347 = s1 ? tmp2473 : tmp3346;
  assign tmp3344 = s2 ? tmp3345 : tmp3347;
  assign tmp3339 = s3 ? tmp3340 : tmp3344;
  assign tmp3352 = l1 ? tmp116 : tmp316;
  assign tmp3351 = s0 ? tmp3352 : 1;
  assign tmp3350 = s1 ? tmp3351 : tmp3346;
  assign tmp3354 = s0 ? tmp3341 : 1;
  assign tmp3353 = s1 ? tmp3354 : tmp135;
  assign tmp3349 = s2 ? tmp3350 : tmp3353;
  assign tmp3358 = l1 ? tmp2485 : tmp316;
  assign tmp3357 = s0 ? tmp3346 : tmp3358;
  assign tmp3359 = s0 ? tmp2410 : tmp3346;
  assign tmp3356 = s1 ? tmp3357 : tmp3359;
  assign tmp3355 = s2 ? tmp2404 : tmp3356;
  assign tmp3348 = s3 ? tmp3349 : tmp3355;
  assign tmp3338 = s4 ? tmp3339 : tmp3348;
  assign tmp3365 = s0 ? tmp3343 : 1;
  assign tmp3364 = s1 ? tmp3365 : tmp2493;
  assign tmp3367 = s0 ? tmp3358 : tmp135;
  assign tmp3366 = s1 ? tmp3343 : tmp3367;
  assign tmp3363 = s2 ? tmp3364 : tmp3366;
  assign tmp3369 = s1 ? tmp2499 : tmp2455;
  assign tmp3370 = ~(s1 ? tmp2425 : tmp3357);
  assign tmp3368 = ~(s2 ? tmp3369 : tmp3370);
  assign tmp3362 = s3 ? tmp3363 : tmp3368;
  assign tmp3374 = s0 ? tmp2433 : tmp3346;
  assign tmp3373 = s1 ? tmp3374 : tmp2434;
  assign tmp3372 = s2 ? tmp3373 : tmp3352;
  assign tmp3378 = ~(l1 ? tmp2485 : tmp203);
  assign tmp3377 = s0 ? tmp172 : tmp3378;
  assign tmp3376 = s1 ? tmp3377 : tmp2455;
  assign tmp3375 = ~(s2 ? tmp3376 : tmp2441);
  assign tmp3371 = s3 ? tmp3372 : tmp3375;
  assign tmp3361 = s4 ? tmp3362 : tmp3371;
  assign tmp3383 = s0 ? tmp2410 : tmp31;
  assign tmp3382 = s1 ? tmp3383 : 0;
  assign tmp3381 = s2 ? tmp3382 : tmp244;
  assign tmp3380 = s3 ? tmp3381 : tmp2580;
  assign tmp3386 = l1 ? tmp74 : tmp173;
  assign tmp3385 = s2 ? tmp2454 : tmp3386;
  assign tmp3384 = ~(s3 ? tmp3385 : tmp2586);
  assign tmp3379 = s4 ? tmp3380 : tmp3384;
  assign tmp3360 = s5 ? tmp3361 : tmp3379;
  assign tmp3337 = s6 ? tmp3338 : tmp3360;
  assign tmp3336 = s7 ? tmp2661 : tmp3337;
  assign tmp3335 = ~(s8 ? tmp3336 : tmp2664);
  assign tmp3333 = s9 ? tmp3334 : tmp3335;
  assign tmp3331 = s10 ? tmp3332 : tmp3333;
  assign tmp3330 = s12 ? tmp2167 : tmp3331;
  assign tmp3329 = s13 ? tmp3330 : tmp2666;
  assign tmp3328 = s14 ? tmp1671 : tmp3329;
  assign tmp2999 = s15 ? tmp3000 : tmp3328;
  assign tmp2 = s16 ? tmp3 : tmp2999;
  assign tmp3394 = s8 ? tmp3105 : tmp834;
  assign tmp3393 = s9 ? tmp3105 : tmp3394;
  assign tmp3397 = ~(s7 ? tmp3106 : tmp774);
  assign tmp3396 = ~(s8 ? tmp884 : tmp3397);
  assign tmp3395 = s9 ? tmp882 : tmp3396;
  assign tmp3392 = s10 ? tmp3393 : tmp3395;
  assign tmp3402 = ~(s6 ? tmp1050 : tmp1074);
  assign tmp3401 = s7 ? 1 : tmp3402;
  assign tmp3400 = s8 ? tmp3214 : tmp3401;
  assign tmp3399 = s9 ? tmp3214 : tmp3400;
  assign tmp3404 = s7 ? tmp3215 : tmp968;
  assign tmp3403 = s9 ? tmp1045 : tmp3404;
  assign tmp3398 = s10 ? tmp3399 : tmp3403;
  assign tmp3391 = s12 ? tmp3392 : tmp3398;
  assign tmp3390 = s13 ? tmp3391 : tmp1110;
  assign tmp3389 = s14 ? tmp5 : tmp3390;
  assign tmp3388 = s15 ? tmp3389 : tmp1670;
  assign tmp3387 = s16 ? tmp3388 : tmp2999;
  assign tmp1 = ~(s17 ? tmp2 : tmp3387);
  assign recovery__1 = tmp1;

  assign tmp3420 = l4 ? 1 : 0;
  assign tmp3419 = ~(l3 ? tmp3420 : 1);
  assign tmp3418 = l2 ? 1 : tmp3419;
  assign tmp3422 = l3 ? 1 : 0;
  assign tmp3424 = ~(l4 ? 1 : 0);
  assign tmp3423 = ~(l3 ? 1 : tmp3424);
  assign tmp3421 = ~(l2 ? tmp3422 : tmp3423);
  assign tmp3417 = l1 ? tmp3418 : tmp3421;
  assign tmp3427 = l2 ? tmp3422 : 0;
  assign tmp3426 = l1 ? 1 : tmp3427;
  assign tmp3429 = l2 ? 1 : tmp3424;
  assign tmp3428 = ~(l1 ? tmp3429 : tmp3421);
  assign tmp3425 = ~(s0 ? tmp3426 : tmp3428);
  assign tmp3416 = s1 ? tmp3417 : tmp3425;
  assign tmp3434 = l2 ? 1 : 0;
  assign tmp3436 = ~(l3 ? 1 : 0);
  assign tmp3435 = ~(l2 ? 1 : tmp3436);
  assign tmp3433 = l1 ? tmp3434 : tmp3435;
  assign tmp3438 = l2 ? tmp3420 : tmp3423;
  assign tmp3437 = ~(l1 ? tmp3420 : tmp3438);
  assign tmp3432 = s0 ? tmp3433 : tmp3437;
  assign tmp3441 = ~(l2 ? tmp3422 : tmp3436);
  assign tmp3440 = l1 ? tmp3418 : tmp3441;
  assign tmp3439 = s0 ? tmp3440 : tmp3437;
  assign tmp3431 = s1 ? tmp3432 : tmp3439;
  assign tmp3444 = ~(l1 ? 1 : tmp3434);
  assign tmp3443 = s0 ? tmp3440 : tmp3444;
  assign tmp3446 = l1 ? tmp3420 : tmp3438;
  assign tmp3448 = l2 ? tmp3422 : tmp3423;
  assign tmp3447 = l1 ? tmp3420 : tmp3448;
  assign tmp3445 = ~(s0 ? tmp3446 : tmp3447);
  assign tmp3442 = s1 ? tmp3443 : tmp3445;
  assign tmp3430 = s2 ? tmp3431 : tmp3442;
  assign tmp3415 = s3 ? tmp3416 : tmp3430;
  assign tmp3453 = l1 ? tmp3434 : tmp3421;
  assign tmp3452 = s0 ? tmp3453 : tmp3444;
  assign tmp3454 = ~(s0 ? tmp3447 : tmp3446);
  assign tmp3451 = s1 ? tmp3452 : tmp3454;
  assign tmp3457 = ~(l1 ? 1 : 0);
  assign tmp3456 = s0 ? tmp3417 : tmp3457;
  assign tmp3459 = l1 ? 1 : tmp3422;
  assign tmp3460 = l1 ? 1 : 0;
  assign tmp3458 = ~(s0 ? tmp3459 : tmp3460);
  assign tmp3455 = s1 ? tmp3456 : tmp3458;
  assign tmp3450 = s2 ? tmp3451 : tmp3455;
  assign tmp3463 = s0 ? tmp3459 : tmp3426;
  assign tmp3464 = s0 ? tmp3460 : 0;
  assign tmp3462 = s1 ? tmp3463 : tmp3464;
  assign tmp3466 = ~(s0 ? 1 : tmp3437);
  assign tmp3465 = s1 ? tmp3446 : tmp3466;
  assign tmp3461 = ~(s2 ? tmp3462 : tmp3465);
  assign tmp3449 = s3 ? tmp3450 : tmp3461;
  assign tmp3414 = s4 ? tmp3415 : tmp3449;
  assign tmp3473 = l1 ? tmp3429 : tmp3421;
  assign tmp3472 = s0 ? tmp3473 : tmp3444;
  assign tmp3475 = l1 ? 1 : tmp3434;
  assign tmp3476 = ~(l1 ? tmp3434 : tmp3435);
  assign tmp3474 = ~(s0 ? tmp3475 : tmp3476);
  assign tmp3471 = s1 ? tmp3472 : tmp3474;
  assign tmp3480 = ~(l3 ? 1 : tmp3420);
  assign tmp3479 = ~(l1 ? tmp3429 : tmp3480);
  assign tmp3478 = s0 ? tmp3475 : tmp3479;
  assign tmp3481 = s0 ? tmp3446 : tmp3434;
  assign tmp3477 = ~(s1 ? tmp3478 : tmp3481);
  assign tmp3470 = s2 ? tmp3471 : tmp3477;
  assign tmp3486 = l2 ? 1 : tmp3422;
  assign tmp3485 = ~(l1 ? tmp3486 : tmp3441);
  assign tmp3484 = s0 ? tmp3434 : tmp3485;
  assign tmp3487 = s0 ? tmp3434 : tmp3420;
  assign tmp3483 = s1 ? tmp3484 : tmp3487;
  assign tmp3488 = ~(s1 ? 1 : tmp3424);
  assign tmp3482 = ~(s2 ? tmp3483 : tmp3488);
  assign tmp3469 = s3 ? tmp3470 : tmp3482;
  assign tmp3494 = l2 ? tmp3422 : tmp3420;
  assign tmp3493 = ~(l1 ? tmp3420 : tmp3494);
  assign tmp3492 = s0 ? 1 : tmp3493;
  assign tmp3495 = ~(s0 ? 1 : tmp3460);
  assign tmp3491 = s1 ? tmp3492 : tmp3495;
  assign tmp3497 = s0 ? 1 : tmp3460;
  assign tmp3499 = l1 ? tmp3434 : tmp3480;
  assign tmp3498 = ~(s0 ? tmp3499 : 0);
  assign tmp3496 = ~(s1 ? tmp3497 : tmp3498);
  assign tmp3490 = s2 ? tmp3491 : tmp3496;
  assign tmp3503 = l1 ? tmp3486 : tmp3429;
  assign tmp3502 = s0 ? tmp3499 : tmp3503;
  assign tmp3504 = ~(s0 ? tmp3460 : tmp3420);
  assign tmp3501 = s1 ? tmp3502 : tmp3504;
  assign tmp3500 = s2 ? tmp3501 : 1;
  assign tmp3489 = s3 ? tmp3490 : tmp3500;
  assign tmp3468 = s4 ? tmp3469 : tmp3489;
  assign tmp3509 = s0 ? tmp3420 : 0;
  assign tmp3508 = s1 ? tmp3509 : 0;
  assign tmp3512 = l1 ? tmp3434 : 0;
  assign tmp3511 = s0 ? 1 : tmp3512;
  assign tmp3510 = ~(s1 ? tmp3511 : tmp3512);
  assign tmp3507 = s2 ? tmp3508 : tmp3510;
  assign tmp3515 = s0 ? tmp3512 : 1;
  assign tmp3514 = s1 ? tmp3515 : 1;
  assign tmp3518 = l1 ? tmp3434 : tmp3424;
  assign tmp3517 = s0 ? 1 : tmp3518;
  assign tmp3516 = s1 ? 1 : tmp3517;
  assign tmp3513 = ~(s2 ? tmp3514 : tmp3516);
  assign tmp3506 = s3 ? tmp3507 : tmp3513;
  assign tmp3522 = s0 ? tmp3518 : 1;
  assign tmp3521 = s1 ? tmp3522 : 1;
  assign tmp3525 = l1 ? tmp3429 : tmp3480;
  assign tmp3524 = s0 ? 1 : tmp3525;
  assign tmp3523 = s1 ? tmp3524 : tmp3512;
  assign tmp3520 = s2 ? tmp3521 : tmp3523;
  assign tmp3530 = ~(l2 ? 1 : tmp3424);
  assign tmp3529 = ~(l1 ? tmp3420 : tmp3530);
  assign tmp3528 = s0 ? 1 : tmp3529;
  assign tmp3527 = s1 ? 1 : tmp3528;
  assign tmp3531 = s1 ? tmp3517 : 1;
  assign tmp3526 = s2 ? tmp3527 : tmp3531;
  assign tmp3519 = ~(s3 ? tmp3520 : tmp3526);
  assign tmp3505 = ~(s4 ? tmp3506 : tmp3519);
  assign tmp3467 = s5 ? tmp3468 : tmp3505;
  assign tmp3413 = s6 ? tmp3414 : tmp3467;
  assign tmp3538 = l3 ? tmp3420 : 1;
  assign tmp3537 = l2 ? tmp3420 : tmp3538;
  assign tmp3536 = l1 ? tmp3537 : tmp3448;
  assign tmp3539 = s0 ? tmp3426 : tmp3447;
  assign tmp3535 = s1 ? tmp3536 : tmp3539;
  assign tmp3544 = l2 ? tmp3420 : 1;
  assign tmp3545 = l2 ? tmp3422 : tmp3436;
  assign tmp3543 = l1 ? tmp3544 : tmp3545;
  assign tmp3548 = l3 ? tmp3420 : 0;
  assign tmp3547 = l2 ? tmp3548 : tmp3423;
  assign tmp3546 = l1 ? tmp3420 : tmp3547;
  assign tmp3542 = s0 ? tmp3543 : tmp3546;
  assign tmp3550 = l1 ? tmp3537 : tmp3545;
  assign tmp3549 = s0 ? tmp3550 : tmp3546;
  assign tmp3541 = s1 ? tmp3542 : tmp3549;
  assign tmp3552 = s0 ? tmp3550 : tmp3426;
  assign tmp3553 = s0 ? tmp3546 : tmp3447;
  assign tmp3551 = s1 ? tmp3552 : tmp3553;
  assign tmp3540 = s2 ? tmp3541 : tmp3551;
  assign tmp3534 = s3 ? tmp3535 : tmp3540;
  assign tmp3558 = l1 ? tmp3544 : tmp3448;
  assign tmp3557 = s0 ? tmp3558 : tmp3475;
  assign tmp3559 = s0 ? tmp3447 : tmp3546;
  assign tmp3556 = s1 ? tmp3557 : tmp3559;
  assign tmp3561 = s0 ? tmp3536 : tmp3460;
  assign tmp3562 = s0 ? tmp3459 : tmp3460;
  assign tmp3560 = s1 ? tmp3561 : tmp3562;
  assign tmp3555 = s2 ? tmp3556 : tmp3560;
  assign tmp3566 = ~(l1 ? tmp3420 : tmp3547);
  assign tmp3565 = ~(s0 ? 1 : tmp3566);
  assign tmp3564 = s1 ? tmp3546 : tmp3565;
  assign tmp3563 = s2 ? tmp3462 : tmp3564;
  assign tmp3554 = s3 ? tmp3555 : tmp3563;
  assign tmp3533 = s4 ? tmp3534 : tmp3554;
  assign tmp3572 = s0 ? tmp3447 : tmp3475;
  assign tmp3573 = s0 ? tmp3475 : tmp3543;
  assign tmp3571 = s1 ? tmp3572 : tmp3573;
  assign tmp3576 = l1 ? tmp3420 : tmp3494;
  assign tmp3575 = s0 ? tmp3475 : tmp3576;
  assign tmp3577 = s0 ? tmp3546 : tmp3426;
  assign tmp3574 = s1 ? tmp3575 : tmp3577;
  assign tmp3570 = s2 ? tmp3571 : tmp3574;
  assign tmp3582 = l2 ? tmp3420 : tmp3436;
  assign tmp3581 = l1 ? tmp3582 : tmp3545;
  assign tmp3580 = s0 ? tmp3426 : tmp3581;
  assign tmp3585 = l2 ? tmp3548 : tmp3420;
  assign tmp3584 = l1 ? tmp3420 : tmp3585;
  assign tmp3583 = s0 ? tmp3426 : tmp3584;
  assign tmp3579 = s1 ? tmp3580 : tmp3583;
  assign tmp3587 = ~(l1 ? tmp3420 : tmp3585);
  assign tmp3586 = ~(s1 ? 1 : tmp3587);
  assign tmp3578 = s2 ? tmp3579 : tmp3586;
  assign tmp3569 = s3 ? tmp3570 : tmp3578;
  assign tmp3592 = l1 ? tmp3544 : tmp3494;
  assign tmp3591 = s0 ? tmp3592 : 1;
  assign tmp3590 = ~(s1 ? tmp3497 : tmp3591);
  assign tmp3589 = s2 ? tmp3491 : tmp3590;
  assign tmp3597 = ~(l2 ? tmp3422 : tmp3420);
  assign tmp3596 = l1 ? tmp3434 : tmp3597;
  assign tmp3598 = ~(l1 ? tmp3582 : tmp3530);
  assign tmp3595 = s0 ? tmp3596 : tmp3598;
  assign tmp3594 = s1 ? tmp3595 : tmp3504;
  assign tmp3593 = s2 ? tmp3594 : 1;
  assign tmp3588 = ~(s3 ? tmp3589 : tmp3593);
  assign tmp3568 = s4 ? tmp3569 : tmp3588;
  assign tmp3603 = s0 ? tmp3584 : 0;
  assign tmp3602 = s1 ? tmp3603 : 0;
  assign tmp3607 = ~(l2 ? tmp3422 : 1);
  assign tmp3606 = l1 ? tmp3434 : tmp3607;
  assign tmp3605 = s0 ? 1 : tmp3606;
  assign tmp3608 = s0 ? tmp3512 : tmp3606;
  assign tmp3604 = ~(s1 ? tmp3605 : tmp3608);
  assign tmp3601 = s2 ? tmp3602 : tmp3604;
  assign tmp3600 = s3 ? tmp3601 : tmp3513;
  assign tmp3613 = l1 ? tmp3429 : tmp3597;
  assign tmp3612 = s0 ? 1 : tmp3613;
  assign tmp3614 = s0 ? tmp3606 : tmp3512;
  assign tmp3611 = s1 ? tmp3612 : tmp3614;
  assign tmp3610 = s2 ? tmp3521 : tmp3611;
  assign tmp3609 = ~(s3 ? tmp3610 : tmp3526);
  assign tmp3599 = s4 ? tmp3600 : tmp3609;
  assign tmp3567 = s5 ? tmp3568 : tmp3599;
  assign tmp3532 = ~(s6 ? tmp3533 : tmp3567);
  assign tmp3412 = s8 ? tmp3413 : tmp3532;
  assign tmp3616 = s6 ? tmp3533 : tmp3567;
  assign tmp3622 = ~(l2 ? tmp3422 : 0);
  assign tmp3621 = l1 ? tmp3418 : tmp3622;
  assign tmp3624 = l1 ? tmp3434 : tmp3622;
  assign tmp3625 = l1 ? tmp3429 : tmp3622;
  assign tmp3623 = s0 ? tmp3624 : tmp3625;
  assign tmp3620 = s1 ? tmp3621 : tmp3623;
  assign tmp3630 = ~(l2 ? tmp3548 : 0);
  assign tmp3629 = l1 ? tmp3429 : tmp3630;
  assign tmp3628 = s0 ? tmp3624 : tmp3629;
  assign tmp3631 = s0 ? tmp3621 : tmp3629;
  assign tmp3627 = s1 ? tmp3628 : tmp3631;
  assign tmp3633 = s0 ? tmp3621 : tmp3624;
  assign tmp3634 = s0 ? tmp3629 : tmp3625;
  assign tmp3632 = s1 ? tmp3633 : tmp3634;
  assign tmp3626 = s2 ? tmp3627 : tmp3632;
  assign tmp3619 = s3 ? tmp3620 : tmp3626;
  assign tmp3640 = ~(l2 ? 1 : 0);
  assign tmp3639 = l1 ? tmp3434 : tmp3640;
  assign tmp3638 = s0 ? tmp3624 : tmp3639;
  assign tmp3641 = s0 ? tmp3625 : tmp3629;
  assign tmp3637 = s1 ? tmp3638 : tmp3641;
  assign tmp3644 = l1 ? tmp3434 : 1;
  assign tmp3643 = s0 ? tmp3621 : tmp3644;
  assign tmp3646 = l1 ? tmp3434 : tmp3436;
  assign tmp3645 = s0 ? tmp3646 : tmp3644;
  assign tmp3642 = s1 ? tmp3643 : tmp3645;
  assign tmp3636 = s2 ? tmp3637 : tmp3642;
  assign tmp3649 = s0 ? tmp3646 : tmp3624;
  assign tmp3650 = s0 ? tmp3644 : 1;
  assign tmp3648 = s1 ? tmp3649 : tmp3650;
  assign tmp3652 = s0 ? 1 : tmp3629;
  assign tmp3651 = s1 ? tmp3629 : tmp3652;
  assign tmp3647 = s2 ? tmp3648 : tmp3651;
  assign tmp3635 = s3 ? tmp3636 : tmp3647;
  assign tmp3618 = s4 ? tmp3619 : tmp3635;
  assign tmp3658 = s0 ? tmp3625 : tmp3444;
  assign tmp3660 = ~(l1 ? tmp3434 : tmp3622);
  assign tmp3659 = ~(s0 ? tmp3475 : tmp3660);
  assign tmp3657 = s1 ? tmp3658 : tmp3659;
  assign tmp3663 = ~(l1 ? tmp3429 : tmp3622);
  assign tmp3662 = s0 ? tmp3475 : tmp3663;
  assign tmp3665 = l1 ? 1 : tmp3622;
  assign tmp3664 = ~(s0 ? tmp3629 : tmp3665);
  assign tmp3661 = ~(s1 ? tmp3662 : tmp3664);
  assign tmp3656 = s2 ? tmp3657 : tmp3661;
  assign tmp3669 = l1 ? tmp3486 : tmp3622;
  assign tmp3668 = s0 ? tmp3665 : tmp3669;
  assign tmp3672 = l2 ? tmp3548 : 0;
  assign tmp3671 = ~(l1 ? tmp3420 : tmp3672);
  assign tmp3670 = s0 ? tmp3665 : tmp3671;
  assign tmp3667 = s1 ? tmp3668 : tmp3670;
  assign tmp3674 = ~(l2 ? tmp3548 : tmp3420);
  assign tmp3673 = s1 ? 1 : tmp3674;
  assign tmp3666 = s2 ? tmp3667 : tmp3673;
  assign tmp3655 = s3 ? tmp3656 : tmp3666;
  assign tmp3678 = s0 ? 1 : tmp3625;
  assign tmp3679 = s0 ? tmp3512 : tmp3644;
  assign tmp3677 = s1 ? tmp3678 : tmp3679;
  assign tmp3681 = s0 ? tmp3624 : tmp3512;
  assign tmp3680 = s1 ? tmp3679 : tmp3681;
  assign tmp3676 = s2 ? tmp3677 : tmp3680;
  assign tmp3685 = l1 ? tmp3486 : 1;
  assign tmp3684 = s0 ? tmp3624 : tmp3685;
  assign tmp3686 = s0 ? tmp3644 : tmp3424;
  assign tmp3683 = s1 ? tmp3684 : tmp3686;
  assign tmp3682 = s2 ? tmp3683 : 1;
  assign tmp3675 = s3 ? tmp3676 : tmp3682;
  assign tmp3654 = s4 ? tmp3655 : tmp3675;
  assign tmp3692 = l1 ? tmp3420 : tmp3672;
  assign tmp3691 = s0 ? tmp3692 : 0;
  assign tmp3690 = s1 ? tmp3691 : 0;
  assign tmp3694 = s0 ? 1 : tmp3646;
  assign tmp3695 = s0 ? tmp3434 : tmp3646;
  assign tmp3693 = ~(s1 ? tmp3694 : tmp3695);
  assign tmp3689 = s2 ? tmp3690 : tmp3693;
  assign tmp3698 = s0 ? tmp3434 : 1;
  assign tmp3697 = s1 ? tmp3698 : 1;
  assign tmp3700 = s0 ? 1 : tmp3644;
  assign tmp3699 = s1 ? 1 : tmp3700;
  assign tmp3696 = ~(s2 ? tmp3697 : tmp3699);
  assign tmp3688 = s3 ? tmp3689 : tmp3696;
  assign tmp3703 = s1 ? tmp3650 : 1;
  assign tmp3705 = s0 ? tmp3646 : tmp3434;
  assign tmp3704 = s1 ? tmp3678 : tmp3705;
  assign tmp3702 = s2 ? tmp3703 : tmp3704;
  assign tmp3709 = ~(l1 ? tmp3420 : 0);
  assign tmp3708 = s0 ? 1 : tmp3709;
  assign tmp3707 = s1 ? 1 : tmp3708;
  assign tmp3710 = s1 ? tmp3700 : 1;
  assign tmp3706 = s2 ? tmp3707 : tmp3710;
  assign tmp3701 = ~(s3 ? tmp3702 : tmp3706);
  assign tmp3687 = ~(s4 ? tmp3688 : tmp3701);
  assign tmp3653 = s5 ? tmp3654 : tmp3687;
  assign tmp3617 = ~(s6 ? tmp3618 : tmp3653);
  assign tmp3615 = ~(s8 ? tmp3616 : tmp3617);
  assign tmp3411 = s9 ? tmp3412 : tmp3615;
  assign tmp3715 = s0 ? tmp3624 : tmp3473;
  assign tmp3714 = s1 ? tmp3417 : tmp3715;
  assign tmp3719 = l1 ? tmp3434 : tmp3441;
  assign tmp3721 = ~(l2 ? tmp3548 : tmp3423);
  assign tmp3720 = l1 ? tmp3429 : tmp3721;
  assign tmp3718 = s0 ? tmp3719 : tmp3720;
  assign tmp3722 = s0 ? tmp3440 : tmp3720;
  assign tmp3717 = s1 ? tmp3718 : tmp3722;
  assign tmp3724 = s0 ? tmp3440 : tmp3624;
  assign tmp3725 = s0 ? tmp3720 : tmp3473;
  assign tmp3723 = s1 ? tmp3724 : tmp3725;
  assign tmp3716 = s2 ? tmp3717 : tmp3723;
  assign tmp3713 = s3 ? tmp3714 : tmp3716;
  assign tmp3729 = s0 ? tmp3453 : tmp3639;
  assign tmp3730 = s0 ? tmp3473 : tmp3720;
  assign tmp3728 = s1 ? tmp3729 : tmp3730;
  assign tmp3732 = s0 ? tmp3417 : tmp3644;
  assign tmp3731 = s1 ? tmp3732 : tmp3645;
  assign tmp3727 = s2 ? tmp3728 : tmp3731;
  assign tmp3735 = s0 ? 1 : tmp3720;
  assign tmp3734 = s1 ? tmp3720 : tmp3735;
  assign tmp3733 = s2 ? tmp3648 : tmp3734;
  assign tmp3726 = s3 ? tmp3727 : tmp3733;
  assign tmp3712 = s4 ? tmp3713 : tmp3726;
  assign tmp3742 = ~(l1 ? tmp3434 : tmp3441);
  assign tmp3741 = ~(s0 ? tmp3475 : tmp3742);
  assign tmp3740 = s1 ? tmp3472 : tmp3741;
  assign tmp3745 = ~(l1 ? tmp3429 : tmp3597);
  assign tmp3744 = s0 ? tmp3475 : tmp3745;
  assign tmp3746 = ~(s0 ? tmp3720 : tmp3665);
  assign tmp3743 = ~(s1 ? tmp3744 : tmp3746);
  assign tmp3739 = s2 ? tmp3740 : tmp3743;
  assign tmp3750 = l1 ? tmp3486 : tmp3441;
  assign tmp3749 = s0 ? tmp3665 : tmp3750;
  assign tmp3751 = s0 ? tmp3665 : tmp3587;
  assign tmp3748 = s1 ? tmp3749 : tmp3751;
  assign tmp3747 = s2 ? tmp3748 : tmp3673;
  assign tmp3738 = s3 ? tmp3739 : tmp3747;
  assign tmp3754 = s1 ? tmp3612 : tmp3679;
  assign tmp3756 = s0 ? tmp3596 : tmp3512;
  assign tmp3755 = s1 ? tmp3679 : tmp3756;
  assign tmp3753 = s2 ? tmp3754 : tmp3755;
  assign tmp3759 = s0 ? tmp3596 : tmp3503;
  assign tmp3758 = s1 ? tmp3759 : tmp3686;
  assign tmp3757 = s2 ? tmp3758 : 1;
  assign tmp3752 = s3 ? tmp3753 : tmp3757;
  assign tmp3737 = s4 ? tmp3738 : tmp3752;
  assign tmp3760 = ~(s4 ? tmp3600 : tmp3609);
  assign tmp3736 = s5 ? tmp3737 : tmp3760;
  assign tmp3711 = s6 ? tmp3712 : tmp3736;
  assign tmp3410 = s10 ? tmp3411 : tmp3711;
  assign tmp3771 = ~(l3 ? tmp3420 : 0);
  assign tmp3770 = l2 ? 1 : tmp3771;
  assign tmp3772 = ~(l2 ? tmp3422 : tmp3548);
  assign tmp3769 = l1 ? tmp3770 : tmp3772;
  assign tmp3775 = l2 ? tmp3422 : 1;
  assign tmp3774 = l1 ? tmp3422 : tmp3775;
  assign tmp3776 = ~(l1 ? tmp3770 : tmp3436);
  assign tmp3773 = ~(s0 ? tmp3774 : tmp3776);
  assign tmp3768 = s1 ? tmp3769 : tmp3773;
  assign tmp3781 = l2 ? 1 : tmp3436;
  assign tmp3782 = ~(l2 ? 1 : tmp3422);
  assign tmp3780 = l1 ? tmp3781 : tmp3782;
  assign tmp3783 = ~(l2 ? tmp3420 : tmp3548);
  assign tmp3779 = s0 ? tmp3780 : tmp3783;
  assign tmp3785 = l1 ? tmp3770 : tmp3436;
  assign tmp3784 = s0 ? tmp3785 : tmp3783;
  assign tmp3778 = s1 ? tmp3779 : tmp3784;
  assign tmp3787 = s0 ? tmp3785 : 0;
  assign tmp3789 = l2 ? tmp3420 : tmp3548;
  assign tmp3790 = ~(l1 ? tmp3770 : tmp3772);
  assign tmp3788 = ~(s0 ? tmp3789 : tmp3790);
  assign tmp3786 = s1 ? tmp3787 : tmp3788;
  assign tmp3777 = s2 ? tmp3778 : tmp3786;
  assign tmp3767 = s3 ? tmp3768 : tmp3777;
  assign tmp3795 = l1 ? tmp3781 : tmp3436;
  assign tmp3796 = ~(l1 ? tmp3422 : 1);
  assign tmp3794 = s0 ? tmp3795 : tmp3796;
  assign tmp3797 = s0 ? tmp3769 : tmp3783;
  assign tmp3793 = s1 ? tmp3794 : tmp3797;
  assign tmp3799 = s0 ? tmp3769 : 0;
  assign tmp3800 = ~(s0 ? tmp3422 : 1);
  assign tmp3798 = s1 ? tmp3799 : tmp3800;
  assign tmp3792 = s2 ? tmp3793 : tmp3798;
  assign tmp3803 = s0 ? 1 : 0;
  assign tmp3802 = s1 ? tmp3774 : tmp3803;
  assign tmp3805 = ~(s0 ? 1 : tmp3783);
  assign tmp3804 = s1 ? tmp3789 : tmp3805;
  assign tmp3801 = ~(s2 ? tmp3802 : tmp3804);
  assign tmp3791 = s3 ? tmp3792 : tmp3801;
  assign tmp3766 = s4 ? tmp3767 : tmp3791;
  assign tmp3812 = ~(l1 ? tmp3781 : tmp3782);
  assign tmp3811 = ~(s0 ? 1 : tmp3812);
  assign tmp3810 = s1 ? tmp3787 : tmp3811;
  assign tmp3815 = ~(l1 ? tmp3770 : tmp3622);
  assign tmp3814 = s0 ? 1 : tmp3815;
  assign tmp3816 = s0 ? tmp3789 : 1;
  assign tmp3813 = ~(s1 ? tmp3814 : tmp3816);
  assign tmp3809 = s2 ? tmp3810 : tmp3813;
  assign tmp3820 = ~(l1 ? 1 : tmp3436);
  assign tmp3819 = s0 ? 1 : tmp3820;
  assign tmp3822 = l2 ? tmp3420 : 0;
  assign tmp3821 = s0 ? 1 : tmp3822;
  assign tmp3818 = s1 ? tmp3819 : tmp3821;
  assign tmp3823 = ~(s1 ? 1 : tmp3783);
  assign tmp3817 = ~(s2 ? tmp3818 : tmp3823);
  assign tmp3808 = s3 ? tmp3809 : tmp3817;
  assign tmp3828 = l1 ? tmp3770 : tmp3622;
  assign tmp3827 = s0 ? 1 : tmp3828;
  assign tmp3830 = l1 ? tmp3422 : 1;
  assign tmp3829 = ~(s0 ? tmp3830 : 0);
  assign tmp3826 = s1 ? tmp3827 : tmp3829;
  assign tmp3832 = s0 ? tmp3830 : 0;
  assign tmp3834 = l1 ? tmp3781 : tmp3622;
  assign tmp3833 = ~(s0 ? tmp3834 : tmp3796);
  assign tmp3831 = ~(s1 ? tmp3832 : tmp3833);
  assign tmp3825 = s2 ? tmp3826 : tmp3831;
  assign tmp3837 = s0 ? tmp3665 : 1;
  assign tmp3836 = s1 ? tmp3837 : 1;
  assign tmp3835 = s2 ? tmp3836 : 1;
  assign tmp3824 = s3 ? tmp3825 : tmp3835;
  assign tmp3807 = s4 ? tmp3808 : tmp3824;
  assign tmp3842 = s0 ? tmp3822 : 0;
  assign tmp3841 = s1 ? tmp3842 : 0;
  assign tmp3845 = l1 ? 1 : tmp3640;
  assign tmp3844 = s0 ? 1 : tmp3845;
  assign tmp3843 = ~(s1 ? tmp3844 : tmp3845);
  assign tmp3840 = s2 ? tmp3841 : tmp3843;
  assign tmp3839 = s3 ? tmp3840 : 0;
  assign tmp3849 = s0 ? 1 : tmp3665;
  assign tmp3848 = s1 ? tmp3849 : tmp3845;
  assign tmp3847 = s2 ? 1 : tmp3848;
  assign tmp3846 = ~(s3 ? tmp3847 : 1);
  assign tmp3838 = ~(s4 ? tmp3839 : tmp3846);
  assign tmp3806 = s5 ? tmp3807 : tmp3838;
  assign tmp3765 = s6 ? tmp3766 : tmp3806;
  assign tmp3855 = l2 ? tmp3422 : tmp3548;
  assign tmp3854 = l1 ? tmp3789 : tmp3855;
  assign tmp3857 = l1 ? tmp3486 : tmp3775;
  assign tmp3858 = l1 ? tmp3789 : tmp3422;
  assign tmp3856 = s0 ? tmp3857 : tmp3858;
  assign tmp3853 = s1 ? tmp3854 : tmp3856;
  assign tmp3863 = l2 ? tmp3420 : tmp3422;
  assign tmp3862 = l1 ? tmp3863 : tmp3422;
  assign tmp3864 = l1 ? tmp3789 : tmp3548;
  assign tmp3861 = s0 ? tmp3862 : tmp3864;
  assign tmp3865 = s0 ? tmp3858 : tmp3864;
  assign tmp3860 = s1 ? tmp3861 : tmp3865;
  assign tmp3868 = l1 ? 1 : tmp3775;
  assign tmp3867 = s0 ? tmp3858 : tmp3868;
  assign tmp3869 = s0 ? tmp3864 : tmp3854;
  assign tmp3866 = s1 ? tmp3867 : tmp3869;
  assign tmp3859 = s2 ? tmp3860 : tmp3866;
  assign tmp3852 = s3 ? tmp3853 : tmp3859;
  assign tmp3873 = s0 ? tmp3862 : tmp3685;
  assign tmp3874 = s0 ? tmp3854 : tmp3864;
  assign tmp3872 = s1 ? tmp3873 : tmp3874;
  assign tmp3876 = s0 ? tmp3854 : 1;
  assign tmp3878 = l1 ? tmp3486 : tmp3422;
  assign tmp3877 = s0 ? tmp3878 : 1;
  assign tmp3875 = s1 ? tmp3876 : tmp3877;
  assign tmp3871 = s2 ? tmp3872 : tmp3875;
  assign tmp3880 = s1 ? tmp3857 : tmp3803;
  assign tmp3883 = ~(l1 ? tmp3789 : tmp3548);
  assign tmp3882 = ~(s0 ? 1 : tmp3883);
  assign tmp3881 = s1 ? tmp3864 : tmp3882;
  assign tmp3879 = s2 ? tmp3880 : tmp3881;
  assign tmp3870 = s3 ? tmp3871 : tmp3879;
  assign tmp3851 = s4 ? tmp3852 : tmp3870;
  assign tmp3889 = s0 ? tmp3858 : 1;
  assign tmp3890 = s0 ? 1 : tmp3862;
  assign tmp3888 = s1 ? tmp3889 : tmp3890;
  assign tmp3892 = s0 ? 1 : tmp3858;
  assign tmp3894 = l1 ? tmp3822 : tmp3548;
  assign tmp3893 = s0 ? tmp3894 : tmp3868;
  assign tmp3891 = s1 ? tmp3892 : tmp3893;
  assign tmp3887 = s2 ? tmp3888 : tmp3891;
  assign tmp3898 = l1 ? tmp3822 : tmp3422;
  assign tmp3897 = s0 ? tmp3868 : tmp3898;
  assign tmp3900 = ~(l1 ? 1 : tmp3771);
  assign tmp3899 = s0 ? tmp3868 : tmp3900;
  assign tmp3896 = s1 ? tmp3897 : tmp3899;
  assign tmp3901 = ~(s1 ? 1 : tmp3883);
  assign tmp3895 = s2 ? tmp3896 : tmp3901;
  assign tmp3886 = s3 ? tmp3887 : tmp3895;
  assign tmp3906 = ~(l1 ? tmp3789 : tmp3427);
  assign tmp3905 = s0 ? 1 : tmp3906;
  assign tmp3907 = ~(s0 ? tmp3685 : tmp3512);
  assign tmp3904 = s1 ? tmp3905 : tmp3907;
  assign tmp3909 = s0 ? tmp3685 : tmp3512;
  assign tmp3908 = ~(s1 ? tmp3909 : tmp3873);
  assign tmp3903 = s2 ? tmp3904 : tmp3908;
  assign tmp3913 = l1 ? 1 : tmp3436;
  assign tmp3914 = ~(l1 ? tmp3822 : 0);
  assign tmp3912 = s0 ? tmp3913 : tmp3914;
  assign tmp3915 = ~(s0 ? tmp3512 : 0);
  assign tmp3911 = s1 ? tmp3912 : tmp3915;
  assign tmp3910 = s2 ? tmp3911 : 1;
  assign tmp3902 = ~(s3 ? tmp3903 : tmp3910);
  assign tmp3885 = s4 ? tmp3886 : tmp3902;
  assign tmp3921 = l1 ? 1 : tmp3771;
  assign tmp3920 = s0 ? tmp3921 : 1;
  assign tmp3919 = s1 ? tmp3920 : 1;
  assign tmp3922 = s0 ? 1 : tmp3913;
  assign tmp3918 = s2 ? tmp3919 : tmp3922;
  assign tmp3917 = s3 ? tmp3918 : 1;
  assign tmp3926 = s0 ? tmp3913 : 1;
  assign tmp3925 = s1 ? tmp3922 : tmp3926;
  assign tmp3924 = s2 ? 1 : tmp3925;
  assign tmp3923 = s3 ? tmp3924 : 1;
  assign tmp3916 = ~(s4 ? tmp3917 : tmp3923);
  assign tmp3884 = s5 ? tmp3885 : tmp3916;
  assign tmp3850 = ~(s6 ? tmp3851 : tmp3884);
  assign tmp3764 = s8 ? tmp3765 : tmp3850;
  assign tmp3928 = s6 ? tmp3851 : tmp3884;
  assign tmp3933 = l1 ? tmp3770 : tmp3597;
  assign tmp3932 = s1 ? tmp3933 : tmp3773;
  assign tmp3937 = l1 ? tmp3781 : tmp3607;
  assign tmp3938 = ~(l1 ? tmp3548 : tmp3585);
  assign tmp3936 = s0 ? tmp3937 : tmp3938;
  assign tmp3940 = l1 ? tmp3770 : tmp3607;
  assign tmp3939 = s0 ? tmp3940 : tmp3938;
  assign tmp3935 = s1 ? tmp3936 : tmp3939;
  assign tmp3942 = s0 ? tmp3940 : tmp3607;
  assign tmp3944 = l1 ? tmp3548 : tmp3585;
  assign tmp3945 = l1 ? tmp3548 : tmp3494;
  assign tmp3943 = ~(s0 ? tmp3944 : tmp3945);
  assign tmp3941 = s1 ? tmp3942 : tmp3943;
  assign tmp3934 = s2 ? tmp3935 : tmp3941;
  assign tmp3931 = s3 ? tmp3932 : tmp3934;
  assign tmp3949 = ~(s0 ? tmp3945 : tmp3944);
  assign tmp3948 = s1 ? tmp3794 : tmp3949;
  assign tmp3951 = s0 ? tmp3933 : tmp3512;
  assign tmp3953 = ~(l1 ? tmp3434 : 0);
  assign tmp3952 = ~(s0 ? tmp3422 : tmp3953);
  assign tmp3950 = s1 ? tmp3951 : tmp3952;
  assign tmp3947 = s2 ? tmp3948 : tmp3950;
  assign tmp3956 = ~(s0 ? tmp3512 : 1);
  assign tmp3955 = s1 ? tmp3774 : tmp3956;
  assign tmp3958 = ~(s0 ? 1 : tmp3938);
  assign tmp3957 = s1 ? tmp3944 : tmp3958;
  assign tmp3954 = ~(s2 ? tmp3955 : tmp3957);
  assign tmp3946 = s3 ? tmp3947 : tmp3954;
  assign tmp3930 = s4 ? tmp3931 : tmp3946;
  assign tmp3965 = ~(l1 ? tmp3781 : tmp3607);
  assign tmp3964 = ~(s0 ? 1 : tmp3965);
  assign tmp3963 = s1 ? tmp3787 : tmp3964;
  assign tmp3968 = l1 ? 1 : tmp3674;
  assign tmp3967 = ~(s0 ? tmp3968 : tmp3607);
  assign tmp3966 = ~(s1 ? tmp3814 : tmp3967);
  assign tmp3962 = s2 ? tmp3963 : tmp3966;
  assign tmp3972 = ~(l1 ? 1 : tmp3607);
  assign tmp3971 = s0 ? tmp3775 : tmp3972;
  assign tmp3974 = ~(l1 ? 1 : tmp3630);
  assign tmp3973 = s0 ? tmp3775 : tmp3974;
  assign tmp3970 = s1 ? tmp3971 : tmp3973;
  assign tmp3976 = ~(l1 ? tmp3548 : tmp3672);
  assign tmp3975 = ~(s1 ? 1 : tmp3976);
  assign tmp3969 = ~(s2 ? tmp3970 : tmp3975);
  assign tmp3961 = s3 ? tmp3962 : tmp3969;
  assign tmp3981 = ~(l1 ? tmp3548 : tmp3427);
  assign tmp3980 = s0 ? 1 : tmp3981;
  assign tmp3979 = s1 ? tmp3980 : tmp3829;
  assign tmp3978 = s2 ? tmp3979 : tmp3831;
  assign tmp3977 = s3 ? tmp3978 : tmp3835;
  assign tmp3960 = s4 ? tmp3961 : tmp3977;
  assign tmp3987 = l1 ? 1 : tmp3630;
  assign tmp3986 = s0 ? tmp3987 : 1;
  assign tmp3985 = s1 ? tmp3986 : 1;
  assign tmp3984 = s2 ? tmp3985 : tmp3922;
  assign tmp3983 = s3 ? tmp3984 : 1;
  assign tmp3990 = s1 ? tmp3849 : tmp3926;
  assign tmp3989 = s2 ? 1 : tmp3990;
  assign tmp3988 = s3 ? tmp3989 : 1;
  assign tmp3982 = s4 ? tmp3983 : tmp3988;
  assign tmp3959 = s5 ? tmp3960 : tmp3982;
  assign tmp3929 = ~(s6 ? tmp3930 : tmp3959);
  assign tmp3927 = ~(s8 ? tmp3928 : tmp3929);
  assign tmp3763 = s9 ? tmp3764 : tmp3927;
  assign tmp3996 = s0 ? tmp3795 : tmp3771;
  assign tmp3997 = s0 ? tmp3785 : tmp3771;
  assign tmp3995 = s1 ? tmp3996 : tmp3997;
  assign tmp3999 = s0 ? tmp3785 : tmp3607;
  assign tmp4001 = l1 ? tmp3548 : tmp3855;
  assign tmp4000 = ~(s0 ? tmp3548 : tmp4001);
  assign tmp3998 = s1 ? tmp3999 : tmp4000;
  assign tmp3994 = s2 ? tmp3995 : tmp3998;
  assign tmp3993 = s3 ? tmp3768 : tmp3994;
  assign tmp4005 = ~(s0 ? tmp4001 : tmp3548);
  assign tmp4004 = s1 ? tmp3794 : tmp4005;
  assign tmp4007 = s0 ? tmp3769 : tmp3512;
  assign tmp4006 = s1 ? tmp4007 : tmp3952;
  assign tmp4003 = s2 ? tmp4004 : tmp4006;
  assign tmp4010 = ~(s0 ? 1 : tmp3771);
  assign tmp4009 = s1 ? tmp3548 : tmp4010;
  assign tmp4008 = ~(s2 ? tmp3955 : tmp4009);
  assign tmp4002 = s3 ? tmp4003 : tmp4008;
  assign tmp3992 = s4 ? tmp3993 : tmp4002;
  assign tmp4017 = ~(l1 ? tmp3781 : tmp3436);
  assign tmp4016 = ~(s0 ? 1 : tmp4017);
  assign tmp4015 = s1 ? tmp3787 : tmp4016;
  assign tmp4019 = s0 ? 1 : tmp3776;
  assign tmp4020 = s0 ? tmp3548 : tmp3775;
  assign tmp4018 = ~(s1 ? tmp4019 : tmp4020);
  assign tmp4014 = s2 ? tmp4015 : tmp4018;
  assign tmp4023 = s0 ? tmp3775 : tmp3820;
  assign tmp4024 = s0 ? tmp3775 : tmp3900;
  assign tmp4022 = s1 ? tmp4023 : tmp4024;
  assign tmp4025 = ~(s1 ? 1 : tmp3771);
  assign tmp4021 = ~(s2 ? tmp4022 : tmp4025);
  assign tmp4013 = s3 ? tmp4014 : tmp4021;
  assign tmp4029 = ~(s0 ? tmp3795 : tmp3796);
  assign tmp4028 = ~(s1 ? tmp3832 : tmp4029);
  assign tmp4027 = s2 ? tmp3979 : tmp4028;
  assign tmp4031 = s1 ? tmp3926 : 1;
  assign tmp4030 = s2 ? tmp4031 : 1;
  assign tmp4026 = s3 ? tmp4027 : tmp4030;
  assign tmp4012 = s4 ? tmp4013 : tmp4026;
  assign tmp4032 = s4 ? tmp3917 : tmp3923;
  assign tmp4011 = s5 ? tmp4012 : tmp4032;
  assign tmp3991 = s6 ? tmp3992 : tmp4011;
  assign tmp3762 = s10 ? tmp3763 : tmp3991;
  assign tmp4041 = l1 ? tmp3422 : tmp3640;
  assign tmp4042 = ~(l1 ? tmp3770 : tmp3781);
  assign tmp4040 = ~(s0 ? tmp4041 : tmp4042);
  assign tmp4039 = s1 ? tmp3770 : tmp4040;
  assign tmp4045 = s0 ? tmp3781 : tmp3770;
  assign tmp4047 = l1 ? tmp3770 : tmp3781;
  assign tmp4046 = s0 ? tmp4047 : tmp3770;
  assign tmp4044 = s1 ? tmp4045 : tmp4046;
  assign tmp4050 = ~(l1 ? 1 : tmp3640);
  assign tmp4049 = s0 ? tmp4047 : tmp4050;
  assign tmp4048 = s1 ? tmp4049 : tmp3770;
  assign tmp4043 = s2 ? tmp4044 : tmp4048;
  assign tmp4038 = s3 ? tmp4039 : tmp4043;
  assign tmp4055 = ~(l1 ? tmp3422 : tmp3640);
  assign tmp4054 = s0 ? tmp3781 : tmp4055;
  assign tmp4053 = s1 ? tmp4054 : tmp3770;
  assign tmp4057 = s0 ? tmp3770 : 0;
  assign tmp4059 = l1 ? tmp3422 : 0;
  assign tmp4058 = ~(s0 ? tmp4059 : 1);
  assign tmp4056 = s1 ? tmp4057 : tmp4058;
  assign tmp4052 = s2 ? tmp4053 : tmp4056;
  assign tmp4061 = s1 ? tmp4041 : tmp3803;
  assign tmp4063 = s0 ? 1 : tmp3770;
  assign tmp4062 = ~(s1 ? tmp3770 : tmp4063);
  assign tmp4060 = ~(s2 ? tmp4061 : tmp4062);
  assign tmp4051 = s3 ? tmp4052 : tmp4060;
  assign tmp4037 = s4 ? tmp4038 : tmp4051;
  assign tmp4069 = ~(s0 ? tmp3845 : tmp3435);
  assign tmp4068 = s1 ? tmp4049 : tmp4069;
  assign tmp4072 = ~(l1 ? tmp3770 : 1);
  assign tmp4071 = s0 ? tmp3845 : tmp4072;
  assign tmp4074 = l1 ? 1 : tmp3770;
  assign tmp4073 = ~(s0 ? tmp4074 : tmp3434);
  assign tmp4070 = ~(s1 ? tmp4071 : tmp4073);
  assign tmp4067 = s2 ? tmp4068 : tmp4070;
  assign tmp4078 = l1 ? 1 : tmp3781;
  assign tmp4077 = s0 ? tmp3434 : tmp4078;
  assign tmp4076 = s1 ? tmp4077 : tmp3698;
  assign tmp4081 = l1 ? tmp3770 : 1;
  assign tmp4080 = s0 ? tmp4081 : 1;
  assign tmp4079 = s1 ? 1 : tmp4080;
  assign tmp4075 = s2 ? tmp4076 : tmp4079;
  assign tmp4066 = s3 ? tmp4067 : tmp4075;
  assign tmp4085 = s0 ? 1 : tmp4081;
  assign tmp4086 = ~(s0 ? tmp4059 : 0);
  assign tmp4084 = s1 ? tmp4085 : tmp4086;
  assign tmp4088 = s0 ? tmp4059 : 0;
  assign tmp4090 = l1 ? tmp3781 : 1;
  assign tmp4091 = ~(l1 ? tmp3422 : 0);
  assign tmp4089 = ~(s0 ? tmp4090 : tmp4091);
  assign tmp4087 = ~(s1 ? tmp4088 : tmp4089);
  assign tmp4083 = s2 ? tmp4084 : tmp4087;
  assign tmp4082 = s3 ? tmp4083 : 1;
  assign tmp4065 = s4 ? tmp4066 : tmp4082;
  assign tmp4064 = s5 ? tmp4065 : 1;
  assign tmp4036 = s6 ? tmp4037 : tmp4064;
  assign tmp4097 = ~(l2 ? 1 : tmp3771);
  assign tmp4096 = l1 ? tmp3789 : tmp4097;
  assign tmp4099 = l1 ? tmp3486 : tmp3640;
  assign tmp4100 = l1 ? tmp3789 : tmp3435;
  assign tmp4098 = s0 ? tmp4099 : tmp4100;
  assign tmp4095 = s1 ? tmp4096 : tmp4098;
  assign tmp4104 = l1 ? tmp3863 : tmp3435;
  assign tmp4103 = s0 ? tmp4104 : tmp4096;
  assign tmp4105 = s0 ? tmp4100 : tmp4096;
  assign tmp4102 = s1 ? tmp4103 : tmp4105;
  assign tmp4107 = s0 ? tmp4100 : tmp3845;
  assign tmp4106 = s1 ? tmp4107 : tmp4096;
  assign tmp4101 = s2 ? tmp4102 : tmp4106;
  assign tmp4094 = s3 ? tmp4095 : tmp4101;
  assign tmp4111 = s0 ? tmp4104 : tmp4099;
  assign tmp4110 = s1 ? tmp4111 : tmp4096;
  assign tmp4113 = s0 ? tmp4096 : 1;
  assign tmp4115 = l1 ? tmp3486 : 0;
  assign tmp4114 = s0 ? tmp4115 : 1;
  assign tmp4112 = s1 ? tmp4113 : tmp4114;
  assign tmp4109 = s2 ? tmp4110 : tmp4112;
  assign tmp4117 = s1 ? tmp4099 : tmp3803;
  assign tmp4120 = ~(l1 ? tmp3789 : tmp4097);
  assign tmp4119 = ~(s0 ? 1 : tmp4120);
  assign tmp4118 = s1 ? tmp4096 : tmp4119;
  assign tmp4116 = s2 ? tmp4117 : tmp4118;
  assign tmp4108 = s3 ? tmp4109 : tmp4116;
  assign tmp4093 = s4 ? tmp4094 : tmp4108;
  assign tmp4126 = s0 ? tmp3845 : tmp4104;
  assign tmp4125 = s1 ? tmp4107 : tmp4126;
  assign tmp4129 = l1 ? tmp3789 : 0;
  assign tmp4128 = s0 ? tmp3845 : tmp4129;
  assign tmp4131 = l1 ? tmp3822 : tmp4097;
  assign tmp4130 = s0 ? tmp4131 : tmp3845;
  assign tmp4127 = s1 ? tmp4128 : tmp4130;
  assign tmp4124 = s2 ? tmp4125 : tmp4127;
  assign tmp4135 = l1 ? tmp3822 : tmp3435;
  assign tmp4134 = s0 ? tmp3845 : tmp4135;
  assign tmp4136 = s0 ? tmp3845 : 0;
  assign tmp4133 = s1 ? tmp4134 : tmp4136;
  assign tmp4139 = l1 ? tmp3822 : 0;
  assign tmp4138 = ~(s0 ? tmp4129 : tmp4139);
  assign tmp4137 = ~(s1 ? 1 : tmp4138);
  assign tmp4132 = s2 ? tmp4133 : tmp4137;
  assign tmp4123 = s3 ? tmp4124 : tmp4132;
  assign tmp4144 = ~(l1 ? tmp3789 : 0);
  assign tmp4143 = s0 ? 1 : tmp4144;
  assign tmp4145 = ~(s0 ? tmp4115 : tmp3512);
  assign tmp4142 = s1 ? tmp4143 : tmp4145;
  assign tmp4147 = s0 ? tmp4115 : tmp3512;
  assign tmp4149 = l1 ? tmp3863 : 0;
  assign tmp4148 = s0 ? tmp4149 : tmp4115;
  assign tmp4146 = ~(s1 ? tmp4147 : tmp4148);
  assign tmp4141 = s2 ? tmp4142 : tmp4146;
  assign tmp4152 = s0 ? 1 : tmp3914;
  assign tmp4151 = s1 ? tmp4152 : tmp3915;
  assign tmp4150 = s2 ? tmp4151 : 1;
  assign tmp4140 = ~(s3 ? tmp4141 : tmp4150);
  assign tmp4122 = s4 ? tmp4123 : tmp4140;
  assign tmp4121 = s5 ? tmp4122 : 0;
  assign tmp4092 = ~(s6 ? tmp4093 : tmp4121);
  assign tmp4035 = s8 ? tmp4036 : tmp4092;
  assign tmp4154 = s6 ? tmp4093 : tmp4121;
  assign tmp4159 = l1 ? tmp3770 : tmp3429;
  assign tmp4158 = s1 ? tmp4159 : tmp4040;
  assign tmp4163 = l1 ? tmp3781 : tmp3434;
  assign tmp4164 = ~(l1 ? tmp3548 : tmp3530);
  assign tmp4162 = s0 ? tmp4163 : tmp4164;
  assign tmp4166 = l1 ? tmp3770 : tmp3434;
  assign tmp4165 = s0 ? tmp4166 : tmp4164;
  assign tmp4161 = s1 ? tmp4162 : tmp4165;
  assign tmp4168 = s0 ? tmp4166 : tmp3434;
  assign tmp4167 = s1 ? tmp4168 : tmp4164;
  assign tmp4160 = s2 ? tmp4161 : tmp4167;
  assign tmp4157 = s3 ? tmp4158 : tmp4160;
  assign tmp4171 = s1 ? tmp4054 : tmp4164;
  assign tmp4173 = s0 ? tmp4159 : tmp3512;
  assign tmp4174 = ~(s0 ? tmp4059 : tmp3953);
  assign tmp4172 = s1 ? tmp4173 : tmp4174;
  assign tmp4170 = s2 ? tmp4171 : tmp4172;
  assign tmp4176 = s1 ? tmp4041 : tmp3956;
  assign tmp4178 = l1 ? tmp3548 : tmp3530;
  assign tmp4179 = ~(s0 ? 1 : tmp4164);
  assign tmp4177 = s1 ? tmp4178 : tmp4179;
  assign tmp4175 = ~(s2 ? tmp4176 : tmp4177);
  assign tmp4169 = s3 ? tmp4170 : tmp4175;
  assign tmp4156 = s4 ? tmp4157 : tmp4169;
  assign tmp4186 = ~(l1 ? tmp3781 : tmp3434);
  assign tmp4185 = ~(s0 ? tmp3845 : tmp4186);
  assign tmp4184 = s1 ? tmp4049 : tmp4185;
  assign tmp4189 = l1 ? 1 : tmp3429;
  assign tmp4188 = ~(s0 ? tmp4189 : tmp3475);
  assign tmp4187 = ~(s1 ? tmp4071 : tmp4188);
  assign tmp4183 = s2 ? tmp4184 : tmp4187;
  assign tmp4192 = s0 ? tmp3475 : 1;
  assign tmp4191 = s1 ? tmp3475 : tmp4192;
  assign tmp4195 = l1 ? tmp3548 : 0;
  assign tmp4194 = ~(s0 ? tmp4195 : 0);
  assign tmp4193 = s1 ? 1 : tmp4194;
  assign tmp4190 = s2 ? tmp4191 : tmp4193;
  assign tmp4182 = s3 ? tmp4183 : tmp4190;
  assign tmp4200 = ~(l1 ? tmp3548 : 0);
  assign tmp4199 = s0 ? 1 : tmp4200;
  assign tmp4198 = s1 ? tmp4199 : tmp4086;
  assign tmp4197 = s2 ? tmp4198 : tmp4087;
  assign tmp4196 = s3 ? tmp4197 : 1;
  assign tmp4181 = s4 ? tmp4182 : tmp4196;
  assign tmp4180 = s5 ? tmp4181 : 1;
  assign tmp4155 = ~(s6 ? tmp4156 : tmp4180);
  assign tmp4153 = ~(s8 ? tmp4154 : tmp4155);
  assign tmp4034 = s9 ? tmp4035 : tmp4153;
  assign tmp4207 = ~(l1 ? tmp3548 : tmp4097);
  assign tmp4206 = s0 ? tmp3781 : tmp4207;
  assign tmp4208 = s0 ? tmp4047 : tmp4207;
  assign tmp4205 = s1 ? tmp4206 : tmp4208;
  assign tmp4210 = s0 ? tmp4047 : tmp3434;
  assign tmp4209 = s1 ? tmp4210 : tmp4207;
  assign tmp4204 = s2 ? tmp4205 : tmp4209;
  assign tmp4203 = s3 ? tmp4039 : tmp4204;
  assign tmp4213 = s1 ? tmp4054 : tmp4207;
  assign tmp4215 = s0 ? tmp3770 : tmp3512;
  assign tmp4214 = s1 ? tmp4215 : tmp4174;
  assign tmp4212 = s2 ? tmp4213 : tmp4214;
  assign tmp4218 = l1 ? tmp3548 : tmp4097;
  assign tmp4219 = ~(s0 ? 1 : tmp4207);
  assign tmp4217 = s1 ? tmp4218 : tmp4219;
  assign tmp4216 = ~(s2 ? tmp4176 : tmp4217);
  assign tmp4211 = s3 ? tmp4212 : tmp4216;
  assign tmp4202 = s4 ? tmp4203 : tmp4211;
  assign tmp4225 = ~(s0 ? tmp4074 : tmp3475);
  assign tmp4224 = ~(s1 ? tmp4071 : tmp4225);
  assign tmp4223 = s2 ? tmp4068 : tmp4224;
  assign tmp4228 = s0 ? tmp3475 : tmp4078;
  assign tmp4227 = s1 ? tmp4228 : tmp4192;
  assign tmp4226 = s2 ? tmp4227 : tmp4193;
  assign tmp4222 = s3 ? tmp4223 : tmp4226;
  assign tmp4221 = s4 ? tmp4222 : tmp4196;
  assign tmp4220 = s5 ? tmp4221 : 1;
  assign tmp4201 = s6 ? tmp4202 : tmp4220;
  assign tmp4033 = s10 ? tmp4034 : tmp4201;
  assign tmp3761 = s12 ? tmp3762 : tmp4033;
  assign tmp3409 = s13 ? tmp3410 : tmp3761;
  assign tmp4238 = l1 ? 1 : tmp3772;
  assign tmp4240 = l1 ? 1 : tmp3607;
  assign tmp4239 = s0 ? tmp4240 : tmp3913;
  assign tmp4237 = s1 ? tmp4238 : tmp4239;
  assign tmp4244 = l1 ? 1 : tmp3782;
  assign tmp4245 = l1 ? 1 : tmp3783;
  assign tmp4243 = s0 ? tmp4244 : tmp4245;
  assign tmp4246 = s0 ? tmp3913 : tmp4245;
  assign tmp4242 = s1 ? tmp4243 : tmp4246;
  assign tmp4248 = s0 ? tmp3913 : tmp3460;
  assign tmp4249 = s0 ? tmp4245 : tmp4238;
  assign tmp4247 = s1 ? tmp4248 : tmp4249;
  assign tmp4241 = s2 ? tmp4242 : tmp4247;
  assign tmp4236 = s3 ? tmp4237 : tmp4241;
  assign tmp4253 = s0 ? tmp4238 : tmp4245;
  assign tmp4252 = s1 ? tmp4248 : tmp4253;
  assign tmp4255 = s0 ? tmp4238 : tmp3460;
  assign tmp4254 = s1 ? tmp4255 : tmp4248;
  assign tmp4251 = s2 ? tmp4252 : tmp4254;
  assign tmp4258 = s0 ? tmp3460 : 1;
  assign tmp4257 = s1 ? tmp4240 : tmp4258;
  assign tmp4260 = s0 ? tmp4245 : tmp3783;
  assign tmp4261 = s0 ? 1 : tmp4245;
  assign tmp4259 = s1 ? tmp4260 : tmp4261;
  assign tmp4256 = s2 ? tmp4257 : tmp4259;
  assign tmp4250 = s3 ? tmp4251 : tmp4256;
  assign tmp4235 = s4 ? tmp4236 : tmp4250;
  assign tmp4267 = s0 ? tmp3460 : tmp4244;
  assign tmp4266 = s1 ? tmp4248 : tmp4267;
  assign tmp4269 = s0 ? tmp3460 : tmp3665;
  assign tmp4270 = ~(s0 ? tmp3789 : 1);
  assign tmp4268 = s1 ? tmp4269 : tmp4270;
  assign tmp4265 = s2 ? tmp4266 : tmp4268;
  assign tmp4275 = ~(l2 ? tmp3420 : 0);
  assign tmp4274 = l1 ? 1 : tmp4275;
  assign tmp4273 = s0 ? tmp4274 : 1;
  assign tmp4272 = ~(s1 ? 1 : tmp4273);
  assign tmp4271 = ~(s2 ? tmp3818 : tmp4272);
  assign tmp4264 = s3 ? tmp4265 : tmp4271;
  assign tmp4278 = s1 ? tmp3849 : tmp4258;
  assign tmp4280 = s0 ? tmp3665 : tmp3460;
  assign tmp4279 = s1 ? tmp4258 : tmp4280;
  assign tmp4277 = s2 ? tmp4278 : tmp4279;
  assign tmp4276 = s3 ? tmp4277 : tmp3835;
  assign tmp4263 = s4 ? tmp4264 : tmp4276;
  assign tmp4262 = s5 ? tmp4263 : tmp3838;
  assign tmp4234 = s6 ? tmp4235 : tmp4262;
  assign tmp4287 = l3 ? 1 : tmp3420;
  assign tmp4286 = ~(l2 ? tmp4287 : tmp3548);
  assign tmp4285 = l1 ? 1 : tmp4286;
  assign tmp4290 = ~(l2 ? tmp4287 : 1);
  assign tmp4289 = l1 ? 1 : tmp4290;
  assign tmp4292 = ~(l2 ? tmp4287 : tmp3422);
  assign tmp4291 = l1 ? 1 : tmp4292;
  assign tmp4288 = s0 ? tmp4289 : tmp4291;
  assign tmp4284 = s1 ? tmp4285 : tmp4288;
  assign tmp4295 = s0 ? tmp4291 : tmp4245;
  assign tmp4294 = s1 ? tmp4243 : tmp4295;
  assign tmp4297 = s0 ? tmp4291 : tmp3460;
  assign tmp4298 = s0 ? tmp4245 : tmp4285;
  assign tmp4296 = s1 ? tmp4297 : tmp4298;
  assign tmp4293 = s2 ? tmp4294 : tmp4296;
  assign tmp4283 = s3 ? tmp4284 : tmp4293;
  assign tmp4302 = s0 ? tmp4285 : tmp4245;
  assign tmp4301 = s1 ? tmp4297 : tmp4302;
  assign tmp4304 = s0 ? tmp4285 : tmp3460;
  assign tmp4306 = l1 ? 1 : tmp3480;
  assign tmp4305 = s0 ? tmp4306 : tmp3460;
  assign tmp4303 = s1 ? tmp4304 : tmp4305;
  assign tmp4300 = s2 ? tmp4301 : tmp4303;
  assign tmp4308 = s1 ? tmp4289 : tmp4258;
  assign tmp4311 = ~(l1 ? 1 : tmp3783);
  assign tmp4310 = ~(s0 ? tmp3420 : tmp4311);
  assign tmp4309 = s1 ? tmp4245 : tmp4310;
  assign tmp4307 = s2 ? tmp4308 : tmp4309;
  assign tmp4299 = s3 ? tmp4300 : tmp4307;
  assign tmp4282 = s4 ? tmp4283 : tmp4299;
  assign tmp4316 = s1 ? tmp4297 : tmp4267;
  assign tmp4320 = ~(l2 ? tmp4287 : 0);
  assign tmp4319 = l1 ? 1 : tmp4320;
  assign tmp4318 = s0 ? tmp3460 : tmp4319;
  assign tmp4321 = s0 ? tmp4245 : tmp3460;
  assign tmp4317 = s1 ? tmp4318 : tmp4321;
  assign tmp4315 = s2 ? tmp4316 : tmp4317;
  assign tmp4324 = s0 ? tmp3460 : tmp4291;
  assign tmp4325 = s0 ? tmp3460 : tmp4275;
  assign tmp4323 = s1 ? tmp4324 : tmp4325;
  assign tmp4327 = ~(l1 ? 1 : tmp4275);
  assign tmp4326 = ~(s1 ? tmp3509 : tmp4327);
  assign tmp4322 = s2 ? tmp4323 : tmp4326;
  assign tmp4314 = s3 ? tmp4315 : tmp4322;
  assign tmp4331 = s0 ? 1 : tmp4319;
  assign tmp4333 = l1 ? 1 : tmp3424;
  assign tmp4332 = s0 ? tmp3460 : tmp4333;
  assign tmp4330 = s1 ? tmp4331 : tmp4332;
  assign tmp4335 = s0 ? tmp4319 : tmp3460;
  assign tmp4334 = s1 ? tmp4332 : tmp4335;
  assign tmp4329 = s2 ? tmp4330 : tmp4334;
  assign tmp4338 = s0 ? tmp4319 : tmp4274;
  assign tmp4339 = s0 ? tmp4333 : 1;
  assign tmp4337 = s1 ? tmp4338 : tmp4339;
  assign tmp4336 = s2 ? tmp4337 : 1;
  assign tmp4328 = s3 ? tmp4329 : tmp4336;
  assign tmp4313 = s4 ? tmp4314 : tmp4328;
  assign tmp4344 = ~(s0 ? 1 : tmp4333);
  assign tmp4343 = s1 ? tmp3842 : tmp4344;
  assign tmp4346 = s0 ? tmp4333 : tmp3845;
  assign tmp4345 = ~(s1 ? tmp4346 : tmp3845);
  assign tmp4342 = s2 ? tmp4343 : tmp4345;
  assign tmp4341 = s3 ? tmp4342 : 0;
  assign tmp4350 = s0 ? 1 : tmp3424;
  assign tmp4349 = s1 ? 1 : tmp4350;
  assign tmp4351 = s1 ? tmp4331 : tmp3845;
  assign tmp4348 = s2 ? tmp4349 : tmp4351;
  assign tmp4353 = s1 ? tmp4339 : 1;
  assign tmp4352 = s2 ? tmp4353 : 1;
  assign tmp4347 = ~(s3 ? tmp4348 : tmp4352);
  assign tmp4340 = ~(s4 ? tmp4341 : tmp4347);
  assign tmp4312 = s5 ? tmp4313 : tmp4340;
  assign tmp4281 = s6 ? tmp4282 : tmp4312;
  assign tmp4233 = s8 ? tmp4234 : tmp4281;
  assign tmp4360 = ~(l2 ? tmp4287 : tmp3420);
  assign tmp4359 = l1 ? 1 : tmp4360;
  assign tmp4361 = s0 ? tmp4289 : tmp4306;
  assign tmp4358 = s1 ? tmp4359 : tmp4361;
  assign tmp4364 = s0 ? tmp4289 : tmp4333;
  assign tmp4363 = s1 ? tmp4332 : tmp4364;
  assign tmp4366 = s0 ? tmp4289 : tmp3460;
  assign tmp4367 = s0 ? tmp4333 : tmp4359;
  assign tmp4365 = s1 ? tmp4366 : tmp4367;
  assign tmp4362 = s2 ? tmp4363 : tmp4365;
  assign tmp4357 = s3 ? tmp4358 : tmp4362;
  assign tmp4371 = s0 ? tmp4359 : tmp4333;
  assign tmp4370 = s1 ? tmp4305 : tmp4371;
  assign tmp4373 = s0 ? tmp4359 : tmp3460;
  assign tmp4372 = s1 ? tmp4373 : tmp4305;
  assign tmp4369 = s2 ? tmp4370 : tmp4372;
  assign tmp4377 = ~(l1 ? 1 : tmp3424);
  assign tmp4376 = ~(s0 ? tmp3420 : tmp4377);
  assign tmp4375 = s1 ? tmp4333 : tmp4376;
  assign tmp4374 = s2 ? tmp4308 : tmp4375;
  assign tmp4368 = s3 ? tmp4369 : tmp4374;
  assign tmp4356 = s4 ? tmp4357 : tmp4368;
  assign tmp4382 = s1 ? tmp4305 : tmp3460;
  assign tmp4384 = s0 ? tmp3460 : tmp4306;
  assign tmp4385 = s0 ? tmp4333 : tmp3460;
  assign tmp4383 = s1 ? tmp4384 : tmp4385;
  assign tmp4381 = s2 ? tmp4382 : tmp4383;
  assign tmp4388 = s0 ? tmp3460 : tmp4289;
  assign tmp4387 = s1 ? tmp4388 : tmp4332;
  assign tmp4389 = ~(s1 ? tmp3509 : tmp4377);
  assign tmp4386 = s2 ? tmp4387 : tmp4389;
  assign tmp4380 = s3 ? tmp4381 : tmp4386;
  assign tmp4392 = s1 ? tmp4332 : tmp4305;
  assign tmp4391 = s2 ? tmp4330 : tmp4392;
  assign tmp4395 = s0 ? tmp4306 : tmp4274;
  assign tmp4394 = s1 ? tmp4395 : tmp4339;
  assign tmp4393 = s2 ? tmp4394 : 1;
  assign tmp4390 = s3 ? tmp4391 : tmp4393;
  assign tmp4379 = s4 ? tmp4380 : tmp4390;
  assign tmp4400 = s0 ? 1 : tmp4333;
  assign tmp4399 = s1 ? tmp4339 : tmp4400;
  assign tmp4401 = s1 ? tmp4385 : tmp3460;
  assign tmp4398 = s2 ? tmp4399 : tmp4401;
  assign tmp4397 = s3 ? tmp4398 : 1;
  assign tmp4405 = s0 ? 1 : tmp4306;
  assign tmp4404 = s1 ? tmp4405 : tmp3460;
  assign tmp4403 = s2 ? tmp4349 : tmp4404;
  assign tmp4402 = s3 ? tmp4403 : tmp4352;
  assign tmp4396 = s4 ? tmp4397 : tmp4402;
  assign tmp4378 = s5 ? tmp4379 : tmp4396;
  assign tmp4355 = s6 ? tmp4356 : tmp4378;
  assign tmp4354 = s8 ? tmp4281 : tmp4355;
  assign tmp4232 = s9 ? tmp4233 : tmp4354;
  assign tmp4231 = s10 ? tmp4232 : tmp4281;
  assign tmp4415 = l3 ? 1 : tmp3424;
  assign tmp4414 = l2 ? tmp3422 : tmp4415;
  assign tmp4413 = l1 ? tmp3486 : tmp4414;
  assign tmp4418 = l2 ? 1 : tmp4415;
  assign tmp4417 = l1 ? tmp4418 : tmp4414;
  assign tmp4416 = s0 ? tmp3422 : tmp4417;
  assign tmp4412 = s1 ? tmp4413 : tmp4416;
  assign tmp4420 = s0 ? tmp3878 : tmp4417;
  assign tmp4421 = s1 ? tmp3877 : tmp4417;
  assign tmp4419 = s2 ? tmp4420 : tmp4421;
  assign tmp4411 = s3 ? tmp4412 : tmp4419;
  assign tmp4425 = s0 ? tmp4413 : tmp3830;
  assign tmp4424 = s1 ? tmp4425 : tmp4417;
  assign tmp4427 = s0 ? tmp4413 : 1;
  assign tmp4428 = s0 ? tmp3422 : 1;
  assign tmp4426 = s1 ? tmp4427 : tmp4428;
  assign tmp4423 = s2 ? tmp4424 : tmp4426;
  assign tmp4431 = s0 ? 1 : tmp3775;
  assign tmp4430 = s1 ? tmp3422 : tmp4431;
  assign tmp4435 = ~(l2 ? tmp3422 : tmp4415);
  assign tmp4434 = ~(l1 ? tmp3420 : tmp4435);
  assign tmp4433 = s0 ? tmp4417 : tmp4434;
  assign tmp4436 = s0 ? tmp3868 : tmp4417;
  assign tmp4432 = s1 ? tmp4433 : tmp4436;
  assign tmp4429 = s2 ? tmp4430 : tmp4432;
  assign tmp4422 = s3 ? tmp4423 : tmp4429;
  assign tmp4410 = s4 ? tmp4411 : tmp4422;
  assign tmp4442 = s0 ? tmp4417 : 1;
  assign tmp4443 = s0 ? 1 : tmp3878;
  assign tmp4441 = s1 ? tmp4442 : tmp4443;
  assign tmp4447 = l2 ? tmp3422 : tmp3424;
  assign tmp4446 = l1 ? tmp4418 : tmp4447;
  assign tmp4445 = s0 ? 1 : tmp4446;
  assign tmp4449 = l1 ? tmp3420 : tmp4435;
  assign tmp4448 = ~(s0 ? tmp4449 : 0);
  assign tmp4444 = s1 ? tmp4445 : tmp4448;
  assign tmp4440 = s2 ? tmp4441 : tmp4444;
  assign tmp4454 = ~(l2 ? tmp3422 : tmp3424);
  assign tmp4453 = ~(l1 ? tmp3420 : tmp4454);
  assign tmp4452 = s0 ? 1 : tmp4453;
  assign tmp4451 = s1 ? tmp4443 : tmp4452;
  assign tmp4456 = s0 ? tmp3868 : 1;
  assign tmp4457 = s0 ? tmp4446 : tmp4453;
  assign tmp4455 = s1 ? tmp4456 : tmp4457;
  assign tmp4450 = s2 ? tmp4451 : tmp4455;
  assign tmp4439 = s3 ? tmp4440 : tmp4450;
  assign tmp4461 = s0 ? tmp3868 : tmp4446;
  assign tmp4460 = s1 ? tmp4461 : tmp3832;
  assign tmp4464 = l1 ? tmp3486 : tmp4447;
  assign tmp4463 = s0 ? tmp4464 : tmp3830;
  assign tmp4462 = s1 ? tmp3832 : tmp4463;
  assign tmp4459 = s2 ? tmp4460 : tmp4462;
  assign tmp4468 = l1 ? tmp3434 : tmp4447;
  assign tmp4470 = ~(l2 ? 1 : tmp3420);
  assign tmp4469 = l1 ? tmp3486 : tmp4470;
  assign tmp4467 = s0 ? tmp4468 : tmp4469;
  assign tmp4472 = l1 ? tmp3420 : tmp4454;
  assign tmp4471 = ~(s0 ? 1 : tmp4472);
  assign tmp4466 = s1 ? tmp4467 : tmp4471;
  assign tmp4474 = s0 ? tmp3775 : 1;
  assign tmp4473 = s1 ? 1 : tmp4474;
  assign tmp4465 = s2 ? tmp4466 : tmp4473;
  assign tmp4458 = s3 ? tmp4459 : tmp4465;
  assign tmp4438 = s4 ? tmp4439 : tmp4458;
  assign tmp4479 = s0 ? tmp4472 : 0;
  assign tmp4478 = s1 ? tmp4479 : tmp3495;
  assign tmp4481 = s0 ? tmp3460 : tmp3434;
  assign tmp4482 = s0 ? tmp3512 : tmp3434;
  assign tmp4480 = ~(s1 ? tmp4481 : tmp4482);
  assign tmp4477 = s2 ? tmp4478 : tmp4480;
  assign tmp4486 = l1 ? tmp3434 : tmp4470;
  assign tmp4485 = s0 ? tmp3845 : tmp4486;
  assign tmp4484 = s1 ? tmp3844 : tmp4485;
  assign tmp4483 = ~(s2 ? tmp3514 : tmp4484);
  assign tmp4476 = s3 ? tmp4477 : tmp4483;
  assign tmp4490 = s0 ? tmp4486 : 1;
  assign tmp4491 = s0 ? 1 : tmp3868;
  assign tmp4489 = s1 ? tmp4490 : tmp4491;
  assign tmp4494 = l1 ? tmp3429 : tmp4447;
  assign tmp4493 = s0 ? 1 : tmp4494;
  assign tmp4495 = s0 ? tmp3434 : tmp3512;
  assign tmp4492 = s1 ? tmp4493 : tmp4495;
  assign tmp4488 = s2 ? tmp4489 : tmp4492;
  assign tmp4500 = l2 ? 1 : tmp3420;
  assign tmp4499 = ~(l1 ? tmp3420 : tmp4500);
  assign tmp4498 = s0 ? 1 : tmp4499;
  assign tmp4497 = s1 ? tmp4258 : tmp4498;
  assign tmp4501 = s1 ? tmp4485 : 1;
  assign tmp4496 = s2 ? tmp4497 : tmp4501;
  assign tmp4487 = ~(s3 ? tmp4488 : tmp4496);
  assign tmp4475 = ~(s4 ? tmp4476 : tmp4487);
  assign tmp4437 = s5 ? tmp4438 : tmp4475;
  assign tmp4409 = s6 ? tmp4410 : tmp4437;
  assign tmp4507 = l2 ? tmp3420 : tmp4415;
  assign tmp4506 = l1 ? tmp3486 : tmp4507;
  assign tmp4509 = l1 ? tmp3486 : tmp3544;
  assign tmp4510 = l1 ? tmp4418 : tmp4507;
  assign tmp4508 = s0 ? tmp4509 : tmp4510;
  assign tmp4505 = s1 ? tmp4506 : tmp4508;
  assign tmp4515 = l2 ? tmp4287 : tmp4415;
  assign tmp4514 = l1 ? tmp4418 : tmp4515;
  assign tmp4513 = s0 ? tmp3486 : tmp4514;
  assign tmp4517 = l1 ? tmp3486 : tmp3863;
  assign tmp4516 = s0 ? tmp4517 : tmp4514;
  assign tmp4512 = s1 ? tmp4513 : tmp4516;
  assign tmp4519 = s0 ? tmp4517 : 1;
  assign tmp4520 = s0 ? tmp4514 : tmp4510;
  assign tmp4518 = s1 ? tmp4519 : tmp4520;
  assign tmp4511 = s2 ? tmp4512 : tmp4518;
  assign tmp4504 = s3 ? tmp4505 : tmp4511;
  assign tmp4524 = s0 ? tmp4506 : tmp3685;
  assign tmp4525 = s0 ? tmp4510 : tmp4514;
  assign tmp4523 = s1 ? tmp4524 : tmp4525;
  assign tmp4527 = s0 ? tmp4506 : 1;
  assign tmp4529 = l1 ? tmp3486 : tmp3420;
  assign tmp4528 = s0 ? tmp4529 : 1;
  assign tmp4526 = s1 ? tmp4527 : tmp4528;
  assign tmp4522 = s2 ? tmp4523 : tmp4526;
  assign tmp4532 = s0 ? tmp4529 : tmp4509;
  assign tmp4531 = s1 ? tmp4532 : tmp4431;
  assign tmp4535 = l1 ? tmp3429 : tmp4515;
  assign tmp4534 = s0 ? tmp4514 : tmp4535;
  assign tmp4538 = l2 ? tmp4287 : 1;
  assign tmp4537 = l1 ? 1 : tmp4538;
  assign tmp4536 = s0 ? tmp4537 : tmp4514;
  assign tmp4533 = s1 ? tmp4534 : tmp4536;
  assign tmp4530 = s2 ? tmp4531 : tmp4533;
  assign tmp4521 = s3 ? tmp4522 : tmp4530;
  assign tmp4503 = s4 ? tmp4504 : tmp4521;
  assign tmp4544 = s0 ? tmp4510 : 1;
  assign tmp4545 = s0 ? 1 : tmp3486;
  assign tmp4543 = s1 ? tmp4544 : tmp4545;
  assign tmp4549 = l2 ? tmp3420 : tmp3424;
  assign tmp4548 = l1 ? tmp4418 : tmp4549;
  assign tmp4547 = s0 ? 1 : tmp4548;
  assign tmp4550 = s0 ? tmp4535 : 1;
  assign tmp4546 = s1 ? tmp4547 : tmp4550;
  assign tmp4542 = s2 ? tmp4543 : tmp4546;
  assign tmp4553 = s0 ? 1 : tmp4517;
  assign tmp4556 = ~(l2 ? tmp4287 : tmp3424);
  assign tmp4555 = ~(l1 ? tmp3420 : tmp4556);
  assign tmp4554 = s0 ? 1 : tmp4555;
  assign tmp4552 = s1 ? tmp4553 : tmp4554;
  assign tmp4558 = s0 ? tmp4537 : 1;
  assign tmp4561 = l2 ? tmp4287 : tmp3424;
  assign tmp4560 = l1 ? tmp4418 : tmp4561;
  assign tmp4562 = l1 ? tmp3429 : tmp4561;
  assign tmp4559 = s0 ? tmp4560 : tmp4562;
  assign tmp4557 = s1 ? tmp4558 : tmp4559;
  assign tmp4551 = s2 ? tmp4552 : tmp4557;
  assign tmp4541 = s3 ? tmp4542 : tmp4551;
  assign tmp4566 = s0 ? tmp3868 : tmp4548;
  assign tmp4567 = s0 ? tmp3685 : tmp3822;
  assign tmp4565 = s1 ? tmp4566 : tmp4567;
  assign tmp4570 = l1 ? tmp3486 : tmp4549;
  assign tmp4569 = s0 ? tmp4570 : tmp3685;
  assign tmp4568 = s1 ? tmp4567 : tmp4569;
  assign tmp4564 = s2 ? tmp4565 : tmp4568;
  assign tmp4574 = l1 ? tmp3434 : tmp4549;
  assign tmp4573 = s0 ? tmp4574 : tmp4570;
  assign tmp4575 = s0 ? tmp3822 : tmp4453;
  assign tmp4572 = s1 ? tmp4573 : tmp4575;
  assign tmp4571 = s2 ? tmp4572 : tmp4473;
  assign tmp4563 = s3 ? tmp4564 : tmp4571;
  assign tmp4540 = s4 ? tmp4541 : tmp4563;
  assign tmp4581 = l1 ? tmp3420 : tmp4556;
  assign tmp4580 = s0 ? tmp4581 : 0;
  assign tmp4583 = l1 ? 1 : tmp3420;
  assign tmp4582 = ~(s0 ? 1 : tmp4583);
  assign tmp4579 = s1 ? tmp4580 : tmp4582;
  assign tmp4585 = s0 ? tmp4583 : tmp3434;
  assign tmp4584 = ~(s1 ? tmp4585 : tmp4482);
  assign tmp4578 = s2 ? tmp4579 : tmp4584;
  assign tmp4577 = s3 ? tmp4578 : tmp4483;
  assign tmp4589 = s0 ? 1 : tmp4537;
  assign tmp4588 = s1 ? tmp4490 : tmp4589;
  assign tmp4592 = l1 ? tmp3429 : tmp4549;
  assign tmp4591 = s0 ? 1 : tmp4592;
  assign tmp4590 = s1 ? tmp4591 : tmp4495;
  assign tmp4587 = s2 ? tmp4588 : tmp4590;
  assign tmp4595 = s0 ? tmp4583 : 1;
  assign tmp4594 = s1 ? tmp4595 : tmp4498;
  assign tmp4593 = s2 ? tmp4594 : tmp4501;
  assign tmp4586 = ~(s3 ? tmp4587 : tmp4593);
  assign tmp4576 = ~(s4 ? tmp4577 : tmp4586);
  assign tmp4539 = s5 ? tmp4540 : tmp4576;
  assign tmp4502 = s6 ? tmp4503 : tmp4539;
  assign tmp4408 = s8 ? tmp4409 : tmp4502;
  assign tmp4407 = s9 ? tmp4408 : tmp4502;
  assign tmp4406 = s10 ? tmp4407 : tmp4502;
  assign tmp4230 = s12 ? tmp4231 : tmp4406;
  assign tmp4604 = l1 ? tmp3422 : tmp3421;
  assign tmp4606 = l1 ? tmp3422 : tmp3622;
  assign tmp4608 = l2 ? 1 : tmp3423;
  assign tmp4607 = ~(l1 ? tmp4608 : tmp3448);
  assign tmp4605 = s0 ? tmp4606 : tmp4607;
  assign tmp4603 = s1 ? tmp4604 : tmp4605;
  assign tmp4613 = ~(l2 ? tmp3420 : tmp3423);
  assign tmp4612 = ~(l1 ? tmp4414 : tmp4613);
  assign tmp4611 = s0 ? tmp3781 : tmp4612;
  assign tmp4615 = l1 ? tmp3781 : tmp3545;
  assign tmp4614 = s0 ? tmp4615 : tmp4612;
  assign tmp4610 = s1 ? tmp4611 : tmp4614;
  assign tmp4617 = s0 ? tmp4615 : tmp3434;
  assign tmp4619 = l1 ? tmp4414 : tmp4613;
  assign tmp4620 = l1 ? tmp4414 : tmp3421;
  assign tmp4618 = ~(s0 ? tmp4619 : tmp4620);
  assign tmp4616 = s1 ? tmp4617 : tmp4618;
  assign tmp4609 = ~(s2 ? tmp4610 : tmp4616);
  assign tmp4602 = s3 ? tmp4603 : tmp4609;
  assign tmp4625 = l1 ? tmp3781 : tmp3448;
  assign tmp4624 = s0 ? tmp4625 : tmp3781;
  assign tmp4626 = ~(s0 ? tmp4620 : tmp4619);
  assign tmp4623 = s1 ? tmp4624 : tmp4626;
  assign tmp4628 = s0 ? tmp4604 : 1;
  assign tmp4630 = l1 ? tmp3422 : tmp3436;
  assign tmp4629 = s0 ? tmp4630 : 1;
  assign tmp4627 = ~(s1 ? tmp4628 : tmp4629);
  assign tmp4622 = s2 ? tmp4623 : tmp4627;
  assign tmp4633 = s0 ? tmp4630 : tmp4606;
  assign tmp4632 = s1 ? tmp4633 : 1;
  assign tmp4636 = l1 ? tmp4447 : tmp4613;
  assign tmp4635 = s0 ? tmp4619 : tmp4636;
  assign tmp4638 = l1 ? tmp3775 : 1;
  assign tmp4637 = s0 ? tmp4638 : tmp4619;
  assign tmp4634 = s1 ? tmp4635 : tmp4637;
  assign tmp4631 = ~(s2 ? tmp4632 : tmp4634);
  assign tmp4621 = ~(s3 ? tmp4622 : tmp4631);
  assign tmp4601 = s4 ? tmp4602 : tmp4621;
  assign tmp4645 = l1 ? tmp4608 : tmp3448;
  assign tmp4644 = s0 ? tmp4645 : tmp3434;
  assign tmp4643 = s1 ? tmp4644 : tmp3781;
  assign tmp4648 = l1 ? tmp4608 : tmp4287;
  assign tmp4647 = s0 ? tmp3434 : tmp4648;
  assign tmp4649 = ~(s0 ? tmp4636 : tmp3640);
  assign tmp4646 = s1 ? tmp4647 : tmp4649;
  assign tmp4642 = s2 ? tmp4643 : tmp4646;
  assign tmp4652 = s0 ? tmp3434 : tmp4615;
  assign tmp4654 = ~(l1 ? tmp4447 : tmp3424);
  assign tmp4653 = s0 ? tmp3434 : tmp4654;
  assign tmp4651 = s1 ? tmp4652 : tmp4653;
  assign tmp4656 = s0 ? tmp4638 : 1;
  assign tmp4658 = l1 ? tmp4414 : tmp3424;
  assign tmp4659 = l1 ? tmp4447 : tmp3424;
  assign tmp4657 = s0 ? tmp4658 : tmp4659;
  assign tmp4655 = ~(s1 ? tmp4656 : tmp4657);
  assign tmp4650 = s2 ? tmp4651 : tmp4655;
  assign tmp4641 = s3 ? tmp4642 : tmp4650;
  assign tmp4664 = l1 ? tmp4414 : tmp3597;
  assign tmp4663 = s0 ? 1 : tmp4664;
  assign tmp4665 = s0 ? tmp4059 : tmp3457;
  assign tmp4662 = s1 ? tmp4663 : tmp4665;
  assign tmp4668 = l1 ? tmp3781 : tmp4287;
  assign tmp4667 = ~(s0 ? tmp4668 : tmp4091);
  assign tmp4666 = s1 ? tmp4665 : tmp4667;
  assign tmp4661 = s2 ? tmp4662 : tmp4666;
  assign tmp4672 = l1 ? 1 : tmp4287;
  assign tmp4673 = ~(l1 ? tmp3422 : tmp3429);
  assign tmp4671 = s0 ? tmp4672 : tmp4673;
  assign tmp4674 = s0 ? tmp3460 : tmp4654;
  assign tmp4670 = s1 ? tmp4671 : tmp4674;
  assign tmp4669 = ~(s2 ? tmp4670 : 0);
  assign tmp4660 = ~(s3 ? tmp4661 : tmp4669);
  assign tmp4640 = s4 ? tmp4641 : tmp4660;
  assign tmp4679 = s0 ? tmp4659 : 1;
  assign tmp4680 = s0 ? 1 : tmp3953;
  assign tmp4678 = s1 ? tmp4679 : tmp4680;
  assign tmp4681 = ~(s1 ? tmp3515 : 1);
  assign tmp4677 = s2 ? tmp4678 : tmp4681;
  assign tmp4683 = s1 ? tmp3803 : 0;
  assign tmp4686 = ~(l1 ? 1 : tmp3420);
  assign tmp4685 = s0 ? 1 : tmp4686;
  assign tmp4684 = ~(s1 ? 1 : tmp4685);
  assign tmp4682 = ~(s2 ? tmp4683 : tmp4684);
  assign tmp4676 = s3 ? tmp4677 : tmp4682;
  assign tmp4690 = s0 ? tmp4583 : tmp3512;
  assign tmp4692 = ~(l1 ? tmp3775 : 1);
  assign tmp4691 = s0 ? tmp3512 : tmp4692;
  assign tmp4689 = s1 ? tmp4690 : tmp4691;
  assign tmp4695 = ~(l1 ? tmp4500 : tmp4287);
  assign tmp4694 = s0 ? 1 : tmp4695;
  assign tmp4693 = ~(s1 ? tmp4694 : 0);
  assign tmp4688 = s2 ? tmp4689 : tmp4693;
  assign tmp4699 = l1 ? tmp4447 : tmp3429;
  assign tmp4698 = ~(s0 ? 1 : tmp4699);
  assign tmp4697 = s1 ? tmp3512 : tmp4698;
  assign tmp4700 = ~(s1 ? tmp4685 : tmp4680);
  assign tmp4696 = s2 ? tmp4697 : tmp4700;
  assign tmp4687 = ~(s3 ? tmp4688 : tmp4696);
  assign tmp4675 = ~(s4 ? tmp4676 : tmp4687);
  assign tmp4639 = ~(s5 ? tmp4640 : tmp4675);
  assign tmp4600 = s6 ? tmp4601 : tmp4639;
  assign tmp4706 = l2 ? tmp4287 : tmp3422;
  assign tmp4707 = ~(l2 ? tmp4287 : tmp3423);
  assign tmp4705 = l1 ? tmp4706 : tmp4707;
  assign tmp4709 = l1 ? tmp3486 : tmp4320;
  assign tmp4710 = l1 ? tmp4507 : tmp4707;
  assign tmp4708 = s0 ? tmp4709 : tmp4710;
  assign tmp4704 = s1 ? tmp4705 : tmp4708;
  assign tmp4714 = l1 ? tmp4515 : tmp4613;
  assign tmp4713 = s0 ? tmp4104 : tmp4714;
  assign tmp4717 = ~(l2 ? tmp4287 : tmp3436);
  assign tmp4716 = l1 ? tmp3863 : tmp4717;
  assign tmp4715 = s0 ? tmp4716 : tmp4714;
  assign tmp4712 = s1 ? tmp4713 : tmp4715;
  assign tmp4719 = s0 ? tmp4716 : tmp3845;
  assign tmp4721 = l1 ? tmp4515 : tmp4707;
  assign tmp4720 = s0 ? tmp4714 : tmp4721;
  assign tmp4718 = s1 ? tmp4719 : tmp4720;
  assign tmp4711 = s2 ? tmp4712 : tmp4718;
  assign tmp4703 = s3 ? tmp4704 : tmp4711;
  assign tmp4726 = l1 ? tmp3863 : tmp4707;
  assign tmp4725 = s0 ? tmp4726 : tmp4099;
  assign tmp4727 = s0 ? tmp4721 : tmp4714;
  assign tmp4724 = s1 ? tmp4725 : tmp4727;
  assign tmp4729 = s0 ? tmp4705 : 1;
  assign tmp4731 = l1 ? tmp3486 : tmp3480;
  assign tmp4730 = s0 ? tmp4731 : 1;
  assign tmp4728 = s1 ? tmp4729 : tmp4730;
  assign tmp4723 = s2 ? tmp4724 : tmp4728;
  assign tmp4734 = s0 ? tmp4731 : tmp4709;
  assign tmp4733 = s1 ? tmp4734 : 1;
  assign tmp4737 = l1 ? tmp4561 : tmp4613;
  assign tmp4736 = s0 ? tmp4714 : tmp4737;
  assign tmp4739 = l1 ? tmp3775 : tmp3424;
  assign tmp4738 = s0 ? tmp4739 : tmp4714;
  assign tmp4735 = s1 ? tmp4736 : tmp4738;
  assign tmp4732 = s2 ? tmp4733 : tmp4735;
  assign tmp4722 = s3 ? tmp4723 : tmp4732;
  assign tmp4702 = s4 ? tmp4703 : tmp4722;
  assign tmp4745 = s0 ? tmp4710 : tmp3640;
  assign tmp4747 = ~(l1 ? tmp3863 : tmp3435);
  assign tmp4746 = ~(s0 ? tmp3434 : tmp4747);
  assign tmp4744 = s1 ? tmp4745 : tmp4746;
  assign tmp4750 = ~(l1 ? tmp4507 : tmp3480);
  assign tmp4749 = s0 ? tmp3434 : tmp4750;
  assign tmp4751 = ~(s0 ? tmp4737 : tmp3845);
  assign tmp4748 = ~(s1 ? tmp4749 : tmp4751);
  assign tmp4743 = s2 ? tmp4744 : tmp4748;
  assign tmp4754 = s0 ? tmp3845 : tmp4716;
  assign tmp4755 = s0 ? tmp3845 : tmp4659;
  assign tmp4753 = s1 ? tmp4754 : tmp4755;
  assign tmp4757 = s0 ? tmp4739 : 1;
  assign tmp4759 = l1 ? tmp4515 : tmp3424;
  assign tmp4760 = l1 ? tmp4561 : tmp3424;
  assign tmp4758 = s0 ? tmp4759 : tmp4760;
  assign tmp4756 = s1 ? tmp4757 : tmp4758;
  assign tmp4752 = s2 ? tmp4753 : tmp4756;
  assign tmp4742 = s3 ? tmp4743 : tmp4752;
  assign tmp4765 = l1 ? tmp4515 : tmp4360;
  assign tmp4764 = s0 ? 1 : tmp4765;
  assign tmp4766 = s0 ? tmp4115 : tmp3518;
  assign tmp4763 = s1 ? tmp4764 : tmp4766;
  assign tmp4769 = l1 ? tmp3863 : tmp3480;
  assign tmp4768 = s0 ? tmp4769 : tmp4115;
  assign tmp4767 = s1 ? tmp4766 : tmp4768;
  assign tmp4762 = s2 ? tmp4763 : tmp4767;
  assign tmp4773 = ~(l1 ? tmp4706 : tmp3424);
  assign tmp4772 = s0 ? tmp4672 : tmp4773;
  assign tmp4774 = ~(s0 ? tmp3518 : tmp4659);
  assign tmp4771 = s1 ? tmp4772 : tmp4774;
  assign tmp4770 = ~(s2 ? tmp4771 : 0);
  assign tmp4761 = s3 ? tmp4762 : tmp4770;
  assign tmp4741 = s4 ? tmp4742 : tmp4761;
  assign tmp4780 = ~(l1 ? tmp3434 : tmp3420);
  assign tmp4779 = s0 ? 1 : tmp4780;
  assign tmp4778 = s1 ? tmp4679 : tmp4779;
  assign tmp4783 = l1 ? tmp3434 : tmp3420;
  assign tmp4782 = s0 ? tmp4783 : 1;
  assign tmp4781 = ~(s1 ? tmp4782 : 1);
  assign tmp4777 = s2 ? tmp4778 : tmp4781;
  assign tmp4776 = s3 ? tmp4777 : tmp4682;
  assign tmp4788 = ~(l1 ? tmp3775 : tmp3424);
  assign tmp4787 = s0 ? tmp3512 : tmp4788;
  assign tmp4786 = s1 ? tmp4690 : tmp4787;
  assign tmp4785 = s2 ? tmp4786 : tmp4693;
  assign tmp4791 = s0 ? tmp4783 : tmp3512;
  assign tmp4790 = s1 ? tmp4791 : tmp4698;
  assign tmp4789 = s2 ? tmp4790 : tmp4700;
  assign tmp4784 = ~(s3 ? tmp4785 : tmp4789);
  assign tmp4775 = s4 ? tmp4776 : tmp4784;
  assign tmp4740 = s5 ? tmp4741 : tmp4775;
  assign tmp4701 = s6 ? tmp4702 : tmp4740;
  assign tmp4599 = s8 ? tmp4600 : tmp4701;
  assign tmp4797 = l1 ? tmp4706 : tmp3622;
  assign tmp4799 = l1 ? tmp4507 : tmp3622;
  assign tmp4798 = s0 ? tmp3669 : tmp4799;
  assign tmp4796 = s1 ? tmp4797 : tmp4798;
  assign tmp4803 = l2 ? tmp4415 : tmp3436;
  assign tmp4804 = ~(l1 ? tmp4515 : tmp3630);
  assign tmp4802 = s0 ? tmp4803 : tmp4804;
  assign tmp4806 = l1 ? tmp3863 : tmp3622;
  assign tmp4807 = l1 ? tmp4515 : tmp3630;
  assign tmp4805 = ~(s0 ? tmp4806 : tmp4807);
  assign tmp4801 = s1 ? tmp4802 : tmp4805;
  assign tmp4809 = s0 ? tmp4806 : tmp3622;
  assign tmp4811 = l1 ? tmp4515 : tmp3622;
  assign tmp4810 = s0 ? tmp4807 : tmp4811;
  assign tmp4808 = ~(s1 ? tmp4809 : tmp4810);
  assign tmp4800 = ~(s2 ? tmp4801 : tmp4808);
  assign tmp4795 = s3 ? tmp4796 : tmp4800;
  assign tmp4815 = s0 ? tmp4806 : tmp4099;
  assign tmp4816 = s0 ? tmp4811 : tmp4807;
  assign tmp4814 = s1 ? tmp4815 : tmp4816;
  assign tmp4818 = s0 ? tmp4797 : 1;
  assign tmp4820 = l1 ? tmp3486 : tmp3436;
  assign tmp4819 = s0 ? tmp4820 : 1;
  assign tmp4817 = s1 ? tmp4818 : tmp4819;
  assign tmp4813 = s2 ? tmp4814 : tmp4817;
  assign tmp4823 = s0 ? tmp4820 : tmp3669;
  assign tmp4822 = s1 ? tmp4823 : 1;
  assign tmp4826 = l1 ? tmp4561 : tmp3630;
  assign tmp4825 = s0 ? tmp4807 : tmp4826;
  assign tmp4827 = s0 ? tmp4638 : tmp4807;
  assign tmp4824 = s1 ? tmp4825 : tmp4827;
  assign tmp4821 = s2 ? tmp4822 : tmp4824;
  assign tmp4812 = s3 ? tmp4813 : tmp4821;
  assign tmp4794 = s4 ? tmp4795 : tmp4812;
  assign tmp4833 = s0 ? tmp4799 : tmp3640;
  assign tmp4834 = ~(s0 ? tmp3434 : tmp4803);
  assign tmp4832 = s1 ? tmp4833 : tmp4834;
  assign tmp4837 = ~(l1 ? tmp4507 : tmp3622);
  assign tmp4836 = s0 ? tmp3434 : tmp4837;
  assign tmp4838 = ~(s0 ? tmp4826 : tmp3665);
  assign tmp4835 = ~(s1 ? tmp4836 : tmp4838);
  assign tmp4831 = s2 ? tmp4832 : tmp4835;
  assign tmp4841 = s0 ? tmp3665 : tmp4806;
  assign tmp4843 = l1 ? tmp4447 : tmp3630;
  assign tmp4842 = s0 ? tmp3665 : tmp4843;
  assign tmp4840 = s1 ? tmp4841 : tmp4842;
  assign tmp4846 = l1 ? tmp4561 : 1;
  assign tmp4845 = s0 ? tmp4807 : tmp4846;
  assign tmp4844 = s1 ? tmp4656 : tmp4845;
  assign tmp4839 = s2 ? tmp4840 : tmp4844;
  assign tmp4830 = s3 ? tmp4831 : tmp4839;
  assign tmp4850 = s0 ? 1 : tmp4811;
  assign tmp4851 = s0 ? tmp4115 : tmp3644;
  assign tmp4849 = s1 ? tmp4850 : tmp4851;
  assign tmp4853 = s0 ? tmp4806 : tmp4115;
  assign tmp4852 = s1 ? tmp4851 : tmp4853;
  assign tmp4848 = s2 ? tmp4849 : tmp4852;
  assign tmp4857 = ~(l1 ? tmp4706 : 1);
  assign tmp4856 = s0 ? tmp3426 : tmp4857;
  assign tmp4859 = l1 ? tmp4447 : 1;
  assign tmp4858 = ~(s0 ? tmp3644 : tmp4859);
  assign tmp4855 = s1 ? tmp4856 : tmp4858;
  assign tmp4854 = ~(s2 ? tmp4855 : 0);
  assign tmp4847 = s3 ? tmp4848 : tmp4854;
  assign tmp4829 = s4 ? tmp4830 : tmp4847;
  assign tmp4864 = s0 ? tmp4843 : 1;
  assign tmp4863 = s1 ? tmp4864 : tmp4680;
  assign tmp4866 = s0 ? tmp3512 : tmp3459;
  assign tmp4867 = s0 ? 1 : tmp3459;
  assign tmp4865 = ~(s1 ? tmp4866 : tmp4867);
  assign tmp4862 = s2 ? tmp4863 : tmp4865;
  assign tmp4870 = s0 ? 1 : tmp3457;
  assign tmp4869 = ~(s1 ? 1 : tmp4870);
  assign tmp4868 = ~(s2 ? tmp4683 : tmp4869);
  assign tmp4861 = s3 ? tmp4862 : tmp4868;
  assign tmp4874 = s0 ? tmp3460 : tmp3512;
  assign tmp4873 = s1 ? tmp4874 : tmp4691;
  assign tmp4877 = ~(l1 ? tmp4500 : tmp3427);
  assign tmp4876 = s0 ? 1 : tmp4877;
  assign tmp4878 = ~(s0 ? tmp3459 : 1);
  assign tmp4875 = ~(s1 ? tmp4876 : tmp4878);
  assign tmp4872 = s2 ? tmp4873 : tmp4875;
  assign tmp4881 = ~(s0 ? 1 : tmp4859);
  assign tmp4880 = s1 ? tmp3512 : tmp4881;
  assign tmp4882 = ~(s1 ? tmp4870 : tmp4680);
  assign tmp4879 = s2 ? tmp4880 : tmp4882;
  assign tmp4871 = ~(s3 ? tmp4872 : tmp4879);
  assign tmp4860 = s4 ? tmp4861 : tmp4871;
  assign tmp4828 = s5 ? tmp4829 : tmp4860;
  assign tmp4793 = s6 ? tmp4794 : tmp4828;
  assign tmp4792 = s8 ? tmp4701 : tmp4793;
  assign tmp4598 = s9 ? tmp4599 : tmp4792;
  assign tmp4887 = l1 ? tmp4706 : tmp3421;
  assign tmp4889 = l1 ? tmp4507 : tmp3421;
  assign tmp4888 = s0 ? tmp3669 : tmp4889;
  assign tmp4886 = s1 ? tmp4887 : tmp4888;
  assign tmp4893 = ~(l1 ? tmp4515 : tmp3721);
  assign tmp4892 = s0 ? tmp4803 : tmp4893;
  assign tmp4895 = l1 ? tmp3863 : tmp3441;
  assign tmp4896 = l1 ? tmp4515 : tmp3721;
  assign tmp4894 = ~(s0 ? tmp4895 : tmp4896);
  assign tmp4891 = s1 ? tmp4892 : tmp4894;
  assign tmp4898 = s0 ? tmp4895 : tmp3622;
  assign tmp4900 = l1 ? tmp4515 : tmp3421;
  assign tmp4899 = s0 ? tmp4896 : tmp4900;
  assign tmp4897 = ~(s1 ? tmp4898 : tmp4899);
  assign tmp4890 = ~(s2 ? tmp4891 : tmp4897);
  assign tmp4885 = s3 ? tmp4886 : tmp4890;
  assign tmp4905 = l1 ? tmp3863 : tmp3421;
  assign tmp4904 = s0 ? tmp4905 : tmp4099;
  assign tmp4906 = s0 ? tmp4900 : tmp4896;
  assign tmp4903 = s1 ? tmp4904 : tmp4906;
  assign tmp4908 = s0 ? tmp4887 : 1;
  assign tmp4907 = s1 ? tmp4908 : tmp4819;
  assign tmp4902 = s2 ? tmp4903 : tmp4907;
  assign tmp4912 = l1 ? tmp4561 : tmp3721;
  assign tmp4911 = s0 ? tmp4896 : tmp4912;
  assign tmp4913 = s0 ? tmp4638 : tmp4896;
  assign tmp4910 = s1 ? tmp4911 : tmp4913;
  assign tmp4909 = s2 ? tmp4822 : tmp4910;
  assign tmp4901 = s3 ? tmp4902 : tmp4909;
  assign tmp4884 = s4 ? tmp4885 : tmp4901;
  assign tmp4919 = s0 ? tmp4889 : tmp3640;
  assign tmp4918 = s1 ? tmp4919 : tmp4834;
  assign tmp4922 = ~(l1 ? tmp4507 : tmp3597);
  assign tmp4921 = s0 ? tmp3434 : tmp4922;
  assign tmp4923 = ~(s0 ? tmp4912 : tmp3665);
  assign tmp4920 = ~(s1 ? tmp4921 : tmp4923);
  assign tmp4917 = s2 ? tmp4918 : tmp4920;
  assign tmp4926 = s0 ? tmp3665 : tmp4895;
  assign tmp4928 = l1 ? tmp4447 : tmp3674;
  assign tmp4927 = s0 ? tmp3665 : tmp4928;
  assign tmp4925 = s1 ? tmp4926 : tmp4927;
  assign tmp4931 = l1 ? tmp4515 : tmp3674;
  assign tmp4932 = l1 ? tmp4561 : tmp3429;
  assign tmp4930 = s0 ? tmp4931 : tmp4932;
  assign tmp4929 = s1 ? tmp4656 : tmp4930;
  assign tmp4924 = s2 ? tmp4925 : tmp4929;
  assign tmp4916 = s3 ? tmp4917 : tmp4924;
  assign tmp4937 = l1 ? tmp4515 : tmp3597;
  assign tmp4936 = s0 ? 1 : tmp4937;
  assign tmp4935 = s1 ? tmp4936 : tmp4851;
  assign tmp4940 = l1 ? tmp3863 : tmp3597;
  assign tmp4939 = s0 ? tmp4940 : tmp4115;
  assign tmp4938 = s1 ? tmp4851 : tmp4939;
  assign tmp4934 = s2 ? tmp4935 : tmp4938;
  assign tmp4944 = l1 ? 1 : tmp3494;
  assign tmp4945 = ~(l1 ? tmp4706 : tmp3429);
  assign tmp4943 = s0 ? tmp4944 : tmp4945;
  assign tmp4946 = ~(s0 ? tmp3644 : tmp4659);
  assign tmp4942 = s1 ? tmp4943 : tmp4946;
  assign tmp4941 = ~(s2 ? tmp4942 : 0);
  assign tmp4933 = s3 ? tmp4934 : tmp4941;
  assign tmp4915 = s4 ? tmp4916 : tmp4933;
  assign tmp4951 = s0 ? tmp4928 : 1;
  assign tmp4950 = s1 ? tmp4951 : tmp4680;
  assign tmp4953 = s0 ? tmp3512 : tmp3868;
  assign tmp4952 = ~(s1 ? tmp4953 : tmp4491);
  assign tmp4949 = s2 ? tmp4950 : tmp4952;
  assign tmp4948 = s3 ? tmp4949 : tmp4682;
  assign tmp4958 = ~(l1 ? tmp4500 : tmp3494);
  assign tmp4957 = s0 ? 1 : tmp4958;
  assign tmp4959 = ~(s0 ? tmp3868 : 1);
  assign tmp4956 = ~(s1 ? tmp4957 : tmp4959);
  assign tmp4955 = s2 ? tmp4689 : tmp4956;
  assign tmp4954 = ~(s3 ? tmp4955 : tmp4696);
  assign tmp4947 = s4 ? tmp4948 : tmp4954;
  assign tmp4914 = s5 ? tmp4915 : tmp4947;
  assign tmp4883 = s6 ? tmp4884 : tmp4914;
  assign tmp4597 = s10 ? tmp4598 : tmp4883;
  assign tmp4967 = l1 ? tmp3422 : tmp4418;
  assign tmp4969 = ~(l1 ? tmp4608 : tmp3423);
  assign tmp4968 = s0 ? tmp3830 : tmp4969;
  assign tmp4966 = s1 ? tmp4967 : tmp4968;
  assign tmp4973 = ~(l1 ? tmp4414 : tmp4415);
  assign tmp4972 = s0 ? tmp3795 : tmp4973;
  assign tmp4974 = s0 ? tmp3780 : tmp4973;
  assign tmp4971 = s1 ? tmp4972 : tmp4974;
  assign tmp4976 = s0 ? tmp3780 : 0;
  assign tmp4978 = l1 ? tmp4414 : tmp4415;
  assign tmp4979 = l1 ? tmp4414 : tmp4418;
  assign tmp4977 = ~(s0 ? tmp4978 : tmp4979);
  assign tmp4975 = s1 ? tmp4976 : tmp4977;
  assign tmp4970 = ~(s2 ? tmp4971 : tmp4975);
  assign tmp4965 = s3 ? tmp4966 : tmp4970;
  assign tmp4984 = l1 ? tmp3781 : tmp3423;
  assign tmp4983 = s0 ? tmp4984 : tmp3796;
  assign tmp4985 = ~(s0 ? tmp4979 : tmp4978);
  assign tmp4982 = s1 ? tmp4983 : tmp4985;
  assign tmp4987 = s0 ? tmp4967 : 1;
  assign tmp4988 = s0 ? tmp3830 : 1;
  assign tmp4986 = ~(s1 ? tmp4987 : tmp4988);
  assign tmp4981 = s2 ? tmp4982 : tmp4986;
  assign tmp4990 = s1 ? tmp3830 : 1;
  assign tmp4993 = l1 ? tmp4447 : tmp4415;
  assign tmp4992 = s0 ? tmp4978 : tmp4993;
  assign tmp4994 = s0 ? tmp4638 : tmp4978;
  assign tmp4991 = s1 ? tmp4992 : tmp4994;
  assign tmp4989 = ~(s2 ? tmp4990 : tmp4991);
  assign tmp4980 = ~(s3 ? tmp4981 : tmp4989);
  assign tmp4964 = s4 ? tmp4965 : tmp4980;
  assign tmp5001 = l1 ? tmp4608 : tmp3423;
  assign tmp5000 = s0 ? tmp5001 : 0;
  assign tmp4999 = s1 ? tmp5000 : tmp3795;
  assign tmp5004 = ~(l1 ? tmp4608 : tmp3530);
  assign tmp5003 = s0 ? 1 : tmp5004;
  assign tmp5005 = s0 ? tmp4993 : 1;
  assign tmp5002 = ~(s1 ? tmp5003 : tmp5005);
  assign tmp4998 = s2 ? tmp4999 : tmp5002;
  assign tmp5008 = s0 ? 1 : tmp3812;
  assign tmp5009 = s0 ? 1 : tmp4699;
  assign tmp5007 = s1 ? tmp5008 : tmp5009;
  assign tmp5012 = l1 ? tmp4414 : tmp3429;
  assign tmp5011 = s0 ? tmp5012 : tmp4659;
  assign tmp5010 = s1 ? tmp4656 : tmp5011;
  assign tmp5006 = ~(s2 ? tmp5007 : tmp5010);
  assign tmp4997 = s3 ? tmp4998 : tmp5006;
  assign tmp5016 = s0 ? 1 : tmp5012;
  assign tmp5017 = s0 ? tmp3830 : tmp3457;
  assign tmp5015 = s1 ? tmp5016 : tmp5017;
  assign tmp5020 = l1 ? tmp3781 : tmp3530;
  assign tmp5019 = ~(s0 ? tmp5020 : tmp3796);
  assign tmp5018 = s1 ? tmp5017 : tmp5019;
  assign tmp5014 = s2 ? tmp5015 : tmp5018;
  assign tmp5024 = l1 ? 1 : tmp3530;
  assign tmp5023 = s0 ? tmp5024 : tmp4673;
  assign tmp5022 = s1 ? tmp5023 : tmp4674;
  assign tmp5021 = ~(s2 ? tmp5022 : 0);
  assign tmp5013 = ~(s3 ? tmp5014 : tmp5021);
  assign tmp4996 = s4 ? tmp4997 : tmp5013;
  assign tmp5029 = s0 ? tmp4699 : 1;
  assign tmp5028 = s1 ? tmp5029 : tmp4680;
  assign tmp5031 = s0 ? tmp3512 : tmp3845;
  assign tmp5030 = ~(s1 ? tmp5031 : tmp3844);
  assign tmp5027 = s2 ? tmp5028 : tmp5030;
  assign tmp5026 = s3 ? tmp5027 : tmp4682;
  assign tmp5036 = ~(l1 ? tmp4500 : tmp3530);
  assign tmp5035 = s0 ? 1 : tmp5036;
  assign tmp5037 = ~(s0 ? tmp3845 : 1);
  assign tmp5034 = ~(s1 ? tmp5035 : tmp5037);
  assign tmp5033 = s2 ? tmp4689 : tmp5034;
  assign tmp5032 = ~(s3 ? tmp5033 : tmp4696);
  assign tmp5025 = ~(s4 ? tmp5026 : tmp5032);
  assign tmp4995 = ~(s5 ? tmp4996 : tmp5025);
  assign tmp4963 = s6 ? tmp4964 : tmp4995;
  assign tmp5042 = l1 ? tmp4706 : tmp4415;
  assign tmp5045 = l2 ? tmp4415 : 1;
  assign tmp5044 = l1 ? tmp3486 : tmp5045;
  assign tmp5046 = l1 ? tmp4507 : tmp4415;
  assign tmp5043 = s0 ? tmp5044 : tmp5046;
  assign tmp5041 = s1 ? tmp5042 : tmp5043;
  assign tmp5050 = l1 ? tmp4515 : tmp4415;
  assign tmp5049 = s0 ? tmp3862 : tmp5050;
  assign tmp5053 = l2 ? tmp4415 : tmp3422;
  assign tmp5052 = l1 ? tmp3863 : tmp5053;
  assign tmp5051 = s0 ? tmp5052 : tmp5050;
  assign tmp5048 = s1 ? tmp5049 : tmp5051;
  assign tmp5055 = s0 ? tmp5052 : tmp3459;
  assign tmp5054 = s1 ? tmp5055 : tmp5050;
  assign tmp5047 = s2 ? tmp5048 : tmp5054;
  assign tmp5040 = s3 ? tmp5041 : tmp5047;
  assign tmp5060 = l1 ? tmp3863 : tmp4415;
  assign tmp5059 = s0 ? tmp5060 : tmp3685;
  assign tmp5058 = s1 ? tmp5059 : tmp5050;
  assign tmp5062 = s0 ? tmp5042 : 1;
  assign tmp5064 = l1 ? tmp3486 : tmp4415;
  assign tmp5063 = s0 ? tmp5064 : 1;
  assign tmp5061 = s1 ? tmp5062 : tmp5063;
  assign tmp5057 = s2 ? tmp5058 : tmp5061;
  assign tmp5067 = s0 ? tmp5064 : tmp5044;
  assign tmp5066 = s1 ? tmp5067 : 1;
  assign tmp5070 = l1 ? tmp4561 : tmp4415;
  assign tmp5069 = s0 ? tmp5050 : tmp5070;
  assign tmp5071 = s0 ? tmp4739 : tmp5050;
  assign tmp5068 = s1 ? tmp5069 : tmp5071;
  assign tmp5065 = s2 ? tmp5066 : tmp5068;
  assign tmp5056 = s3 ? tmp5057 : tmp5065;
  assign tmp5039 = s4 ? tmp5040 : tmp5056;
  assign tmp5077 = s0 ? tmp5046 : 1;
  assign tmp5076 = s1 ? tmp5077 : tmp3890;
  assign tmp5081 = l2 ? tmp4415 : tmp3424;
  assign tmp5080 = l1 ? tmp4507 : tmp5081;
  assign tmp5079 = s0 ? 1 : tmp5080;
  assign tmp5082 = s0 ? tmp5070 : tmp3459;
  assign tmp5078 = s1 ? tmp5079 : tmp5082;
  assign tmp5075 = s2 ? tmp5076 : tmp5078;
  assign tmp5085 = s0 ? tmp3459 : tmp5052;
  assign tmp5087 = l1 ? tmp4447 : tmp5081;
  assign tmp5086 = s0 ? tmp3459 : tmp5087;
  assign tmp5084 = s1 ? tmp5085 : tmp5086;
  assign tmp5090 = l1 ? tmp4515 : tmp5081;
  assign tmp5089 = s0 ? tmp5090 : tmp4760;
  assign tmp5088 = s1 ? tmp4757 : tmp5089;
  assign tmp5083 = s2 ? tmp5084 : tmp5088;
  assign tmp5074 = s3 ? tmp5075 : tmp5083;
  assign tmp5094 = s0 ? 1 : tmp5090;
  assign tmp5095 = s0 ? tmp3685 : tmp3518;
  assign tmp5093 = s1 ? tmp5094 : tmp5095;
  assign tmp5098 = l1 ? tmp3863 : tmp5081;
  assign tmp5097 = s0 ? tmp5098 : tmp3685;
  assign tmp5096 = s1 ? tmp5095 : tmp5097;
  assign tmp5092 = s2 ? tmp5093 : tmp5096;
  assign tmp5103 = ~(l2 ? tmp4415 : tmp3424);
  assign tmp5102 = l1 ? 1 : tmp5103;
  assign tmp5101 = s0 ? tmp5102 : tmp4773;
  assign tmp5100 = s1 ? tmp5101 : tmp4774;
  assign tmp5099 = ~(s2 ? tmp5100 : 0);
  assign tmp5091 = s3 ? tmp5092 : tmp5099;
  assign tmp5073 = s4 ? tmp5074 : tmp5091;
  assign tmp5108 = s0 ? tmp5087 : 1;
  assign tmp5107 = s1 ? tmp5108 : tmp4779;
  assign tmp5110 = s0 ? tmp4783 : tmp3665;
  assign tmp5109 = ~(s1 ? tmp5110 : tmp3849);
  assign tmp5106 = s2 ? tmp5107 : tmp5109;
  assign tmp5105 = s3 ? tmp5106 : tmp4682;
  assign tmp5115 = ~(l1 ? tmp4500 : tmp5103);
  assign tmp5114 = s0 ? 1 : tmp5115;
  assign tmp5116 = ~(s0 ? tmp3665 : 1);
  assign tmp5113 = ~(s1 ? tmp5114 : tmp5116);
  assign tmp5112 = s2 ? tmp4786 : tmp5113;
  assign tmp5111 = ~(s3 ? tmp5112 : tmp4789);
  assign tmp5104 = s4 ? tmp5105 : tmp5111;
  assign tmp5072 = s5 ? tmp5073 : tmp5104;
  assign tmp5038 = s6 ? tmp5039 : tmp5072;
  assign tmp4962 = s8 ? tmp4963 : tmp5038;
  assign tmp5122 = l1 ? tmp4706 : 1;
  assign tmp5124 = l1 ? tmp4507 : 1;
  assign tmp5123 = s0 ? tmp3685 : tmp5124;
  assign tmp5121 = s1 ? tmp5122 : tmp5123;
  assign tmp5127 = l1 ? tmp3863 : 1;
  assign tmp5128 = l1 ? tmp4515 : 1;
  assign tmp5126 = s0 ? tmp5127 : tmp5128;
  assign tmp5130 = s0 ? tmp5127 : 1;
  assign tmp5129 = s1 ? tmp5130 : tmp5128;
  assign tmp5125 = s2 ? tmp5126 : tmp5129;
  assign tmp5120 = s3 ? tmp5121 : tmp5125;
  assign tmp5134 = s0 ? tmp5127 : tmp3685;
  assign tmp5133 = s1 ? tmp5134 : tmp5128;
  assign tmp5136 = s0 ? tmp5122 : 1;
  assign tmp5137 = s0 ? tmp3685 : 1;
  assign tmp5135 = s1 ? tmp5136 : tmp5137;
  assign tmp5132 = s2 ? tmp5133 : tmp5135;
  assign tmp5139 = s1 ? tmp3685 : 1;
  assign tmp5141 = s0 ? tmp5128 : tmp4846;
  assign tmp5142 = s0 ? tmp4638 : tmp5128;
  assign tmp5140 = s1 ? tmp5141 : tmp5142;
  assign tmp5138 = s2 ? tmp5139 : tmp5140;
  assign tmp5131 = s3 ? tmp5132 : tmp5138;
  assign tmp5119 = s4 ? tmp5120 : tmp5131;
  assign tmp5148 = s0 ? tmp5124 : 1;
  assign tmp5149 = s0 ? 1 : tmp5127;
  assign tmp5147 = s1 ? tmp5148 : tmp5149;
  assign tmp5151 = s0 ? 1 : tmp5124;
  assign tmp5152 = s0 ? tmp4846 : 1;
  assign tmp5150 = s1 ? tmp5151 : tmp5152;
  assign tmp5146 = s2 ? tmp5147 : tmp5150;
  assign tmp5155 = s0 ? 1 : tmp4859;
  assign tmp5154 = s1 ? tmp5149 : tmp5155;
  assign tmp5156 = s1 ? tmp4656 : tmp5141;
  assign tmp5153 = s2 ? tmp5154 : tmp5156;
  assign tmp5145 = s3 ? tmp5146 : tmp5153;
  assign tmp5160 = s0 ? 1 : tmp5128;
  assign tmp5161 = s0 ? tmp3685 : tmp3644;
  assign tmp5159 = s1 ? tmp5160 : tmp5161;
  assign tmp5162 = s1 ? tmp5161 : tmp5134;
  assign tmp5158 = s2 ? tmp5159 : tmp5162;
  assign tmp5165 = s0 ? tmp3460 : tmp4857;
  assign tmp5164 = s1 ? tmp5165 : tmp4858;
  assign tmp5163 = ~(s2 ? tmp5164 : 0);
  assign tmp5157 = s3 ? tmp5158 : tmp5163;
  assign tmp5144 = s4 ? tmp5145 : tmp5157;
  assign tmp5170 = s0 ? tmp4859 : 1;
  assign tmp5169 = s1 ? tmp5170 : tmp4680;
  assign tmp5172 = s0 ? tmp3512 : tmp3460;
  assign tmp5171 = ~(s1 ? tmp5172 : tmp3497);
  assign tmp5168 = s2 ? tmp5169 : tmp5171;
  assign tmp5167 = s3 ? tmp5168 : tmp4868;
  assign tmp5177 = ~(l1 ? tmp4500 : 0);
  assign tmp5176 = s0 ? 1 : tmp5177;
  assign tmp5178 = ~(s0 ? tmp3460 : 1);
  assign tmp5175 = ~(s1 ? tmp5176 : tmp5178);
  assign tmp5174 = s2 ? tmp4873 : tmp5175;
  assign tmp5173 = ~(s3 ? tmp5174 : tmp4879);
  assign tmp5166 = s4 ? tmp5167 : tmp5173;
  assign tmp5143 = s5 ? tmp5144 : tmp5166;
  assign tmp5118 = s6 ? tmp5119 : tmp5143;
  assign tmp5117 = s8 ? tmp5038 : tmp5118;
  assign tmp4961 = s9 ? tmp4962 : tmp5117;
  assign tmp5183 = l1 ? tmp4706 : tmp4418;
  assign tmp5185 = l1 ? tmp4507 : tmp4418;
  assign tmp5184 = s0 ? tmp3685 : tmp5185;
  assign tmp5182 = s1 ? tmp5183 : tmp5184;
  assign tmp5188 = l1 ? tmp3863 : tmp3486;
  assign tmp5189 = l1 ? tmp4515 : tmp4418;
  assign tmp5187 = s0 ? tmp5188 : tmp5189;
  assign tmp5191 = s0 ? tmp5188 : 1;
  assign tmp5190 = s1 ? tmp5191 : tmp5189;
  assign tmp5186 = s2 ? tmp5187 : tmp5190;
  assign tmp5181 = s3 ? tmp5182 : tmp5186;
  assign tmp5196 = l1 ? tmp3863 : tmp4418;
  assign tmp5195 = s0 ? tmp5196 : tmp3685;
  assign tmp5194 = s1 ? tmp5195 : tmp5189;
  assign tmp5198 = s0 ? tmp5183 : 1;
  assign tmp5197 = s1 ? tmp5198 : tmp5137;
  assign tmp5193 = s2 ? tmp5194 : tmp5197;
  assign tmp5202 = l1 ? tmp4561 : tmp4418;
  assign tmp5201 = s0 ? tmp5189 : tmp5202;
  assign tmp5203 = s0 ? tmp4638 : tmp5189;
  assign tmp5200 = s1 ? tmp5201 : tmp5203;
  assign tmp5199 = s2 ? tmp5139 : tmp5200;
  assign tmp5192 = s3 ? tmp5193 : tmp5199;
  assign tmp5180 = s4 ? tmp5181 : tmp5192;
  assign tmp5209 = s0 ? tmp5185 : 1;
  assign tmp5210 = s0 ? 1 : tmp5188;
  assign tmp5208 = s1 ? tmp5209 : tmp5210;
  assign tmp5213 = l1 ? tmp4507 : tmp3429;
  assign tmp5212 = s0 ? 1 : tmp5213;
  assign tmp5214 = s0 ? tmp5202 : 1;
  assign tmp5211 = s1 ? tmp5212 : tmp5214;
  assign tmp5207 = s2 ? tmp5208 : tmp5211;
  assign tmp5216 = s1 ? tmp5210 : tmp5009;
  assign tmp5219 = l1 ? tmp4515 : tmp3429;
  assign tmp5218 = s0 ? tmp5219 : tmp4932;
  assign tmp5217 = s1 ? tmp4656 : tmp5218;
  assign tmp5215 = s2 ? tmp5216 : tmp5217;
  assign tmp5206 = s3 ? tmp5207 : tmp5215;
  assign tmp5223 = s0 ? 1 : tmp5219;
  assign tmp5222 = s1 ? tmp5223 : tmp5161;
  assign tmp5226 = l1 ? tmp3863 : tmp3429;
  assign tmp5225 = s0 ? tmp5226 : tmp3685;
  assign tmp5224 = s1 ? tmp5161 : tmp5225;
  assign tmp5221 = s2 ? tmp5222 : tmp5224;
  assign tmp5229 = s0 ? tmp5024 : tmp4945;
  assign tmp5228 = s1 ? tmp5229 : tmp4946;
  assign tmp5227 = ~(s2 ? tmp5228 : 0);
  assign tmp5220 = s3 ? tmp5221 : tmp5227;
  assign tmp5205 = s4 ? tmp5206 : tmp5220;
  assign tmp5230 = s4 ? tmp5026 : tmp5032;
  assign tmp5204 = s5 ? tmp5205 : tmp5230;
  assign tmp5179 = s6 ? tmp5180 : tmp5204;
  assign tmp4960 = s10 ? tmp4961 : tmp5179;
  assign tmp4596 = s12 ? tmp4597 : tmp4960;
  assign tmp4229 = s13 ? tmp4230 : tmp4596;
  assign tmp3408 = s14 ? tmp3409 : tmp4229;
  assign tmp5241 = l1 ? tmp4447 : 0;
  assign tmp5244 = l2 ? 1 : tmp3538;
  assign tmp5243 = l1 ? tmp5244 : 1;
  assign tmp5242 = ~(s0 ? 1 : tmp5243);
  assign tmp5240 = s1 ? tmp5241 : tmp5242;
  assign tmp5249 = l2 ? tmp3422 : tmp3419;
  assign tmp5250 = ~(l2 ? tmp3538 : 1);
  assign tmp5248 = ~(l1 ? tmp5249 : tmp5250);
  assign tmp5247 = s0 ? 1 : tmp5248;
  assign tmp5252 = l1 ? tmp4500 : 1;
  assign tmp5251 = s0 ? tmp5252 : tmp5248;
  assign tmp5246 = s1 ? tmp5247 : tmp5251;
  assign tmp5254 = s0 ? tmp5252 : 1;
  assign tmp5253 = s1 ? tmp5254 : tmp5248;
  assign tmp5245 = ~(s2 ? tmp5246 : tmp5253);
  assign tmp5239 = s3 ? tmp5240 : tmp5245;
  assign tmp5257 = s1 ? 1 : tmp5248;
  assign tmp5259 = s0 ? tmp5241 : 0;
  assign tmp5258 = ~(s1 ? tmp5259 : 0);
  assign tmp5256 = s2 ? tmp5257 : tmp5258;
  assign tmp5263 = ~(l1 ? tmp3486 : tmp3427);
  assign tmp5262 = s0 ? 1 : tmp5263;
  assign tmp5261 = s1 ? 1 : tmp5262;
  assign tmp5266 = l1 ? tmp5249 : tmp5250;
  assign tmp5267 = l1 ? tmp3422 : tmp5250;
  assign tmp5265 = s0 ? tmp5266 : tmp5267;
  assign tmp5269 = l1 ? tmp3422 : tmp3427;
  assign tmp5268 = s0 ? tmp5269 : tmp5266;
  assign tmp5264 = ~(s1 ? tmp5265 : tmp5268);
  assign tmp5260 = s2 ? tmp5261 : tmp5264;
  assign tmp5255 = ~(s3 ? tmp5256 : tmp5260);
  assign tmp5238 = s4 ? tmp5239 : tmp5255;
  assign tmp5275 = s0 ? tmp5243 : 1;
  assign tmp5274 = s1 ? tmp5275 : 1;
  assign tmp5277 = s0 ? 1 : tmp5243;
  assign tmp5278 = ~(s0 ? tmp5267 : 0);
  assign tmp5276 = s1 ? tmp5277 : tmp5278;
  assign tmp5273 = s2 ? tmp5274 : tmp5276;
  assign tmp5281 = s0 ? 1 : tmp4090;
  assign tmp5283 = ~(l1 ? tmp3422 : tmp5250);
  assign tmp5282 = s0 ? 1 : tmp5283;
  assign tmp5280 = s1 ? tmp5281 : tmp5282;
  assign tmp5286 = l1 ? tmp3486 : tmp3434;
  assign tmp5285 = s0 ? tmp5269 : tmp5286;
  assign tmp5287 = s0 ? tmp5266 : tmp5269;
  assign tmp5284 = ~(s1 ? tmp5285 : tmp5287);
  assign tmp5279 = s2 ? tmp5280 : tmp5284;
  assign tmp5272 = s3 ? tmp5273 : tmp5279;
  assign tmp5292 = l1 ? tmp5249 : 0;
  assign tmp5291 = s0 ? tmp3426 : tmp5292;
  assign tmp5290 = s1 ? tmp5291 : 0;
  assign tmp5289 = s2 ? tmp5290 : 0;
  assign tmp5295 = s0 ? 1 : tmp4091;
  assign tmp5297 = ~(l1 ? tmp3422 : tmp3427);
  assign tmp5296 = s0 ? 1 : tmp5297;
  assign tmp5294 = s1 ? tmp5295 : tmp5296;
  assign tmp5300 = l1 ? tmp3486 : tmp3427;
  assign tmp5299 = s0 ? tmp5300 : tmp3475;
  assign tmp5298 = ~(s1 ? tmp3475 : tmp5299);
  assign tmp5293 = ~(s2 ? tmp5294 : tmp5298);
  assign tmp5288 = ~(s3 ? tmp5289 : tmp5293);
  assign tmp5271 = s4 ? tmp5272 : tmp5288;
  assign tmp5305 = s0 ? tmp5267 : 1;
  assign tmp5306 = s0 ? 1 : tmp3640;
  assign tmp5304 = s1 ? tmp5305 : tmp5306;
  assign tmp5307 = ~(s1 ? tmp3698 : 1);
  assign tmp5303 = s2 ? tmp5304 : tmp5307;
  assign tmp5311 = ~(l1 ? tmp3422 : tmp3434);
  assign tmp5310 = s0 ? 1 : tmp5311;
  assign tmp5309 = s1 ? 1 : tmp5310;
  assign tmp5314 = l1 ? tmp3422 : tmp3434;
  assign tmp5313 = s0 ? tmp5314 : tmp3460;
  assign tmp5312 = ~(s1 ? tmp5313 : tmp3464);
  assign tmp5308 = ~(s2 ? tmp5309 : tmp5312);
  assign tmp5302 = s3 ? tmp5303 : tmp5308;
  assign tmp5318 = ~(s0 ? tmp4059 : tmp5269);
  assign tmp5317 = s1 ? tmp5295 : tmp5318;
  assign tmp5321 = ~(l1 ? tmp3781 : 1);
  assign tmp5320 = s0 ? 1 : tmp5321;
  assign tmp5319 = ~(s1 ? tmp5320 : 0);
  assign tmp5316 = s2 ? tmp5317 : tmp5319;
  assign tmp5324 = s0 ? tmp3434 : tmp5311;
  assign tmp5325 = ~(s0 ? tmp5314 : tmp4059);
  assign tmp5323 = s1 ? tmp5324 : tmp5325;
  assign tmp5327 = ~(s0 ? 1 : tmp4091);
  assign tmp5326 = ~(s1 ? tmp3464 : tmp5327);
  assign tmp5322 = s2 ? tmp5323 : tmp5326;
  assign tmp5315 = ~(s3 ? tmp5316 : tmp5322);
  assign tmp5301 = ~(s4 ? tmp5302 : tmp5315);
  assign tmp5270 = ~(s5 ? tmp5271 : tmp5301);
  assign tmp5237 = s6 ? tmp5238 : tmp5270;
  assign tmp5335 = ~(l1 ? tmp3434 : 1);
  assign tmp5334 = s0 ? 1 : tmp5335;
  assign tmp5333 = s1 ? tmp5305 : tmp5334;
  assign tmp5336 = ~(s1 ? tmp3650 : 1);
  assign tmp5332 = s2 ? tmp5333 : tmp5336;
  assign tmp5331 = s3 ? tmp5332 : tmp5308;
  assign tmp5340 = s0 ? tmp3644 : tmp5311;
  assign tmp5339 = s1 ? tmp5340 : tmp5325;
  assign tmp5338 = s2 ? tmp5339 : tmp5326;
  assign tmp5337 = ~(s3 ? tmp5316 : tmp5338);
  assign tmp5330 = ~(s4 ? tmp5331 : tmp5337);
  assign tmp5329 = ~(s5 ? tmp5271 : tmp5330);
  assign tmp5328 = s6 ? tmp5238 : tmp5329;
  assign tmp5236 = s8 ? tmp5237 : tmp5328;
  assign tmp5235 = s9 ? tmp5236 : tmp5328;
  assign tmp5234 = s10 ? tmp5235 : tmp5328;
  assign tmp5349 = ~(l2 ? 1 : tmp3538);
  assign tmp5348 = l1 ? tmp3427 : tmp5349;
  assign tmp5347 = s1 ? tmp5348 : 0;
  assign tmp5352 = ~(l1 ? tmp3427 : tmp3419);
  assign tmp5351 = s0 ? 1 : tmp5352;
  assign tmp5353 = s1 ? 1 : tmp5352;
  assign tmp5350 = ~(s2 ? tmp5351 : tmp5353);
  assign tmp5346 = s3 ? tmp5347 : tmp5350;
  assign tmp5357 = s0 ? tmp5348 : 0;
  assign tmp5356 = ~(s1 ? tmp5357 : 0);
  assign tmp5355 = s2 ? tmp5353 : tmp5356;
  assign tmp5361 = ~(l1 ? tmp3434 : tmp3422);
  assign tmp5360 = s0 ? 1 : tmp5361;
  assign tmp5359 = s1 ? 1 : tmp5360;
  assign tmp5363 = l1 ? tmp3427 : tmp3419;
  assign tmp5365 = l1 ? tmp3427 : tmp3422;
  assign tmp5364 = s0 ? tmp5365 : tmp5363;
  assign tmp5362 = ~(s1 ? tmp5363 : tmp5364);
  assign tmp5358 = s2 ? tmp5359 : tmp5362;
  assign tmp5354 = ~(s3 ? tmp5355 : tmp5358);
  assign tmp5345 = s4 ? tmp5346 : tmp5354;
  assign tmp5371 = ~(s0 ? tmp5363 : 0);
  assign tmp5370 = s1 ? 1 : tmp5371;
  assign tmp5369 = s2 ? 1 : tmp5370;
  assign tmp5376 = ~(l2 ? tmp3538 : tmp3436);
  assign tmp5375 = ~(l1 ? tmp3427 : tmp5376);
  assign tmp5374 = s0 ? 1 : tmp5375;
  assign tmp5373 = s1 ? 1 : tmp5374;
  assign tmp5378 = s0 ? tmp5365 : tmp3644;
  assign tmp5380 = l1 ? tmp3427 : tmp5376;
  assign tmp5379 = s0 ? tmp5380 : tmp5365;
  assign tmp5377 = ~(s1 ? tmp5378 : tmp5379);
  assign tmp5372 = s2 ? tmp5373 : tmp5377;
  assign tmp5368 = s3 ? tmp5369 : tmp5372;
  assign tmp5385 = l1 ? tmp3434 : tmp3422;
  assign tmp5386 = l1 ? tmp3427 : tmp3435;
  assign tmp5384 = s0 ? tmp5385 : tmp5386;
  assign tmp5383 = s1 ? tmp5384 : 0;
  assign tmp5382 = s2 ? tmp5383 : 0;
  assign tmp5390 = ~(l1 ? tmp3427 : tmp3435);
  assign tmp5389 = s0 ? 1 : tmp5390;
  assign tmp5392 = ~(l1 ? tmp3427 : tmp3422);
  assign tmp5391 = s0 ? 1 : tmp5392;
  assign tmp5388 = s1 ? tmp5389 : tmp5391;
  assign tmp5394 = s0 ? tmp5385 : 1;
  assign tmp5393 = ~(s1 ? 1 : tmp5394);
  assign tmp5387 = ~(s2 ? tmp5388 : tmp5393);
  assign tmp5381 = ~(s3 ? tmp5382 : tmp5387);
  assign tmp5367 = s4 ? tmp5368 : tmp5381;
  assign tmp5399 = s0 ? tmp5380 : tmp3644;
  assign tmp5400 = s0 ? tmp3644 : 0;
  assign tmp5398 = s1 ? tmp5399 : tmp5400;
  assign tmp5397 = s2 ? tmp5398 : 0;
  assign tmp5403 = s0 ? 1 : tmp3436;
  assign tmp5404 = ~(s0 ? tmp3422 : tmp3457);
  assign tmp5402 = s1 ? tmp5403 : tmp5404;
  assign tmp5406 = s0 ? tmp3460 : tmp5361;
  assign tmp5407 = ~(s0 ? tmp5385 : 0);
  assign tmp5405 = s1 ? tmp5406 : tmp5407;
  assign tmp5401 = ~(s2 ? tmp5402 : tmp5405);
  assign tmp5396 = s3 ? tmp5397 : tmp5401;
  assign tmp5410 = s1 ? 1 : tmp5391;
  assign tmp5411 = ~(s1 ? tmp5400 : 0);
  assign tmp5409 = s2 ? tmp5410 : tmp5411;
  assign tmp5414 = s0 ? 1 : tmp4244;
  assign tmp5415 = s0 ? tmp3460 : tmp5390;
  assign tmp5413 = s1 ? tmp5414 : tmp5415;
  assign tmp5417 = s0 ? tmp5385 : 0;
  assign tmp5418 = s0 ? tmp3422 : 0;
  assign tmp5416 = ~(s1 ? tmp5417 : tmp5418);
  assign tmp5412 = s2 ? tmp5413 : tmp5416;
  assign tmp5408 = ~(s3 ? tmp5409 : tmp5412);
  assign tmp5395 = ~(s4 ? tmp5396 : tmp5408);
  assign tmp5366 = ~(s5 ? tmp5367 : tmp5395);
  assign tmp5344 = s6 ? tmp5345 : tmp5366;
  assign tmp5422 = s1 ? tmp5363 : 0;
  assign tmp5421 = s3 ? tmp5422 : tmp5350;
  assign tmp5426 = s0 ? tmp5363 : 0;
  assign tmp5425 = ~(s1 ? tmp5426 : 0);
  assign tmp5424 = s2 ? tmp5353 : tmp5425;
  assign tmp5423 = ~(s3 ? tmp5424 : tmp5358);
  assign tmp5420 = s4 ? tmp5421 : tmp5423;
  assign tmp5430 = ~(s2 ? tmp5391 : tmp5393);
  assign tmp5429 = ~(s3 ? tmp5382 : tmp5430);
  assign tmp5428 = s4 ? tmp5368 : tmp5429;
  assign tmp5427 = ~(s5 ? tmp5428 : tmp5395);
  assign tmp5419 = s6 ? tmp5420 : tmp5427;
  assign tmp5343 = s8 ? tmp5344 : tmp5419;
  assign tmp5438 = s0 ? tmp3460 : tmp5392;
  assign tmp5437 = s1 ? tmp5414 : tmp5438;
  assign tmp5436 = s2 ? tmp5437 : tmp5416;
  assign tmp5435 = ~(s3 ? tmp5409 : tmp5436);
  assign tmp5434 = ~(s4 ? tmp5396 : tmp5435);
  assign tmp5433 = ~(s5 ? tmp5367 : tmp5434);
  assign tmp5432 = s6 ? tmp5345 : tmp5433;
  assign tmp5431 = s8 ? tmp5419 : tmp5432;
  assign tmp5342 = s9 ? tmp5343 : tmp5431;
  assign tmp5341 = s10 ? tmp5342 : tmp5419;
  assign tmp5233 = s12 ? tmp5234 : tmp5341;
  assign tmp5447 = l1 ? tmp4447 : tmp3597;
  assign tmp5449 = l1 ? tmp5244 : tmp3494;
  assign tmp5448 = ~(s0 ? tmp3459 : tmp5449);
  assign tmp5446 = s1 ? tmp5447 : tmp5448;
  assign tmp5452 = l1 ? tmp4500 : tmp3775;
  assign tmp5453 = ~(l1 ? tmp5249 : tmp3597);
  assign tmp5451 = s0 ? tmp5452 : tmp5453;
  assign tmp5455 = s0 ? tmp5452 : 1;
  assign tmp5454 = s1 ? tmp5455 : tmp5453;
  assign tmp5450 = ~(s2 ? tmp5451 : tmp5454);
  assign tmp5445 = s3 ? tmp5446 : tmp5450;
  assign tmp5459 = s0 ? tmp4944 : 1;
  assign tmp5458 = s1 ? tmp5459 : tmp5453;
  assign tmp5461 = s0 ? tmp5447 : 0;
  assign tmp5460 = ~(s1 ? tmp5461 : tmp4878);
  assign tmp5457 = s2 ? tmp5458 : tmp5460;
  assign tmp5465 = ~(l1 ? tmp3486 : tmp3622);
  assign tmp5464 = s0 ? 1 : tmp5465;
  assign tmp5463 = s1 ? tmp3459 : tmp5464;
  assign tmp5468 = l1 ? tmp5249 : tmp3597;
  assign tmp5469 = l1 ? tmp3422 : tmp3597;
  assign tmp5467 = s0 ? tmp5468 : tmp5469;
  assign tmp5470 = s0 ? tmp4606 : tmp5468;
  assign tmp5466 = ~(s1 ? tmp5467 : tmp5470);
  assign tmp5462 = s2 ? tmp5463 : tmp5466;
  assign tmp5456 = ~(s3 ? tmp5457 : tmp5462);
  assign tmp5444 = s4 ? tmp5445 : tmp5456;
  assign tmp5476 = s0 ? tmp5449 : 1;
  assign tmp5475 = s1 ? tmp5476 : 1;
  assign tmp5478 = s0 ? 1 : tmp5449;
  assign tmp5479 = ~(s0 ? tmp5469 : 0);
  assign tmp5477 = s1 ? tmp5478 : tmp5479;
  assign tmp5474 = s2 ? tmp5475 : tmp5477;
  assign tmp5483 = l1 ? tmp3781 : tmp3775;
  assign tmp5482 = s0 ? 1 : tmp5483;
  assign tmp5485 = ~(l1 ? tmp3422 : tmp3421);
  assign tmp5484 = s0 ? 1 : tmp5485;
  assign tmp5481 = s1 ? tmp5482 : tmp5484;
  assign tmp5487 = s0 ? tmp4606 : tmp4099;
  assign tmp5489 = l1 ? tmp5249 : tmp3421;
  assign tmp5488 = s0 ? tmp5489 : tmp4604;
  assign tmp5486 = ~(s1 ? tmp5487 : tmp5488);
  assign tmp5480 = s2 ? tmp5481 : tmp5486;
  assign tmp5473 = s3 ? tmp5474 : tmp5480;
  assign tmp5493 = s0 ? tmp3665 : tmp5489;
  assign tmp5492 = s1 ? tmp5493 : tmp3495;
  assign tmp5494 = ~(s1 ? tmp3497 : tmp5459);
  assign tmp5491 = s2 ? tmp5492 : tmp5494;
  assign tmp5498 = ~(l1 ? tmp3422 : tmp4418);
  assign tmp5497 = s0 ? tmp4944 : tmp5498;
  assign tmp5499 = s0 ? tmp3460 : tmp5485;
  assign tmp5496 = s1 ? tmp5497 : tmp5499;
  assign tmp5501 = s0 ? tmp3669 : tmp3845;
  assign tmp5500 = ~(s1 ? tmp3845 : tmp5501);
  assign tmp5495 = ~(s2 ? tmp5496 : tmp5500);
  assign tmp5490 = ~(s3 ? tmp5491 : tmp5495);
  assign tmp5472 = s4 ? tmp5473 : tmp5490;
  assign tmp5506 = s0 ? tmp4604 : tmp3460;
  assign tmp5507 = s0 ? tmp3460 : tmp3953;
  assign tmp5505 = s1 ? tmp5506 : tmp5507;
  assign tmp5504 = s2 ? tmp5505 : tmp4681;
  assign tmp5510 = s0 ? tmp3460 : tmp4055;
  assign tmp5509 = s1 ? tmp3497 : tmp5510;
  assign tmp5512 = s0 ? tmp4041 : 1;
  assign tmp5514 = ~(l1 ? 1 : tmp3530);
  assign tmp5513 = s0 ? 1 : tmp5514;
  assign tmp5511 = ~(s1 ? tmp5512 : tmp5513);
  assign tmp5508 = ~(s2 ? tmp5509 : tmp5511);
  assign tmp5503 = s3 ? tmp5504 : tmp5508;
  assign tmp5518 = s0 ? tmp5024 : tmp3796;
  assign tmp5519 = ~(s0 ? tmp3830 : tmp4606);
  assign tmp5517 = s1 ? tmp5518 : tmp5519;
  assign tmp5522 = ~(l1 ? tmp3781 : tmp3494);
  assign tmp5521 = s0 ? tmp3460 : tmp5522;
  assign tmp5520 = ~(s1 ? tmp5521 : 0);
  assign tmp5516 = s2 ? tmp5517 : tmp5520;
  assign tmp5525 = s0 ? tmp3512 : tmp4055;
  assign tmp5526 = ~(s0 ? tmp4041 : tmp4967);
  assign tmp5524 = s1 ? tmp5525 : tmp5526;
  assign tmp5528 = ~(s0 ? tmp3460 : tmp3796);
  assign tmp5527 = ~(s1 ? tmp5513 : tmp5528);
  assign tmp5523 = s2 ? tmp5524 : tmp5527;
  assign tmp5515 = ~(s3 ? tmp5516 : tmp5523);
  assign tmp5502 = ~(s4 ? tmp5503 : tmp5515);
  assign tmp5471 = ~(s5 ? tmp5472 : tmp5502);
  assign tmp5443 = s6 ? tmp5444 : tmp5471;
  assign tmp5534 = l1 ? 1 : tmp3544;
  assign tmp5535 = l1 ? tmp5244 : tmp3420;
  assign tmp5533 = ~(s0 ? tmp5534 : tmp5535);
  assign tmp5532 = s1 ? tmp4659 : tmp5533;
  assign tmp5538 = l1 ? tmp4500 : tmp3420;
  assign tmp5539 = ~(l1 ? tmp5249 : tmp4360);
  assign tmp5537 = s0 ? tmp5538 : tmp5539;
  assign tmp5541 = s0 ? tmp5538 : 1;
  assign tmp5543 = l1 ? tmp5249 : tmp4360;
  assign tmp5544 = l1 ? tmp5249 : tmp3424;
  assign tmp5542 = ~(s0 ? tmp5543 : tmp5544);
  assign tmp5540 = s1 ? tmp5541 : tmp5542;
  assign tmp5536 = ~(s2 ? tmp5537 : tmp5540);
  assign tmp5531 = s3 ? tmp5532 : tmp5536;
  assign tmp5548 = ~(s0 ? tmp5544 : tmp5543);
  assign tmp5547 = s1 ? tmp4595 : tmp5548;
  assign tmp5550 = s0 ? tmp4659 : 0;
  assign tmp5551 = ~(s0 ? tmp4583 : 1);
  assign tmp5549 = ~(s1 ? tmp5550 : tmp5551);
  assign tmp5546 = s2 ? tmp5547 : tmp5549;
  assign tmp5554 = s0 ? tmp4583 : tmp5534;
  assign tmp5553 = s1 ? tmp5554 : tmp5464;
  assign tmp5557 = l1 ? tmp3422 : tmp4360;
  assign tmp5556 = s0 ? tmp5543 : tmp5557;
  assign tmp5559 = l1 ? tmp3422 : tmp4320;
  assign tmp5558 = s0 ? tmp5559 : tmp5543;
  assign tmp5555 = ~(s1 ? tmp5556 : tmp5558);
  assign tmp5552 = s2 ? tmp5553 : tmp5555;
  assign tmp5545 = ~(s3 ? tmp5546 : tmp5552);
  assign tmp5530 = s4 ? tmp5531 : tmp5545;
  assign tmp5565 = s0 ? tmp5535 : 1;
  assign tmp5564 = s1 ? tmp5565 : 1;
  assign tmp5567 = s0 ? 1 : tmp5535;
  assign tmp5568 = ~(s0 ? tmp5557 : 0);
  assign tmp5566 = s1 ? tmp5567 : tmp5568;
  assign tmp5563 = s2 ? tmp5564 : tmp5566;
  assign tmp5572 = l1 ? tmp3781 : tmp3420;
  assign tmp5571 = s0 ? 1 : tmp5572;
  assign tmp5574 = ~(l1 ? tmp3422 : tmp4707);
  assign tmp5573 = s0 ? 1 : tmp5574;
  assign tmp5570 = s1 ? tmp5571 : tmp5573;
  assign tmp5576 = s0 ? tmp5559 : tmp4099;
  assign tmp5578 = l1 ? tmp5249 : tmp4707;
  assign tmp5579 = l1 ? tmp3422 : tmp4707;
  assign tmp5577 = s0 ? tmp5578 : tmp5579;
  assign tmp5575 = ~(s1 ? tmp5576 : tmp5577);
  assign tmp5569 = s2 ? tmp5570 : tmp5575;
  assign tmp5562 = s3 ? tmp5563 : tmp5569;
  assign tmp5584 = l1 ? tmp5249 : tmp4613;
  assign tmp5583 = s0 ? tmp3665 : tmp5584;
  assign tmp5582 = s1 ? tmp5583 : tmp4582;
  assign tmp5586 = s0 ? 1 : tmp4583;
  assign tmp5585 = ~(s1 ? tmp5586 : tmp4595);
  assign tmp5581 = s2 ? tmp5582 : tmp5585;
  assign tmp5590 = ~(l1 ? tmp3422 : tmp4415);
  assign tmp5589 = s0 ? tmp4583 : tmp5590;
  assign tmp5591 = s0 ? tmp4583 : tmp5485;
  assign tmp5588 = s1 ? tmp5589 : tmp5591;
  assign tmp5587 = ~(s2 ? tmp5588 : tmp5500);
  assign tmp5580 = ~(s3 ? tmp5581 : tmp5587);
  assign tmp5561 = s4 ? tmp5562 : tmp5580;
  assign tmp5596 = s0 ? tmp5579 : tmp3460;
  assign tmp5597 = s0 ? tmp3460 : tmp4780;
  assign tmp5595 = s1 ? tmp5596 : tmp5597;
  assign tmp5594 = s2 ? tmp5595 : tmp4781;
  assign tmp5593 = s3 ? tmp5594 : tmp5508;
  assign tmp5601 = ~(s0 ? tmp3830 : tmp5559);
  assign tmp5600 = s1 ? tmp5518 : tmp5601;
  assign tmp5604 = ~(l1 ? tmp3781 : tmp3420);
  assign tmp5603 = s0 ? tmp3460 : tmp5604;
  assign tmp5602 = ~(s1 ? tmp5603 : 0);
  assign tmp5599 = s2 ? tmp5600 : tmp5602;
  assign tmp5607 = s0 ? tmp4783 : tmp4055;
  assign tmp5606 = s1 ? tmp5607 : tmp5526;
  assign tmp5605 = s2 ? tmp5606 : tmp5527;
  assign tmp5598 = ~(s3 ? tmp5599 : tmp5605);
  assign tmp5592 = ~(s4 ? tmp5593 : tmp5598);
  assign tmp5560 = ~(s5 ? tmp5561 : tmp5592);
  assign tmp5529 = s6 ? tmp5530 : tmp5560;
  assign tmp5442 = s8 ? tmp5443 : tmp5529;
  assign tmp5613 = l1 ? tmp4447 : tmp3783;
  assign tmp5615 = l1 ? tmp5244 : tmp3863;
  assign tmp5614 = ~(s0 ? tmp5534 : tmp5615);
  assign tmp5612 = s1 ? tmp5613 : tmp5614;
  assign tmp5618 = l1 ? tmp4500 : tmp3544;
  assign tmp5619 = ~(l1 ? tmp5249 : tmp4286);
  assign tmp5617 = s0 ? tmp5618 : tmp5619;
  assign tmp5621 = s0 ? tmp5618 : 1;
  assign tmp5623 = l1 ? tmp5249 : tmp4286;
  assign tmp5624 = l1 ? tmp5249 : tmp3783;
  assign tmp5622 = ~(s0 ? tmp5623 : tmp5624);
  assign tmp5620 = s1 ? tmp5621 : tmp5622;
  assign tmp5616 = ~(s2 ? tmp5617 : tmp5620);
  assign tmp5611 = s3 ? tmp5612 : tmp5616;
  assign tmp5629 = l1 ? 1 : tmp3863;
  assign tmp5628 = s0 ? tmp5629 : 1;
  assign tmp5630 = ~(s0 ? tmp5624 : tmp5623);
  assign tmp5627 = s1 ? tmp5628 : tmp5630;
  assign tmp5632 = s0 ? tmp5613 : 0;
  assign tmp5631 = ~(s1 ? tmp5632 : tmp5551);
  assign tmp5626 = s2 ? tmp5627 : tmp5631;
  assign tmp5636 = l1 ? tmp3422 : tmp4286;
  assign tmp5635 = s0 ? tmp5623 : tmp5636;
  assign tmp5637 = s0 ? tmp5559 : tmp5623;
  assign tmp5634 = ~(s1 ? tmp5635 : tmp5637);
  assign tmp5633 = s2 ? tmp5553 : tmp5634;
  assign tmp5625 = ~(s3 ? tmp5626 : tmp5633);
  assign tmp5610 = s4 ? tmp5611 : tmp5625;
  assign tmp5643 = s0 ? tmp5615 : 1;
  assign tmp5642 = s1 ? tmp5643 : 1;
  assign tmp5646 = l1 ? tmp5244 : tmp3822;
  assign tmp5645 = s0 ? 1 : tmp5646;
  assign tmp5647 = ~(s0 ? tmp5636 : 0);
  assign tmp5644 = s1 ? tmp5645 : tmp5647;
  assign tmp5641 = s2 ? tmp5642 : tmp5644;
  assign tmp5651 = l1 ? tmp3781 : tmp3544;
  assign tmp5650 = s0 ? 1 : tmp5651;
  assign tmp5653 = ~(l1 ? tmp3422 : tmp4320);
  assign tmp5652 = s0 ? 1 : tmp5653;
  assign tmp5649 = s1 ? tmp5650 : tmp5652;
  assign tmp5656 = l1 ? tmp5249 : tmp4320;
  assign tmp5655 = s0 ? tmp5656 : tmp5559;
  assign tmp5654 = ~(s1 ? tmp5576 : tmp5655);
  assign tmp5648 = s2 ? tmp5649 : tmp5654;
  assign tmp5640 = s3 ? tmp5641 : tmp5648;
  assign tmp5661 = l1 ? tmp5249 : tmp4275;
  assign tmp5660 = s0 ? tmp3665 : tmp5661;
  assign tmp5659 = s1 ? tmp5660 : tmp4582;
  assign tmp5664 = l1 ? 1 : tmp3822;
  assign tmp5663 = s0 ? tmp5664 : 1;
  assign tmp5662 = ~(s1 ? tmp5586 : tmp5663);
  assign tmp5658 = s2 ? tmp5659 : tmp5662;
  assign tmp5668 = ~(l1 ? tmp3422 : tmp4275);
  assign tmp5667 = s0 ? tmp5664 : tmp5668;
  assign tmp5670 = ~(l1 ? tmp3422 : tmp3622);
  assign tmp5669 = s0 ? tmp4583 : tmp5670;
  assign tmp5666 = s1 ? tmp5667 : tmp5669;
  assign tmp5665 = ~(s2 ? tmp5666 : tmp5500);
  assign tmp5657 = ~(s3 ? tmp5658 : tmp5665);
  assign tmp5639 = s4 ? tmp5640 : tmp5657;
  assign tmp5675 = s0 ? tmp5559 : tmp3460;
  assign tmp5674 = s1 ? tmp5675 : tmp5597;
  assign tmp5673 = s2 ? tmp5674 : tmp4781;
  assign tmp5677 = ~(s1 ? tmp5512 : tmp4870);
  assign tmp5676 = ~(s2 ? tmp5509 : tmp5677);
  assign tmp5672 = s3 ? tmp5673 : tmp5676;
  assign tmp5681 = s0 ? tmp3460 : tmp3796;
  assign tmp5680 = s1 ? tmp5681 : tmp5601;
  assign tmp5684 = ~(l1 ? tmp3781 : tmp3822);
  assign tmp5683 = s0 ? tmp3460 : tmp5684;
  assign tmp5682 = ~(s1 ? tmp5683 : 0);
  assign tmp5679 = s2 ? tmp5680 : tmp5682;
  assign tmp5687 = ~(s0 ? tmp4041 : tmp3830);
  assign tmp5686 = s1 ? tmp5607 : tmp5687;
  assign tmp5688 = ~(s1 ? tmp4870 : tmp5528);
  assign tmp5685 = s2 ? tmp5686 : tmp5688;
  assign tmp5678 = ~(s3 ? tmp5679 : tmp5685);
  assign tmp5671 = ~(s4 ? tmp5672 : tmp5678);
  assign tmp5638 = ~(s5 ? tmp5639 : tmp5671);
  assign tmp5609 = s6 ? tmp5610 : tmp5638;
  assign tmp5608 = s8 ? tmp5529 : tmp5609;
  assign tmp5441 = s9 ? tmp5442 : tmp5608;
  assign tmp5440 = s10 ? tmp5441 : tmp5529;
  assign tmp5696 = l1 ? tmp4500 : tmp5244;
  assign tmp5697 = s0 ? 1 : tmp5252;
  assign tmp5695 = s1 ? tmp5696 : tmp5697;
  assign tmp5701 = l1 ? tmp4500 : tmp3538;
  assign tmp5700 = s0 ? 1 : tmp5701;
  assign tmp5702 = s0 ? tmp5252 : tmp5701;
  assign tmp5699 = s1 ? tmp5700 : tmp5702;
  assign tmp5703 = s1 ? tmp5254 : tmp5701;
  assign tmp5698 = s2 ? tmp5699 : tmp5703;
  assign tmp5694 = s3 ? tmp5695 : tmp5698;
  assign tmp5706 = s1 ? 1 : tmp5701;
  assign tmp5708 = s0 ? tmp5696 : 1;
  assign tmp5707 = s1 ? tmp5708 : 1;
  assign tmp5705 = s2 ? tmp5706 : tmp5707;
  assign tmp5710 = s1 ? 1 : tmp3694;
  assign tmp5713 = l1 ? tmp4608 : tmp3538;
  assign tmp5712 = s0 ? tmp5701 : tmp5713;
  assign tmp5714 = s0 ? tmp3646 : tmp5701;
  assign tmp5711 = s1 ? tmp5712 : tmp5714;
  assign tmp5709 = s2 ? tmp5710 : tmp5711;
  assign tmp5704 = s3 ? tmp5705 : tmp5709;
  assign tmp5693 = s4 ? tmp5694 : tmp5704;
  assign tmp5719 = s1 ? tmp5254 : 1;
  assign tmp5721 = s0 ? tmp5713 : 1;
  assign tmp5720 = s1 ? tmp5697 : tmp5721;
  assign tmp5718 = s2 ? tmp5719 : tmp5720;
  assign tmp5726 = l2 ? tmp3538 : tmp3436;
  assign tmp5725 = l1 ? tmp4608 : tmp5726;
  assign tmp5724 = s0 ? 1 : tmp5725;
  assign tmp5723 = s1 ? tmp5281 : tmp5724;
  assign tmp5728 = s0 ? tmp3646 : tmp3512;
  assign tmp5730 = l1 ? tmp4500 : tmp5726;
  assign tmp5731 = l1 ? tmp4608 : tmp3436;
  assign tmp5729 = s0 ? tmp5730 : tmp5731;
  assign tmp5727 = s1 ? tmp5728 : tmp5729;
  assign tmp5722 = s2 ? tmp5723 : tmp5727;
  assign tmp5717 = s3 ? tmp5718 : tmp5722;
  assign tmp5736 = l1 ? tmp4500 : tmp3781;
  assign tmp5735 = s0 ? tmp3646 : tmp5736;
  assign tmp5734 = s1 ? tmp5735 : 1;
  assign tmp5733 = s2 ? tmp5734 : 1;
  assign tmp5739 = s0 ? 1 : tmp3781;
  assign tmp5740 = s0 ? 1 : tmp5731;
  assign tmp5738 = s1 ? tmp5739 : tmp5740;
  assign tmp5742 = s0 ? tmp3646 : tmp3460;
  assign tmp5741 = s1 ? tmp3460 : tmp5742;
  assign tmp5737 = s2 ? tmp5738 : tmp5741;
  assign tmp5732 = s3 ? tmp5733 : tmp5737;
  assign tmp5716 = s4 ? tmp5717 : tmp5732;
  assign tmp5747 = s0 ? tmp5725 : tmp3512;
  assign tmp5746 = s1 ? tmp5747 : tmp4482;
  assign tmp5745 = s2 ? tmp5746 : tmp3697;
  assign tmp5751 = ~(l1 ? 1 : tmp3422);
  assign tmp5750 = s0 ? 1 : tmp5751;
  assign tmp5749 = s1 ? tmp5750 : tmp4878;
  assign tmp5754 = ~(l1 ? tmp3434 : tmp3436);
  assign tmp5753 = s0 ? 1 : tmp5754;
  assign tmp5755 = ~(s0 ? tmp3646 : 1);
  assign tmp5752 = ~(s1 ? tmp5753 : tmp5755);
  assign tmp5748 = s2 ? tmp5749 : tmp5752;
  assign tmp5744 = s3 ? tmp5745 : tmp5748;
  assign tmp5759 = s0 ? tmp3644 : tmp3646;
  assign tmp5758 = s1 ? tmp3700 : tmp5759;
  assign tmp5762 = l1 ? tmp4608 : 1;
  assign tmp5761 = s0 ? tmp3512 : tmp5762;
  assign tmp5760 = s1 ? tmp5761 : 1;
  assign tmp5757 = s2 ? tmp5758 : tmp5760;
  assign tmp5766 = l1 ? tmp3434 : tmp3782;
  assign tmp5765 = s0 ? tmp3434 : tmp5766;
  assign tmp5768 = ~(l1 ? tmp4608 : tmp3781);
  assign tmp5767 = ~(s0 ? 1 : tmp5768);
  assign tmp5764 = s1 ? tmp5765 : tmp5767;
  assign tmp5770 = s0 ? tmp3646 : 1;
  assign tmp5771 = ~(s0 ? tmp3459 : tmp5335);
  assign tmp5769 = s1 ? tmp5770 : tmp5771;
  assign tmp5763 = s2 ? tmp5764 : tmp5769;
  assign tmp5756 = s3 ? tmp5757 : tmp5763;
  assign tmp5743 = s4 ? tmp5744 : tmp5756;
  assign tmp5715 = s5 ? tmp5716 : tmp5743;
  assign tmp5692 = s6 ? tmp5693 : tmp5715;
  assign tmp5775 = s1 ? tmp5701 : tmp5697;
  assign tmp5774 = s3 ? tmp5775 : tmp5698;
  assign tmp5779 = s0 ? tmp5701 : 1;
  assign tmp5778 = s1 ? tmp5779 : 1;
  assign tmp5777 = s2 ? tmp5706 : tmp5778;
  assign tmp5776 = s3 ? tmp5777 : tmp5709;
  assign tmp5773 = s4 ? tmp5774 : tmp5776;
  assign tmp5785 = s0 ? 1 : tmp3795;
  assign tmp5784 = s1 ? tmp5785 : tmp5740;
  assign tmp5783 = s2 ? tmp5784 : tmp5741;
  assign tmp5782 = s3 ? tmp5733 : tmp5783;
  assign tmp5781 = s4 ? tmp5717 : tmp5782;
  assign tmp5789 = s1 ? tmp5747 : tmp3679;
  assign tmp5788 = s2 ? tmp5789 : tmp3703;
  assign tmp5787 = s3 ? tmp5788 : tmp5748;
  assign tmp5793 = s0 ? tmp3644 : tmp5766;
  assign tmp5792 = s1 ? tmp5793 : tmp5767;
  assign tmp5791 = s2 ? tmp5792 : tmp5769;
  assign tmp5790 = s3 ? tmp5757 : tmp5791;
  assign tmp5786 = s4 ? tmp5787 : tmp5790;
  assign tmp5780 = s5 ? tmp5781 : tmp5786;
  assign tmp5772 = s6 ? tmp5773 : tmp5780;
  assign tmp5691 = s8 ? tmp5692 : tmp5772;
  assign tmp5802 = ~(l1 ? tmp4608 : tmp3436);
  assign tmp5801 = ~(s0 ? 1 : tmp5802);
  assign tmp5800 = s1 ? tmp5793 : tmp5801;
  assign tmp5799 = s2 ? tmp5800 : tmp5769;
  assign tmp5798 = s3 ? tmp5757 : tmp5799;
  assign tmp5797 = s4 ? tmp5787 : tmp5798;
  assign tmp5796 = s5 ? tmp5716 : tmp5797;
  assign tmp5795 = s6 ? tmp5693 : tmp5796;
  assign tmp5794 = s8 ? tmp5772 : tmp5795;
  assign tmp5690 = s9 ? tmp5691 : tmp5794;
  assign tmp5689 = ~(s10 ? tmp5690 : tmp5772);
  assign tmp5439 = s12 ? tmp5440 : tmp5689;
  assign tmp5232 = s13 ? tmp5233 : tmp5439;
  assign tmp5812 = s0 ? tmp3422 : tmp5802;
  assign tmp5811 = s1 ? tmp3422 : tmp5812;
  assign tmp5815 = ~(l1 ? tmp4414 : tmp3422);
  assign tmp5814 = s0 ? tmp3795 : tmp5815;
  assign tmp5817 = s0 ? tmp3795 : 0;
  assign tmp5816 = s1 ? tmp5817 : tmp5815;
  assign tmp5813 = ~(s2 ? tmp5814 : tmp5816);
  assign tmp5810 = s3 ? tmp5811 : tmp5813;
  assign tmp5820 = s1 ? tmp3795 : tmp5815;
  assign tmp5819 = s2 ? tmp5820 : tmp3800;
  assign tmp5822 = s1 ? tmp3422 : tmp4867;
  assign tmp5825 = l1 ? tmp4414 : tmp3422;
  assign tmp5826 = l1 ? tmp4447 : tmp3422;
  assign tmp5824 = s0 ? tmp5825 : tmp5826;
  assign tmp5828 = l1 ? tmp3775 : tmp3422;
  assign tmp5827 = s0 ? tmp5828 : tmp5825;
  assign tmp5823 = s1 ? tmp5824 : tmp5827;
  assign tmp5821 = ~(s2 ? tmp5822 : tmp5823);
  assign tmp5818 = ~(s3 ? tmp5819 : tmp5821);
  assign tmp5809 = s4 ? tmp5810 : tmp5818;
  assign tmp5834 = s0 ? tmp5731 : 0;
  assign tmp5833 = s1 ? tmp5834 : tmp3795;
  assign tmp5837 = ~(l1 ? tmp4608 : tmp3622);
  assign tmp5836 = s0 ? 1 : tmp5837;
  assign tmp5838 = s0 ? tmp5826 : 1;
  assign tmp5835 = ~(s1 ? tmp5836 : tmp5838);
  assign tmp5832 = s2 ? tmp5833 : tmp5835;
  assign tmp5841 = s0 ? 1 : tmp4017;
  assign tmp5842 = s0 ? 1 : tmp5826;
  assign tmp5840 = s1 ? tmp5841 : tmp5842;
  assign tmp5843 = s1 ? tmp5828 : tmp5824;
  assign tmp5839 = ~(s2 ? tmp5840 : tmp5843);
  assign tmp5831 = s3 ? tmp5832 : tmp5839;
  assign tmp5847 = s0 ? tmp3422 : tmp5825;
  assign tmp5846 = s1 ? tmp5847 : tmp3832;
  assign tmp5849 = ~(l1 ? tmp3781 : tmp3622);
  assign tmp5848 = s1 ? tmp3832 : tmp5849;
  assign tmp5845 = s2 ? tmp5846 : tmp5848;
  assign tmp5853 = ~(l1 ? tmp3422 : tmp3435);
  assign tmp5852 = s0 ? tmp3665 : tmp5853;
  assign tmp5855 = ~(l1 ? tmp4447 : tmp3422);
  assign tmp5854 = s0 ? 1 : tmp5855;
  assign tmp5851 = s1 ? tmp5852 : tmp5854;
  assign tmp5857 = s0 ? tmp3459 : 1;
  assign tmp5856 = ~(s1 ? 1 : tmp5857);
  assign tmp5850 = ~(s2 ? tmp5851 : tmp5856);
  assign tmp5844 = ~(s3 ? tmp5845 : tmp5850);
  assign tmp5830 = s4 ? tmp5831 : tmp5844;
  assign tmp5861 = s1 ? tmp5838 : tmp5334;
  assign tmp5863 = s0 ? tmp3644 : tmp3845;
  assign tmp5862 = ~(s1 ? tmp5863 : tmp3844);
  assign tmp5860 = s2 ? tmp5861 : tmp5862;
  assign tmp5867 = l1 ? 1 : tmp3435;
  assign tmp5866 = s0 ? 1 : tmp5867;
  assign tmp5868 = s0 ? tmp5867 : 0;
  assign tmp5865 = ~(s1 ? tmp5866 : tmp5868);
  assign tmp5864 = ~(s2 ? tmp5749 : tmp5865);
  assign tmp5859 = s3 ? tmp5860 : tmp5864;
  assign tmp5873 = ~(l1 ? tmp3775 : tmp3422);
  assign tmp5872 = s0 ? tmp3644 : tmp5873;
  assign tmp5871 = s1 ? tmp3700 : tmp5872;
  assign tmp5876 = ~(l1 ? tmp4500 : tmp3622);
  assign tmp5875 = s0 ? 1 : tmp5876;
  assign tmp5874 = ~(s1 ? tmp5875 : tmp5037);
  assign tmp5870 = s2 ? tmp5871 : tmp5874;
  assign tmp5880 = l1 ? tmp4447 : tmp3435;
  assign tmp5879 = ~(s0 ? 1 : tmp5880);
  assign tmp5878 = s1 ? tmp5759 : tmp5879;
  assign tmp5882 = s0 ? tmp3459 : tmp5335;
  assign tmp5881 = ~(s1 ? tmp5868 : tmp5882);
  assign tmp5877 = s2 ? tmp5878 : tmp5881;
  assign tmp5869 = ~(s3 ? tmp5870 : tmp5877);
  assign tmp5858 = ~(s4 ? tmp5859 : tmp5869);
  assign tmp5829 = ~(s5 ? tmp5830 : tmp5858);
  assign tmp5808 = s6 ? tmp5809 : tmp5829;
  assign tmp5887 = l1 ? tmp4706 : tmp3422;
  assign tmp5889 = l1 ? tmp4507 : tmp3422;
  assign tmp5888 = s0 ? tmp3878 : tmp5889;
  assign tmp5886 = s1 ? tmp5887 : tmp5888;
  assign tmp5892 = l1 ? tmp4515 : tmp3422;
  assign tmp5891 = s0 ? tmp3862 : tmp5892;
  assign tmp5894 = s0 ? tmp3862 : tmp3459;
  assign tmp5893 = s1 ? tmp5894 : tmp5892;
  assign tmp5890 = s2 ? tmp5891 : tmp5893;
  assign tmp5885 = s3 ? tmp5886 : tmp5890;
  assign tmp5897 = s1 ? tmp3862 : tmp5892;
  assign tmp5899 = s0 ? tmp5887 : 1;
  assign tmp5898 = s1 ? tmp5899 : tmp3877;
  assign tmp5896 = s2 ? tmp5897 : tmp5898;
  assign tmp5901 = s1 ? tmp3878 : tmp4867;
  assign tmp5904 = l1 ? tmp4561 : tmp3422;
  assign tmp5903 = s0 ? tmp5892 : tmp5904;
  assign tmp5905 = s0 ? tmp5828 : tmp5892;
  assign tmp5902 = s1 ? tmp5903 : tmp5905;
  assign tmp5900 = s2 ? tmp5901 : tmp5902;
  assign tmp5895 = s3 ? tmp5896 : tmp5900;
  assign tmp5884 = s4 ? tmp5885 : tmp5895;
  assign tmp5911 = s0 ? tmp5889 : 1;
  assign tmp5910 = s1 ? tmp5911 : tmp3890;
  assign tmp5914 = l1 ? tmp4507 : tmp3427;
  assign tmp5913 = s0 ? 1 : tmp5914;
  assign tmp5915 = s0 ? tmp5904 : tmp3459;
  assign tmp5912 = s1 ? tmp5913 : tmp5915;
  assign tmp5909 = s2 ? tmp5910 : tmp5912;
  assign tmp5918 = s0 ? tmp3459 : tmp3862;
  assign tmp5919 = s0 ? tmp3459 : tmp5826;
  assign tmp5917 = s1 ? tmp5918 : tmp5919;
  assign tmp5920 = s1 ? tmp5828 : tmp5903;
  assign tmp5916 = s2 ? tmp5917 : tmp5920;
  assign tmp5908 = s3 ? tmp5909 : tmp5916;
  assign tmp5924 = s0 ? tmp3422 : tmp5892;
  assign tmp5923 = s1 ? tmp5924 : tmp3909;
  assign tmp5926 = l1 ? tmp3863 : tmp3427;
  assign tmp5925 = s1 ? tmp3909 : tmp5926;
  assign tmp5922 = s2 ? tmp5923 : tmp5925;
  assign tmp5930 = ~(l1 ? tmp4706 : tmp3435);
  assign tmp5929 = s0 ? tmp3665 : tmp5930;
  assign tmp5931 = ~(s0 ? tmp3512 : tmp5826);
  assign tmp5928 = s1 ? tmp5929 : tmp5931;
  assign tmp5927 = ~(s2 ? tmp5928 : tmp5856);
  assign tmp5921 = s3 ? tmp5922 : tmp5927;
  assign tmp5907 = s4 ? tmp5908 : tmp5921;
  assign tmp5936 = s0 ? tmp3644 : tmp3665;
  assign tmp5935 = ~(s1 ? tmp5936 : tmp3849);
  assign tmp5934 = s2 ? tmp5861 : tmp5935;
  assign tmp5933 = s3 ? tmp5934 : tmp5864;
  assign tmp5939 = ~(s1 ? tmp5875 : tmp5116);
  assign tmp5938 = s2 ? tmp5871 : tmp5939;
  assign tmp5937 = ~(s3 ? tmp5938 : tmp5877);
  assign tmp5932 = s4 ? tmp5933 : tmp5937;
  assign tmp5906 = s5 ? tmp5907 : tmp5932;
  assign tmp5883 = s6 ? tmp5884 : tmp5906;
  assign tmp5807 = s8 ? tmp5808 : tmp5883;
  assign tmp5945 = l1 ? tmp4706 : tmp3863;
  assign tmp5947 = l1 ? tmp4507 : tmp3863;
  assign tmp5946 = s0 ? tmp4509 : tmp5947;
  assign tmp5944 = s1 ? tmp5945 : tmp5946;
  assign tmp5951 = l1 ? tmp4515 : tmp4706;
  assign tmp5950 = s0 ? tmp5127 : tmp5951;
  assign tmp5953 = l1 ? tmp3863 : tmp3544;
  assign tmp5952 = s0 ? tmp5953 : tmp5951;
  assign tmp5949 = s1 ? tmp5950 : tmp5952;
  assign tmp5955 = s0 ? tmp5953 : 1;
  assign tmp5957 = l1 ? tmp4515 : tmp3863;
  assign tmp5956 = s0 ? tmp5951 : tmp5957;
  assign tmp5954 = s1 ? tmp5955 : tmp5956;
  assign tmp5948 = s2 ? tmp5949 : tmp5954;
  assign tmp5943 = s3 ? tmp5944 : tmp5948;
  assign tmp5961 = s0 ? tmp3863 : tmp3685;
  assign tmp5962 = s0 ? tmp5957 : tmp5951;
  assign tmp5960 = s1 ? tmp5961 : tmp5962;
  assign tmp5964 = s0 ? tmp5945 : 1;
  assign tmp5963 = s1 ? tmp5964 : tmp4528;
  assign tmp5959 = s2 ? tmp5960 : tmp5963;
  assign tmp5966 = s1 ? tmp4532 : tmp4867;
  assign tmp5969 = l1 ? tmp4561 : tmp4706;
  assign tmp5968 = s0 ? tmp5951 : tmp5969;
  assign tmp5971 = l1 ? tmp3775 : tmp4706;
  assign tmp5970 = s0 ? tmp5971 : tmp5951;
  assign tmp5967 = s1 ? tmp5968 : tmp5970;
  assign tmp5965 = s2 ? tmp5966 : tmp5967;
  assign tmp5958 = s3 ? tmp5959 : tmp5965;
  assign tmp5942 = s4 ? tmp5943 : tmp5958;
  assign tmp5977 = s0 ? tmp5947 : 1;
  assign tmp5976 = s1 ? tmp5977 : tmp5149;
  assign tmp5980 = l1 ? tmp4507 : tmp3822;
  assign tmp5979 = s0 ? 1 : tmp5980;
  assign tmp5981 = s0 ? tmp5969 : 1;
  assign tmp5978 = s1 ? tmp5979 : tmp5981;
  assign tmp5975 = s2 ? tmp5976 : tmp5978;
  assign tmp5984 = s0 ? 1 : tmp5953;
  assign tmp5986 = l1 ? tmp4447 : tmp4706;
  assign tmp5985 = s0 ? 1 : tmp5986;
  assign tmp5983 = s1 ? tmp5984 : tmp5985;
  assign tmp5988 = s0 ? tmp5971 : 1;
  assign tmp5987 = s1 ? tmp5988 : tmp5968;
  assign tmp5982 = s2 ? tmp5983 : tmp5987;
  assign tmp5974 = s3 ? tmp5975 : tmp5982;
  assign tmp5992 = s0 ? tmp3422 : tmp5957;
  assign tmp5991 = s1 ? tmp5992 : tmp4567;
  assign tmp5995 = l1 ? tmp3863 : tmp3822;
  assign tmp5994 = s0 ? tmp5995 : tmp3685;
  assign tmp5993 = s1 ? tmp4567 : tmp5994;
  assign tmp5990 = s2 ? tmp5991 : tmp5993;
  assign tmp5999 = ~(l1 ? tmp4706 : tmp3863);
  assign tmp5998 = s0 ? tmp4274 : tmp5999;
  assign tmp6000 = ~(s0 ? tmp3822 : tmp5826);
  assign tmp5997 = s1 ? tmp5998 : tmp6000;
  assign tmp5996 = ~(s2 ? tmp5997 : tmp5856);
  assign tmp5989 = s3 ? tmp5990 : tmp5996;
  assign tmp5973 = s4 ? tmp5974 : tmp5989;
  assign tmp6005 = s0 ? tmp5986 : 1;
  assign tmp6007 = ~(l1 ? tmp3434 : tmp3424);
  assign tmp6006 = s0 ? 1 : tmp6007;
  assign tmp6004 = s1 ? tmp6005 : tmp6006;
  assign tmp6009 = s0 ? tmp3518 : tmp3460;
  assign tmp6008 = ~(s1 ? tmp6009 : tmp3497);
  assign tmp6003 = s2 ? tmp6004 : tmp6008;
  assign tmp6002 = s3 ? tmp6003 : tmp5864;
  assign tmp6014 = ~(l1 ? tmp3775 : tmp4706);
  assign tmp6013 = s0 ? tmp3644 : tmp6014;
  assign tmp6012 = s1 ? tmp3700 : tmp6013;
  assign tmp6017 = ~(l1 ? tmp4500 : tmp4275);
  assign tmp6016 = s0 ? 1 : tmp6017;
  assign tmp6015 = ~(s1 ? tmp6016 : tmp5178);
  assign tmp6011 = s2 ? tmp6012 : tmp6015;
  assign tmp6020 = s0 ? tmp3518 : tmp3646;
  assign tmp6019 = s1 ? tmp6020 : tmp5879;
  assign tmp6018 = s2 ? tmp6019 : tmp5881;
  assign tmp6010 = ~(s3 ? tmp6011 : tmp6018);
  assign tmp6001 = s4 ? tmp6002 : tmp6010;
  assign tmp5972 = s5 ? tmp5973 : tmp6001;
  assign tmp5941 = s6 ? tmp5942 : tmp5972;
  assign tmp5940 = s8 ? tmp5883 : tmp5941;
  assign tmp5806 = s9 ? tmp5807 : tmp5940;
  assign tmp6026 = s0 ? tmp5188 : tmp5951;
  assign tmp6027 = s0 ? tmp3863 : tmp5951;
  assign tmp6025 = s1 ? tmp6026 : tmp6027;
  assign tmp6029 = s0 ? tmp3863 : 1;
  assign tmp6028 = s1 ? tmp6029 : tmp5956;
  assign tmp6024 = s2 ? tmp6025 : tmp6028;
  assign tmp6023 = s3 ? tmp5944 : tmp6024;
  assign tmp6022 = s4 ? tmp6023 : tmp5958;
  assign tmp6034 = s1 ? tmp5977 : tmp5210;
  assign tmp6033 = s2 ? tmp6034 : tmp5978;
  assign tmp6037 = s0 ? 1 : tmp3863;
  assign tmp6036 = s1 ? tmp6037 : tmp5985;
  assign tmp6035 = s2 ? tmp6036 : tmp5987;
  assign tmp6032 = s3 ? tmp6033 : tmp6035;
  assign tmp6031 = s4 ? tmp6032 : tmp5989;
  assign tmp6042 = s0 ? tmp3518 : tmp3845;
  assign tmp6041 = ~(s1 ? tmp6042 : tmp3844);
  assign tmp6040 = s2 ? tmp6004 : tmp6041;
  assign tmp6039 = s3 ? tmp6040 : tmp5864;
  assign tmp6045 = ~(s1 ? tmp6016 : tmp5037);
  assign tmp6044 = s2 ? tmp6012 : tmp6045;
  assign tmp6043 = ~(s3 ? tmp6044 : tmp6018);
  assign tmp6038 = s4 ? tmp6039 : tmp6043;
  assign tmp6030 = s5 ? tmp6031 : tmp6038;
  assign tmp6021 = s6 ? tmp6022 : tmp6030;
  assign tmp5805 = s10 ? tmp5806 : tmp6021;
  assign tmp6053 = l1 ? tmp3494 : tmp4414;
  assign tmp6055 = ~(l1 ? tmp3418 : tmp4435);
  assign tmp6054 = s0 ? tmp3459 : tmp6055;
  assign tmp6052 = s1 ? tmp6053 : tmp6054;
  assign tmp6058 = l1 ? tmp3429 : tmp3436;
  assign tmp6060 = l2 ? tmp3422 : tmp3538;
  assign tmp6059 = ~(l1 ? tmp6060 : tmp4414);
  assign tmp6057 = s0 ? tmp6058 : tmp6059;
  assign tmp6062 = s0 ? tmp6058 : 0;
  assign tmp6061 = s1 ? tmp6062 : tmp6059;
  assign tmp6056 = ~(s2 ? tmp6057 : tmp6061);
  assign tmp6051 = s3 ? tmp6052 : tmp6056;
  assign tmp6067 = l1 ? tmp3434 : tmp4435;
  assign tmp6066 = s0 ? tmp6067 : 0;
  assign tmp6065 = s1 ? tmp6066 : tmp6059;
  assign tmp6069 = s0 ? tmp6053 : 1;
  assign tmp6068 = ~(s1 ? tmp6069 : tmp5857);
  assign tmp6064 = s2 ? tmp6065 : tmp6068;
  assign tmp6071 = s1 ? tmp3459 : tmp5482;
  assign tmp6074 = l1 ? tmp6060 : tmp4414;
  assign tmp6075 = l1 ? tmp3545 : tmp4414;
  assign tmp6073 = s0 ? tmp6074 : tmp6075;
  assign tmp6077 = l1 ? tmp3545 : tmp3775;
  assign tmp6076 = s0 ? tmp6077 : tmp6074;
  assign tmp6072 = s1 ? tmp6073 : tmp6076;
  assign tmp6070 = ~(s2 ? tmp6071 : tmp6072);
  assign tmp6063 = ~(s3 ? tmp6064 : tmp6070);
  assign tmp6050 = s4 ? tmp6051 : tmp6063;
  assign tmp6084 = l1 ? tmp3418 : tmp4435;
  assign tmp6083 = s0 ? tmp6084 : 0;
  assign tmp6085 = ~(s0 ? 1 : tmp5754);
  assign tmp6082 = s1 ? tmp6083 : tmp6085;
  assign tmp6088 = ~(l1 ? tmp3418 : tmp4454);
  assign tmp6087 = s0 ? 1 : tmp6088;
  assign tmp6089 = s0 ? tmp6075 : 1;
  assign tmp6086 = ~(s1 ? tmp6087 : tmp6089);
  assign tmp6081 = s2 ? tmp6082 : tmp6086;
  assign tmp6093 = ~(l1 ? tmp3486 : tmp3436);
  assign tmp6092 = s0 ? 1 : tmp6093;
  assign tmp6095 = l1 ? tmp3545 : tmp4447;
  assign tmp6094 = s0 ? 1 : tmp6095;
  assign tmp6091 = s1 ? tmp6092 : tmp6094;
  assign tmp6097 = s0 ? tmp6077 : tmp4090;
  assign tmp6099 = l1 ? tmp6060 : tmp4447;
  assign tmp6098 = s0 ? tmp6099 : tmp6095;
  assign tmp6096 = s1 ? tmp6097 : tmp6098;
  assign tmp6090 = ~(s2 ? tmp6091 : tmp6096);
  assign tmp6080 = s3 ? tmp6081 : tmp6090;
  assign tmp6104 = l1 ? tmp3434 : tmp3775;
  assign tmp6103 = s0 ? tmp6104 : tmp6099;
  assign tmp6102 = s1 ? tmp6103 : tmp3497;
  assign tmp6107 = l1 ? tmp3434 : tmp4454;
  assign tmp6106 = ~(s0 ? tmp6107 : 0);
  assign tmp6105 = s1 ? tmp3497 : tmp6106;
  assign tmp6101 = s2 ? tmp6102 : tmp6105;
  assign tmp6111 = ~(l1 ? tmp3545 : tmp4470);
  assign tmp6110 = s0 ? tmp6107 : tmp6111;
  assign tmp6112 = ~(s0 ? tmp3460 : tmp6095);
  assign tmp6109 = s1 ? tmp6110 : tmp6112;
  assign tmp6114 = s0 ? tmp5483 : 1;
  assign tmp6113 = ~(s1 ? 1 : tmp6114);
  assign tmp6108 = ~(s2 ? tmp6109 : tmp6113);
  assign tmp6100 = ~(s3 ? tmp6101 : tmp6108);
  assign tmp6079 = s4 ? tmp6080 : tmp6100;
  assign tmp6119 = s0 ? tmp6095 : tmp3434;
  assign tmp6120 = s0 ? tmp3434 : 0;
  assign tmp6118 = s1 ? tmp6119 : tmp6120;
  assign tmp6122 = s0 ? 1 : tmp3639;
  assign tmp6123 = s0 ? tmp3644 : tmp3639;
  assign tmp6121 = ~(s1 ? tmp6122 : tmp6123);
  assign tmp6117 = s2 ? tmp6118 : tmp6121;
  assign tmp6125 = s1 ? tmp5400 : tmp5327;
  assign tmp6128 = ~(l1 ? tmp3434 : tmp3640);
  assign tmp6127 = s0 ? tmp4059 : tmp6128;
  assign tmp6130 = ~(l1 ? tmp3434 : tmp4500);
  assign tmp6129 = ~(s0 ? tmp3639 : tmp6130);
  assign tmp6126 = s1 ? tmp6127 : tmp6129;
  assign tmp6124 = ~(s2 ? tmp6125 : tmp6126);
  assign tmp6116 = s3 ? tmp6117 : tmp6124;
  assign tmp6135 = l1 ? tmp3434 : tmp4500;
  assign tmp6134 = s0 ? tmp6135 : tmp3486;
  assign tmp6137 = ~(l1 ? tmp3545 : tmp3775);
  assign tmp6136 = s0 ? tmp3486 : tmp6137;
  assign tmp6133 = s1 ? tmp6134 : tmp6136;
  assign tmp6140 = ~(l1 ? tmp3486 : tmp4454);
  assign tmp6139 = s0 ? tmp3434 : tmp6140;
  assign tmp6141 = ~(s0 ? tmp3639 : tmp3644);
  assign tmp6138 = ~(s1 ? tmp6139 : tmp6141);
  assign tmp6132 = s2 ? tmp6133 : tmp6138;
  assign tmp6144 = s0 ? 1 : tmp4115;
  assign tmp6145 = s0 ? tmp4059 : tmp6111;
  assign tmp6143 = s1 ? tmp6144 : tmp6145;
  assign tmp6147 = s0 ? tmp3639 : tmp6130;
  assign tmp6148 = s0 ? 1 : tmp3782;
  assign tmp6146 = ~(s1 ? tmp6147 : tmp6148);
  assign tmp6142 = s2 ? tmp6143 : tmp6146;
  assign tmp6131 = ~(s3 ? tmp6132 : tmp6142);
  assign tmp6115 = ~(s4 ? tmp6116 : tmp6131);
  assign tmp6078 = ~(s5 ? tmp6079 : tmp6115);
  assign tmp6049 = s6 ? tmp6050 : tmp6078;
  assign tmp6154 = l2 ? tmp4287 : tmp3420;
  assign tmp6153 = l1 ? tmp6154 : tmp4414;
  assign tmp6156 = l1 ? tmp3537 : tmp4414;
  assign tmp6155 = s0 ? tmp3459 : tmp6156;
  assign tmp6152 = s1 ? tmp6153 : tmp6155;
  assign tmp6159 = l1 ? tmp3420 : tmp3422;
  assign tmp6161 = l2 ? tmp4287 : tmp3538;
  assign tmp6160 = l1 ? tmp6161 : tmp4414;
  assign tmp6158 = s0 ? tmp6159 : tmp6160;
  assign tmp6163 = s0 ? tmp6159 : tmp3459;
  assign tmp6162 = s1 ? tmp6163 : tmp6160;
  assign tmp6157 = s2 ? tmp6158 : tmp6162;
  assign tmp6151 = s3 ? tmp6152 : tmp6157;
  assign tmp6168 = l1 ? tmp3544 : tmp4414;
  assign tmp6167 = s0 ? tmp6168 : 1;
  assign tmp6166 = s1 ? tmp6167 : tmp6160;
  assign tmp6170 = s0 ? tmp6153 : 1;
  assign tmp6169 = s1 ? tmp6170 : tmp5857;
  assign tmp6165 = s2 ? tmp6166 : tmp6169;
  assign tmp6175 = l2 ? tmp4287 : tmp3436;
  assign tmp6174 = l1 ? tmp6175 : tmp4414;
  assign tmp6173 = s0 ? tmp6160 : tmp6174;
  assign tmp6176 = s0 ? tmp6077 : tmp6160;
  assign tmp6172 = s1 ? tmp6173 : tmp6176;
  assign tmp6171 = s2 ? tmp6071 : tmp6172;
  assign tmp6164 = s3 ? tmp6165 : tmp6171;
  assign tmp6150 = s4 ? tmp6151 : tmp6164;
  assign tmp6182 = s0 ? tmp6156 : 1;
  assign tmp6184 = l1 ? tmp3544 : tmp3422;
  assign tmp6183 = s0 ? 1 : tmp6184;
  assign tmp6181 = s1 ? tmp6182 : tmp6183;
  assign tmp6187 = l1 ? tmp3537 : tmp4447;
  assign tmp6186 = s0 ? 1 : tmp6187;
  assign tmp6188 = s0 ? tmp6174 : tmp3459;
  assign tmp6185 = s1 ? tmp6186 : tmp6188;
  assign tmp6180 = s2 ? tmp6181 : tmp6185;
  assign tmp6192 = ~(l1 ? tmp4415 : tmp3436);
  assign tmp6191 = s0 ? tmp3459 : tmp6192;
  assign tmp6193 = s0 ? tmp3459 : tmp6095;
  assign tmp6190 = s1 ? tmp6191 : tmp6193;
  assign tmp6196 = l1 ? tmp6161 : tmp4447;
  assign tmp6197 = l1 ? tmp6175 : tmp4447;
  assign tmp6195 = s0 ? tmp6196 : tmp6197;
  assign tmp6194 = s1 ? tmp6097 : tmp6195;
  assign tmp6189 = s2 ? tmp6190 : tmp6194;
  assign tmp6179 = s3 ? tmp6180 : tmp6189;
  assign tmp6201 = s0 ? tmp6104 : tmp6196;
  assign tmp6200 = s1 ? tmp6201 : tmp3497;
  assign tmp6204 = l1 ? tmp3544 : tmp4447;
  assign tmp6203 = s0 ? tmp6204 : 1;
  assign tmp6202 = s1 ? tmp3497 : tmp6203;
  assign tmp6199 = s2 ? tmp6200 : tmp6202;
  assign tmp6208 = ~(l1 ? tmp6175 : tmp4470);
  assign tmp6207 = s0 ? tmp6107 : tmp6208;
  assign tmp6206 = s1 ? tmp6207 : tmp6112;
  assign tmp6205 = ~(s2 ? tmp6206 : tmp6113);
  assign tmp6198 = s3 ? tmp6199 : tmp6205;
  assign tmp6178 = s4 ? tmp6179 : tmp6198;
  assign tmp6213 = s0 ? 1 : tmp3624;
  assign tmp6214 = s0 ? tmp3644 : tmp3624;
  assign tmp6212 = ~(s1 ? tmp6213 : tmp6214);
  assign tmp6211 = s2 ? tmp6118 : tmp6212;
  assign tmp6210 = s3 ? tmp6211 : tmp6124;
  assign tmp6218 = ~(s0 ? tmp3624 : tmp3644);
  assign tmp6217 = ~(s1 ? tmp6139 : tmp6218);
  assign tmp6216 = s2 ? tmp6133 : tmp6217;
  assign tmp6215 = ~(s3 ? tmp6216 : tmp6142);
  assign tmp6209 = s4 ? tmp6210 : tmp6215;
  assign tmp6177 = s5 ? tmp6178 : tmp6209;
  assign tmp6149 = s6 ? tmp6150 : tmp6177;
  assign tmp6048 = s8 ? tmp6049 : tmp6149;
  assign tmp6224 = l1 ? tmp6154 : tmp3544;
  assign tmp6226 = l1 ? tmp3537 : tmp3544;
  assign tmp6225 = s0 ? tmp5534 : tmp6226;
  assign tmp6223 = s1 ? tmp6224 : tmp6225;
  assign tmp6229 = l1 ? tmp3420 : tmp3544;
  assign tmp6230 = l1 ? tmp6161 : tmp4538;
  assign tmp6228 = s0 ? tmp6229 : tmp6230;
  assign tmp6232 = s0 ? tmp6229 : 1;
  assign tmp6234 = l1 ? tmp6161 : tmp3544;
  assign tmp6233 = s0 ? tmp6230 : tmp6234;
  assign tmp6231 = s1 ? tmp6232 : tmp6233;
  assign tmp6227 = s2 ? tmp6228 : tmp6231;
  assign tmp6222 = s3 ? tmp6223 : tmp6227;
  assign tmp6238 = s0 ? tmp3544 : 1;
  assign tmp6239 = s0 ? tmp6234 : tmp6230;
  assign tmp6237 = s1 ? tmp6238 : tmp6239;
  assign tmp6241 = s0 ? tmp6224 : 1;
  assign tmp6240 = s1 ? tmp6241 : tmp4595;
  assign tmp6236 = s2 ? tmp6237 : tmp6240;
  assign tmp6243 = s1 ? tmp5554 : tmp5482;
  assign tmp6246 = l1 ? tmp6175 : tmp4538;
  assign tmp6245 = s0 ? tmp6230 : tmp6246;
  assign tmp6248 = l1 ? tmp3545 : tmp4538;
  assign tmp6247 = s0 ? tmp6248 : tmp6230;
  assign tmp6244 = s1 ? tmp6245 : tmp6247;
  assign tmp6242 = s2 ? tmp6243 : tmp6244;
  assign tmp6235 = s3 ? tmp6236 : tmp6242;
  assign tmp6221 = s4 ? tmp6222 : tmp6235;
  assign tmp6254 = s0 ? tmp6226 : 1;
  assign tmp6256 = l1 ? tmp3544 : 1;
  assign tmp6255 = s0 ? 1 : tmp6256;
  assign tmp6253 = s1 ? tmp6254 : tmp6255;
  assign tmp6258 = s0 ? 1 : tmp6226;
  assign tmp6259 = s0 ? tmp6246 : 1;
  assign tmp6257 = s1 ? tmp6258 : tmp6259;
  assign tmp6252 = s2 ? tmp6253 : tmp6257;
  assign tmp6264 = ~(l2 ? tmp3420 : 1);
  assign tmp6263 = ~(l1 ? tmp4415 : tmp6264);
  assign tmp6262 = s0 ? 1 : tmp6263;
  assign tmp6265 = s0 ? 1 : tmp6248;
  assign tmp6261 = s1 ? tmp6262 : tmp6265;
  assign tmp6267 = s0 ? tmp6248 : tmp4090;
  assign tmp6266 = s1 ? tmp6267 : tmp6245;
  assign tmp6260 = s2 ? tmp6261 : tmp6266;
  assign tmp6251 = s3 ? tmp6252 : tmp6260;
  assign tmp6271 = s0 ? tmp6104 : tmp6234;
  assign tmp6270 = s1 ? tmp6271 : tmp5586;
  assign tmp6272 = s1 ? tmp5586 : tmp6238;
  assign tmp6269 = s2 ? tmp6270 : tmp6272;
  assign tmp6276 = l1 ? tmp3434 : tmp6264;
  assign tmp6277 = ~(l1 ? tmp6175 : tmp3544);
  assign tmp6275 = s0 ? tmp6276 : tmp6277;
  assign tmp6278 = ~(s0 ? tmp4583 : tmp6077);
  assign tmp6274 = s1 ? tmp6275 : tmp6278;
  assign tmp6273 = ~(s2 ? tmp6274 : tmp6113);
  assign tmp6268 = s3 ? tmp6269 : tmp6273;
  assign tmp6250 = s4 ? tmp6251 : tmp6268;
  assign tmp6283 = s0 ? tmp6248 : tmp3434;
  assign tmp6284 = s0 ? tmp3434 : tmp4377;
  assign tmp6282 = s1 ? tmp6283 : tmp6284;
  assign tmp6286 = s0 ? tmp4333 : tmp3512;
  assign tmp6285 = ~(s1 ? tmp6286 : tmp4495);
  assign tmp6281 = s2 ? tmp6282 : tmp6285;
  assign tmp6288 = s1 ? tmp6120 : tmp5327;
  assign tmp6290 = ~(s0 ? tmp3639 : tmp3640);
  assign tmp6289 = s1 ? tmp6127 : tmp6290;
  assign tmp6287 = ~(s2 ? tmp6288 : tmp6289);
  assign tmp6280 = s3 ? tmp6281 : tmp6287;
  assign tmp6294 = s0 ? tmp3434 : tmp3486;
  assign tmp6296 = ~(l1 ? tmp3545 : tmp4538);
  assign tmp6295 = s0 ? tmp3486 : tmp6296;
  assign tmp6293 = s1 ? tmp6294 : tmp6295;
  assign tmp6299 = ~(l1 ? tmp3486 : tmp6264);
  assign tmp6298 = s0 ? tmp3434 : tmp6299;
  assign tmp6300 = ~(s0 ? tmp3512 : tmp3434);
  assign tmp6297 = ~(s1 ? tmp6298 : tmp6300);
  assign tmp6292 = s2 ? tmp6293 : tmp6297;
  assign tmp6303 = s0 ? tmp4333 : tmp4115;
  assign tmp6305 = ~(l1 ? tmp3545 : tmp3640);
  assign tmp6304 = s0 ? tmp4059 : tmp6305;
  assign tmp6302 = s1 ? tmp6303 : tmp6304;
  assign tmp6307 = s0 ? tmp3639 : tmp3640;
  assign tmp6306 = ~(s1 ? tmp6307 : tmp6148);
  assign tmp6301 = s2 ? tmp6302 : tmp6306;
  assign tmp6291 = ~(s3 ? tmp6292 : tmp6301);
  assign tmp6279 = s4 ? tmp6280 : tmp6291;
  assign tmp6249 = s5 ? tmp6250 : tmp6279;
  assign tmp6220 = s6 ? tmp6221 : tmp6249;
  assign tmp6219 = s8 ? tmp6149 : tmp6220;
  assign tmp6047 = s9 ? tmp6048 : tmp6219;
  assign tmp6312 = l1 ? tmp6154 : tmp4507;
  assign tmp6314 = l1 ? tmp3537 : tmp4507;
  assign tmp6313 = s0 ? tmp5534 : tmp6314;
  assign tmp6311 = s1 ? tmp6312 : tmp6313;
  assign tmp6317 = l1 ? tmp3420 : tmp3863;
  assign tmp6318 = l1 ? tmp6161 : tmp4515;
  assign tmp6316 = s0 ? tmp6317 : tmp6318;
  assign tmp6320 = s0 ? tmp6317 : 1;
  assign tmp6322 = l1 ? tmp6161 : tmp4507;
  assign tmp6321 = s0 ? tmp6318 : tmp6322;
  assign tmp6319 = s1 ? tmp6320 : tmp6321;
  assign tmp6315 = s2 ? tmp6316 : tmp6319;
  assign tmp6310 = s3 ? tmp6311 : tmp6315;
  assign tmp6327 = l1 ? tmp3544 : tmp4507;
  assign tmp6326 = s0 ? tmp6327 : 1;
  assign tmp6328 = s0 ? tmp6322 : tmp6318;
  assign tmp6325 = s1 ? tmp6326 : tmp6328;
  assign tmp6330 = s0 ? tmp6312 : 1;
  assign tmp6329 = s1 ? tmp6330 : tmp4595;
  assign tmp6324 = s2 ? tmp6325 : tmp6329;
  assign tmp6334 = l1 ? tmp6175 : tmp4515;
  assign tmp6333 = s0 ? tmp6318 : tmp6334;
  assign tmp6335 = s0 ? tmp6248 : tmp6318;
  assign tmp6332 = s1 ? tmp6333 : tmp6335;
  assign tmp6331 = s2 ? tmp6243 : tmp6332;
  assign tmp6323 = s3 ? tmp6324 : tmp6331;
  assign tmp6309 = s4 ? tmp6310 : tmp6323;
  assign tmp6341 = s0 ? tmp6314 : 1;
  assign tmp6343 = l1 ? tmp3544 : tmp3486;
  assign tmp6342 = s0 ? 1 : tmp6343;
  assign tmp6340 = s1 ? tmp6341 : tmp6342;
  assign tmp6346 = l1 ? tmp3537 : tmp4549;
  assign tmp6345 = s0 ? 1 : tmp6346;
  assign tmp6347 = s0 ? tmp6334 : 1;
  assign tmp6344 = s1 ? tmp6345 : tmp6347;
  assign tmp6339 = s2 ? tmp6340 : tmp6344;
  assign tmp6352 = ~(l2 ? tmp3420 : tmp3422);
  assign tmp6351 = ~(l1 ? tmp4415 : tmp6352);
  assign tmp6350 = s0 ? 1 : tmp6351;
  assign tmp6354 = l1 ? tmp3545 : tmp4561;
  assign tmp6353 = s0 ? 1 : tmp6354;
  assign tmp6349 = s1 ? tmp6350 : tmp6353;
  assign tmp6357 = l1 ? tmp6161 : tmp4561;
  assign tmp6358 = l1 ? tmp6175 : tmp4561;
  assign tmp6356 = s0 ? tmp6357 : tmp6358;
  assign tmp6355 = s1 ? tmp6267 : tmp6356;
  assign tmp6348 = s2 ? tmp6349 : tmp6355;
  assign tmp6338 = s3 ? tmp6339 : tmp6348;
  assign tmp6363 = l1 ? tmp6161 : tmp4549;
  assign tmp6362 = s0 ? tmp6104 : tmp6363;
  assign tmp6361 = s1 ? tmp6362 : tmp5586;
  assign tmp6366 = l1 ? tmp3544 : tmp4549;
  assign tmp6365 = s0 ? tmp6366 : 1;
  assign tmp6364 = s1 ? tmp5586 : tmp6365;
  assign tmp6360 = s2 ? tmp6361 : tmp6364;
  assign tmp6371 = ~(l2 ? tmp3420 : tmp3424);
  assign tmp6370 = l1 ? tmp3434 : tmp6371;
  assign tmp6372 = ~(l1 ? tmp6175 : tmp4549);
  assign tmp6369 = s0 ? tmp6370 : tmp6372;
  assign tmp6373 = ~(s0 ? tmp4583 : tmp6095);
  assign tmp6368 = s1 ? tmp6369 : tmp6373;
  assign tmp6367 = ~(s2 ? tmp6368 : tmp6113);
  assign tmp6359 = s3 ? tmp6360 : tmp6367;
  assign tmp6337 = s4 ? tmp6338 : tmp6359;
  assign tmp6378 = s0 ? tmp6354 : tmp3434;
  assign tmp6377 = s1 ? tmp6378 : tmp6284;
  assign tmp6380 = s0 ? tmp4333 : tmp3639;
  assign tmp6379 = ~(s1 ? tmp6380 : tmp6123);
  assign tmp6376 = s2 ? tmp6377 : tmp6379;
  assign tmp6375 = s3 ? tmp6376 : tmp6124;
  assign tmp6383 = s1 ? tmp6134 : tmp6295;
  assign tmp6386 = ~(l1 ? tmp3486 : tmp6371);
  assign tmp6385 = s0 ? tmp3434 : tmp6386;
  assign tmp6384 = ~(s1 ? tmp6385 : tmp6141);
  assign tmp6382 = s2 ? tmp6383 : tmp6384;
  assign tmp6388 = s1 ? tmp6303 : tmp6145;
  assign tmp6387 = s2 ? tmp6388 : tmp6146;
  assign tmp6381 = ~(s3 ? tmp6382 : tmp6387);
  assign tmp6374 = s4 ? tmp6375 : tmp6381;
  assign tmp6336 = s5 ? tmp6337 : tmp6374;
  assign tmp6308 = s6 ? tmp6309 : tmp6336;
  assign tmp6046 = s10 ? tmp6047 : tmp6308;
  assign tmp5804 = s12 ? tmp5805 : tmp6046;
  assign tmp6396 = l1 ? 1 : tmp4500;
  assign tmp6399 = l2 ? 1 : tmp4287;
  assign tmp6398 = l1 ? tmp6399 : tmp4500;
  assign tmp6397 = s0 ? 1 : tmp6398;
  assign tmp6395 = s1 ? tmp6396 : tmp6397;
  assign tmp6401 = s1 ? 1 : tmp6398;
  assign tmp6400 = s2 ? tmp6397 : tmp6401;
  assign tmp6394 = s3 ? tmp6395 : tmp6400;
  assign tmp6405 = s0 ? tmp6396 : 1;
  assign tmp6404 = s1 ? tmp6405 : tmp6398;
  assign tmp6406 = s1 ? tmp6405 : 1;
  assign tmp6403 = s2 ? tmp6404 : tmp6406;
  assign tmp6409 = s0 ? 1 : tmp5314;
  assign tmp6408 = s1 ? 1 : tmp6409;
  assign tmp6411 = s0 ? tmp5286 : tmp6398;
  assign tmp6410 = s1 ? tmp6398 : tmp6411;
  assign tmp6407 = s2 ? tmp6408 : tmp6410;
  assign tmp6402 = s3 ? tmp6403 : tmp6407;
  assign tmp6393 = s4 ? tmp6394 : tmp6402;
  assign tmp6417 = s0 ? tmp6398 : 1;
  assign tmp6416 = s1 ? tmp6417 : 1;
  assign tmp6418 = s1 ? tmp6397 : tmp6417;
  assign tmp6415 = s2 ? tmp6416 : tmp6418;
  assign tmp6422 = l1 ? tmp6399 : tmp4608;
  assign tmp6421 = s0 ? 1 : tmp6422;
  assign tmp6420 = s1 ? 1 : tmp6421;
  assign tmp6424 = s0 ? tmp5286 : tmp5314;
  assign tmp6423 = s1 ? tmp6424 : tmp6422;
  assign tmp6419 = s2 ? tmp6420 : tmp6423;
  assign tmp6414 = s3 ? tmp6415 : tmp6419;
  assign tmp6428 = s0 ? tmp3475 : tmp6422;
  assign tmp6427 = s1 ? tmp6428 : 1;
  assign tmp6429 = s1 ? 1 : tmp6405;
  assign tmp6426 = s2 ? tmp6427 : tmp6429;
  assign tmp6433 = l1 ? 1 : tmp4608;
  assign tmp6432 = s0 ? tmp6396 : tmp6433;
  assign tmp6431 = s1 ? tmp6432 : tmp6421;
  assign tmp6435 = s0 ? tmp5314 : tmp3434;
  assign tmp6434 = s1 ? tmp3434 : tmp6435;
  assign tmp6430 = s2 ? tmp6431 : tmp6434;
  assign tmp6425 = s3 ? tmp6426 : tmp6430;
  assign tmp6413 = s4 ? tmp6414 : tmp6425;
  assign tmp6440 = s0 ? tmp6422 : 1;
  assign tmp6439 = s1 ? tmp6440 : 1;
  assign tmp6438 = s2 ? tmp6439 : 1;
  assign tmp6443 = ~(s0 ? 1 : tmp5311);
  assign tmp6442 = s1 ? tmp3803 : tmp6443;
  assign tmp6445 = s0 ? tmp5314 : tmp3475;
  assign tmp6446 = s0 ? tmp3475 : tmp4500;
  assign tmp6444 = s1 ? tmp6445 : tmp6446;
  assign tmp6441 = s2 ? tmp6442 : tmp6444;
  assign tmp6437 = s3 ? tmp6438 : tmp6441;
  assign tmp6450 = s0 ? tmp4500 : tmp4115;
  assign tmp6451 = s0 ? tmp4115 : tmp5286;
  assign tmp6449 = s1 ? tmp6450 : tmp6451;
  assign tmp6452 = s1 ? tmp6397 : 1;
  assign tmp6448 = s2 ? tmp6449 : tmp6452;
  assign tmp6455 = s0 ? 1 : tmp5286;
  assign tmp6456 = s0 ? tmp5314 : tmp6422;
  assign tmp6454 = s1 ? tmp6455 : tmp6456;
  assign tmp6459 = ~(l1 ? tmp3486 : 0);
  assign tmp6458 = ~(s0 ? 1 : tmp6459);
  assign tmp6457 = s1 ? tmp6446 : tmp6458;
  assign tmp6453 = s2 ? tmp6454 : tmp6457;
  assign tmp6447 = s3 ? tmp6448 : tmp6453;
  assign tmp6436 = s4 ? tmp6437 : tmp6447;
  assign tmp6412 = s5 ? tmp6413 : tmp6436;
  assign tmp6392 = s6 ? tmp6393 : tmp6412;
  assign tmp6466 = l2 ? 1 : tmp3548;
  assign tmp6465 = l1 ? 1 : tmp6466;
  assign tmp6468 = l1 ? tmp6399 : tmp3486;
  assign tmp6467 = s0 ? 1 : tmp6468;
  assign tmp6464 = s1 ? tmp6465 : tmp6467;
  assign tmp6471 = l1 ? tmp6399 : tmp6466;
  assign tmp6470 = s0 ? 1 : tmp6471;
  assign tmp6472 = s1 ? 1 : tmp6471;
  assign tmp6469 = s2 ? tmp6470 : tmp6472;
  assign tmp6463 = s3 ? tmp6464 : tmp6469;
  assign tmp6477 = l1 ? 1 : tmp3486;
  assign tmp6476 = s0 ? tmp6477 : 1;
  assign tmp6475 = s1 ? tmp6476 : tmp6471;
  assign tmp6479 = s0 ? tmp6465 : 1;
  assign tmp6478 = s1 ? tmp6479 : 1;
  assign tmp6474 = s2 ? tmp6475 : tmp6478;
  assign tmp6482 = s0 ? tmp5286 : tmp6471;
  assign tmp6481 = s1 ? tmp6471 : tmp6482;
  assign tmp6480 = s2 ? tmp6408 : tmp6481;
  assign tmp6473 = s3 ? tmp6474 : tmp6480;
  assign tmp6462 = s4 ? tmp6463 : tmp6473;
  assign tmp6488 = s0 ? tmp6468 : 1;
  assign tmp6487 = s1 ? tmp6488 : 1;
  assign tmp6491 = l1 ? tmp6399 : tmp3434;
  assign tmp6490 = s0 ? 1 : tmp6491;
  assign tmp6492 = s0 ? tmp6471 : 1;
  assign tmp6489 = s1 ? tmp6490 : tmp6492;
  assign tmp6486 = s2 ? tmp6487 : tmp6489;
  assign tmp6494 = s1 ? 1 : tmp6490;
  assign tmp6495 = s1 ? tmp6424 : tmp6491;
  assign tmp6493 = s2 ? tmp6494 : tmp6495;
  assign tmp6485 = s3 ? tmp6486 : tmp6493;
  assign tmp6499 = s0 ? tmp3475 : tmp6491;
  assign tmp6498 = s1 ? tmp6499 : 1;
  assign tmp6500 = s1 ? 1 : tmp4192;
  assign tmp6497 = s2 ? tmp6498 : tmp6500;
  assign tmp6502 = s1 ? tmp3475 : tmp6490;
  assign tmp6501 = s2 ? tmp6502 : tmp6434;
  assign tmp6496 = s3 ? tmp6497 : tmp6501;
  assign tmp6484 = s4 ? tmp6485 : tmp6496;
  assign tmp6507 = s0 ? tmp6491 : 1;
  assign tmp6506 = s1 ? tmp6507 : 1;
  assign tmp6505 = s2 ? tmp6506 : 1;
  assign tmp6509 = s1 ? tmp6445 : tmp3475;
  assign tmp6508 = s2 ? tmp6442 : tmp6509;
  assign tmp6504 = s3 ? tmp6505 : tmp6508;
  assign tmp6513 = s0 ? tmp3475 : tmp4115;
  assign tmp6512 = s1 ? tmp6513 : tmp6451;
  assign tmp6514 = s1 ? tmp6490 : 1;
  assign tmp6511 = s2 ? tmp6512 : tmp6514;
  assign tmp6517 = s0 ? tmp5314 : tmp6491;
  assign tmp6516 = s1 ? tmp6455 : tmp6517;
  assign tmp6518 = s1 ? tmp3475 : tmp6458;
  assign tmp6515 = s2 ? tmp6516 : tmp6518;
  assign tmp6510 = s3 ? tmp6511 : tmp6515;
  assign tmp6503 = s4 ? tmp6504 : tmp6510;
  assign tmp6483 = s5 ? tmp6484 : tmp6503;
  assign tmp6461 = s6 ? tmp6462 : tmp6483;
  assign tmp6460 = s8 ? tmp6392 : tmp6461;
  assign tmp6391 = s9 ? tmp6392 : tmp6460;
  assign tmp6390 = s10 ? tmp6391 : tmp6392;
  assign tmp6526 = l1 ? tmp3494 : tmp3486;
  assign tmp6527 = ~(l1 ? tmp3429 : tmp3782);
  assign tmp6525 = s1 ? tmp6526 : tmp6527;
  assign tmp6531 = ~(l1 ? tmp3494 : tmp3486);
  assign tmp6530 = s0 ? tmp3646 : tmp6531;
  assign tmp6533 = l1 ? tmp3429 : tmp3782;
  assign tmp6532 = s0 ? tmp6533 : tmp6531;
  assign tmp6529 = s1 ? tmp6530 : tmp6532;
  assign tmp6535 = s0 ? tmp6533 : 0;
  assign tmp6534 = s1 ? tmp6535 : tmp6531;
  assign tmp6528 = ~(s2 ? tmp6529 : tmp6534);
  assign tmp6524 = s3 ? tmp6525 : tmp6528;
  assign tmp6539 = s0 ? tmp5766 : 0;
  assign tmp6538 = s1 ? tmp6539 : tmp6531;
  assign tmp6541 = s0 ? tmp6526 : 1;
  assign tmp6540 = ~(s1 ? tmp6541 : 1);
  assign tmp6537 = s2 ? tmp6538 : tmp6540;
  assign tmp6545 = l1 ? tmp3434 : tmp3486;
  assign tmp6544 = s0 ? 1 : tmp6545;
  assign tmp6543 = s1 ? 1 : tmp6544;
  assign tmp6548 = l1 ? tmp3448 : tmp3486;
  assign tmp6547 = s0 ? tmp6526 : tmp6548;
  assign tmp6550 = l1 ? tmp3427 : tmp3486;
  assign tmp6549 = s0 ? tmp6550 : tmp6526;
  assign tmp6546 = s1 ? tmp6547 : tmp6549;
  assign tmp6542 = ~(s2 ? tmp6543 : tmp6546);
  assign tmp6536 = ~(s3 ? tmp6537 : tmp6542);
  assign tmp6523 = s4 ? tmp6524 : tmp6536;
  assign tmp6555 = s1 ? tmp6535 : tmp6085;
  assign tmp6558 = ~(l1 ? tmp3429 : tmp3640);
  assign tmp6557 = s0 ? 1 : tmp6558;
  assign tmp6559 = s0 ? tmp6548 : 1;
  assign tmp6556 = ~(s1 ? tmp6557 : tmp6559);
  assign tmp6554 = s2 ? tmp6555 : tmp6556;
  assign tmp6563 = ~(l1 ? tmp3486 : tmp3782);
  assign tmp6562 = s0 ? 1 : tmp6563;
  assign tmp6564 = s0 ? 1 : tmp6548;
  assign tmp6561 = s1 ? tmp6562 : tmp6564;
  assign tmp6566 = s0 ? tmp6550 : tmp3644;
  assign tmp6565 = s1 ? tmp6566 : tmp6547;
  assign tmp6560 = ~(s2 ? tmp6561 : tmp6565);
  assign tmp6553 = s3 ? tmp6554 : tmp6560;
  assign tmp6570 = s0 ? tmp6545 : tmp6526;
  assign tmp6569 = s1 ? tmp6570 : 1;
  assign tmp6572 = ~(s0 ? tmp3639 : 0);
  assign tmp6571 = s1 ? 1 : tmp6572;
  assign tmp6568 = s2 ? tmp6569 : tmp6571;
  assign tmp6576 = ~(l1 ? tmp3545 : tmp3486);
  assign tmp6575 = s0 ? tmp3639 : tmp6576;
  assign tmp6577 = ~(s0 ? 1 : tmp6548);
  assign tmp6574 = s1 ? tmp6575 : tmp6577;
  assign tmp6579 = s0 ? tmp6545 : 1;
  assign tmp6578 = ~(s1 ? 1 : tmp6579);
  assign tmp6573 = ~(s2 ? tmp6574 : tmp6578);
  assign tmp6567 = ~(s3 ? tmp6568 : tmp6573);
  assign tmp6552 = s4 ? tmp6553 : tmp6567;
  assign tmp6584 = s0 ? tmp6548 : tmp3434;
  assign tmp6585 = s0 ? tmp3434 : tmp3457;
  assign tmp6583 = s1 ? tmp6584 : tmp6585;
  assign tmp6587 = s0 ? tmp3460 : tmp3639;
  assign tmp6586 = ~(s1 ? tmp6587 : tmp6123);
  assign tmp6582 = s2 ? tmp6583 : tmp6586;
  assign tmp6590 = s0 ? tmp3644 : tmp3913;
  assign tmp6589 = s1 ? tmp6590 : tmp4248;
  assign tmp6593 = ~(l1 ? tmp3434 : tmp3486);
  assign tmp6592 = s0 ? tmp3460 : tmp6593;
  assign tmp6594 = ~(s0 ? tmp6545 : tmp6128);
  assign tmp6591 = s1 ? tmp6592 : tmp6594;
  assign tmp6588 = ~(s2 ? tmp6589 : tmp6591);
  assign tmp6581 = s3 ? tmp6582 : tmp6588;
  assign tmp6598 = s0 ? tmp3639 : 1;
  assign tmp6600 = ~(l1 ? tmp3427 : tmp3486);
  assign tmp6599 = s0 ? 1 : tmp6600;
  assign tmp6597 = s1 ? tmp6598 : tmp6599;
  assign tmp6603 = ~(l1 ? tmp4418 : tmp3640);
  assign tmp6602 = s0 ? tmp3434 : tmp6603;
  assign tmp6601 = ~(s1 ? tmp6602 : tmp6141);
  assign tmp6596 = s2 ? tmp6597 : tmp6601;
  assign tmp6606 = s0 ? tmp3460 : tmp3913;
  assign tmp6608 = ~(l1 ? tmp3448 : tmp3486);
  assign tmp6607 = s0 ? tmp3460 : tmp6608;
  assign tmp6605 = s1 ? tmp6606 : tmp6607;
  assign tmp6610 = s0 ? tmp6545 : tmp6128;
  assign tmp6611 = ~(s0 ? tmp3913 : 1);
  assign tmp6609 = ~(s1 ? tmp6610 : tmp6611);
  assign tmp6604 = s2 ? tmp6605 : tmp6609;
  assign tmp6595 = ~(s3 ? tmp6596 : tmp6604);
  assign tmp6580 = ~(s4 ? tmp6581 : tmp6595);
  assign tmp6551 = ~(s5 ? tmp6552 : tmp6580);
  assign tmp6522 = s6 ? tmp6523 : tmp6551;
  assign tmp6616 = l1 ? tmp6154 : tmp5053;
  assign tmp6617 = l1 ? tmp3420 : tmp5053;
  assign tmp6615 = s1 ? tmp6616 : tmp6617;
  assign tmp6620 = s0 ? tmp6184 : tmp6616;
  assign tmp6621 = s0 ? tmp6617 : tmp6616;
  assign tmp6619 = s1 ? tmp6620 : tmp6621;
  assign tmp6623 = s0 ? tmp6617 : tmp3459;
  assign tmp6622 = s1 ? tmp6623 : tmp6616;
  assign tmp6618 = s2 ? tmp6619 : tmp6622;
  assign tmp6614 = s3 ? tmp6615 : tmp6618;
  assign tmp6628 = l1 ? tmp3544 : tmp5053;
  assign tmp6627 = s0 ? tmp6628 : 1;
  assign tmp6626 = s1 ? tmp6627 : tmp6616;
  assign tmp6630 = s0 ? tmp6616 : 1;
  assign tmp6632 = l1 ? 1 : tmp4415;
  assign tmp6631 = s0 ? tmp6632 : 1;
  assign tmp6629 = s1 ? tmp6630 : tmp6631;
  assign tmp6625 = s2 ? tmp6626 : tmp6629;
  assign tmp6636 = l1 ? 1 : tmp5045;
  assign tmp6635 = s0 ? tmp6632 : tmp6636;
  assign tmp6634 = s1 ? tmp6635 : tmp6544;
  assign tmp6640 = l2 ? tmp4287 : tmp3423;
  assign tmp6639 = l1 ? tmp6640 : tmp5053;
  assign tmp6638 = s0 ? tmp6616 : tmp6639;
  assign tmp6643 = ~(l2 ? tmp3420 : tmp3436);
  assign tmp6642 = l1 ? tmp3427 : tmp6643;
  assign tmp6641 = s0 ? tmp6642 : tmp6616;
  assign tmp6637 = s1 ? tmp6638 : tmp6641;
  assign tmp6633 = s2 ? tmp6634 : tmp6637;
  assign tmp6624 = s3 ? tmp6625 : tmp6633;
  assign tmp6613 = s4 ? tmp6614 : tmp6624;
  assign tmp6649 = s0 ? tmp6617 : 1;
  assign tmp6648 = s1 ? tmp6649 : tmp6183;
  assign tmp6653 = l2 ? tmp4415 : 0;
  assign tmp6652 = l1 ? tmp3420 : tmp6653;
  assign tmp6651 = s0 ? 1 : tmp6652;
  assign tmp6654 = s0 ? tmp6639 : tmp3459;
  assign tmp6650 = s1 ? tmp6651 : tmp6654;
  assign tmp6647 = s2 ? tmp6648 : tmp6650;
  assign tmp6659 = ~(l2 ? tmp4415 : tmp3422);
  assign tmp6658 = ~(l1 ? tmp4415 : tmp6659);
  assign tmp6657 = s0 ? tmp3459 : tmp6658;
  assign tmp6661 = l1 ? tmp3448 : tmp5053;
  assign tmp6660 = s0 ? tmp3459 : tmp6661;
  assign tmp6656 = s1 ? tmp6657 : tmp6660;
  assign tmp6663 = s0 ? tmp6642 : tmp3644;
  assign tmp6665 = l1 ? tmp6640 : tmp6643;
  assign tmp6664 = s0 ? tmp6616 : tmp6665;
  assign tmp6662 = s1 ? tmp6663 : tmp6664;
  assign tmp6655 = s2 ? tmp6656 : tmp6662;
  assign tmp6646 = s3 ? tmp6647 : tmp6655;
  assign tmp6669 = s0 ? tmp6545 : tmp6616;
  assign tmp6668 = s1 ? tmp6669 : tmp4400;
  assign tmp6672 = l1 ? tmp3544 : tmp6653;
  assign tmp6671 = s0 ? tmp6672 : 1;
  assign tmp6670 = s1 ? tmp4400 : tmp6671;
  assign tmp6667 = s2 ? tmp6668 : tmp6670;
  assign tmp6677 = ~(l2 ? tmp4415 : 0);
  assign tmp6676 = l1 ? tmp3434 : tmp6677;
  assign tmp6678 = ~(l1 ? tmp6175 : tmp6643);
  assign tmp6675 = s0 ? tmp6676 : tmp6678;
  assign tmp6679 = ~(s0 ? tmp4333 : tmp6548);
  assign tmp6674 = s1 ? tmp6675 : tmp6679;
  assign tmp6673 = ~(s2 ? tmp6674 : tmp6578);
  assign tmp6666 = s3 ? tmp6667 : tmp6673;
  assign tmp6645 = s4 ? tmp6646 : tmp6666;
  assign tmp6684 = s0 ? tmp6661 : tmp3434;
  assign tmp6685 = s0 ? tmp3434 : tmp4686;
  assign tmp6683 = s1 ? tmp6684 : tmp6685;
  assign tmp6687 = s0 ? tmp4583 : tmp3624;
  assign tmp6686 = ~(s1 ? tmp6687 : tmp6214);
  assign tmp6682 = s2 ? tmp6683 : tmp6686;
  assign tmp6681 = s3 ? tmp6682 : tmp6588;
  assign tmp6692 = ~(l1 ? tmp3427 : tmp6643);
  assign tmp6691 = s0 ? 1 : tmp6692;
  assign tmp6690 = s1 ? tmp6598 : tmp6691;
  assign tmp6695 = ~(l1 ? tmp4418 : tmp6677);
  assign tmp6694 = s0 ? tmp3434 : tmp6695;
  assign tmp6693 = ~(s1 ? tmp6694 : tmp6218);
  assign tmp6689 = s2 ? tmp6690 : tmp6693;
  assign tmp6698 = s0 ? tmp4583 : tmp3913;
  assign tmp6697 = s1 ? tmp6698 : tmp6607;
  assign tmp6696 = s2 ? tmp6697 : tmp6609;
  assign tmp6688 = ~(s3 ? tmp6689 : tmp6696);
  assign tmp6680 = s4 ? tmp6681 : tmp6688;
  assign tmp6644 = s5 ? tmp6645 : tmp6680;
  assign tmp6612 = s6 ? tmp6613 : tmp6644;
  assign tmp6521 = s8 ? tmp6522 : tmp6612;
  assign tmp6704 = l1 ? tmp6154 : tmp3486;
  assign tmp6705 = l1 ? tmp3420 : tmp3486;
  assign tmp6703 = s1 ? tmp6704 : tmp6705;
  assign tmp6708 = s0 ? tmp6256 : tmp6704;
  assign tmp6710 = l1 ? tmp3420 : 1;
  assign tmp6709 = s0 ? tmp6710 : tmp6704;
  assign tmp6707 = s1 ? tmp6708 : tmp6709;
  assign tmp6712 = s0 ? tmp6710 : 1;
  assign tmp6711 = s1 ? tmp6712 : tmp6704;
  assign tmp6706 = s2 ? tmp6707 : tmp6711;
  assign tmp6702 = s3 ? tmp6703 : tmp6706;
  assign tmp6716 = s0 ? tmp6343 : 1;
  assign tmp6715 = s1 ? tmp6716 : tmp6704;
  assign tmp6718 = s0 ? tmp6704 : 1;
  assign tmp6717 = s1 ? tmp6718 : 1;
  assign tmp6714 = s2 ? tmp6715 : tmp6717;
  assign tmp6722 = l1 ? tmp6640 : tmp3486;
  assign tmp6721 = s0 ? tmp6704 : tmp6722;
  assign tmp6723 = s0 ? tmp6550 : tmp6704;
  assign tmp6720 = s1 ? tmp6721 : tmp6723;
  assign tmp6719 = s2 ? tmp6543 : tmp6720;
  assign tmp6713 = s3 ? tmp6714 : tmp6719;
  assign tmp6701 = s4 ? tmp6702 : tmp6713;
  assign tmp6729 = s0 ? tmp6705 : 1;
  assign tmp6728 = s1 ? tmp6729 : tmp6255;
  assign tmp6732 = l1 ? tmp3420 : tmp3434;
  assign tmp6731 = s0 ? 1 : tmp6732;
  assign tmp6733 = s0 ? tmp6722 : 1;
  assign tmp6730 = s1 ? tmp6731 : tmp6733;
  assign tmp6727 = s2 ? tmp6728 : tmp6730;
  assign tmp6737 = ~(l1 ? tmp4415 : 0);
  assign tmp6736 = s0 ? 1 : tmp6737;
  assign tmp6735 = s1 ? tmp6736 : tmp6564;
  assign tmp6738 = s1 ? tmp6566 : tmp6721;
  assign tmp6734 = s2 ? tmp6735 : tmp6738;
  assign tmp6726 = s3 ? tmp6727 : tmp6734;
  assign tmp6742 = s0 ? tmp6545 : tmp6704;
  assign tmp6741 = s1 ? tmp6742 : 1;
  assign tmp6745 = l1 ? tmp3544 : tmp3434;
  assign tmp6744 = s0 ? tmp6745 : 1;
  assign tmp6743 = s1 ? 1 : tmp6744;
  assign tmp6740 = s2 ? tmp6741 : tmp6743;
  assign tmp6749 = ~(l1 ? tmp6175 : tmp3486);
  assign tmp6748 = s0 ? tmp3639 : tmp6749;
  assign tmp6747 = s1 ? tmp6748 : tmp6577;
  assign tmp6746 = ~(s2 ? tmp6747 : tmp6578);
  assign tmp6739 = s3 ? tmp6740 : tmp6746;
  assign tmp6725 = s4 ? tmp6726 : tmp6739;
  assign tmp6753 = ~(s1 ? tmp4874 : tmp4495);
  assign tmp6752 = s2 ? tmp6583 : tmp6753;
  assign tmp6756 = s0 ? tmp3434 : tmp3913;
  assign tmp6755 = s1 ? tmp6756 : tmp4248;
  assign tmp6754 = ~(s2 ? tmp6755 : tmp6591);
  assign tmp6751 = s3 ? tmp6752 : tmp6754;
  assign tmp6759 = ~(s1 ? tmp6602 : tmp6300);
  assign tmp6758 = s2 ? tmp6597 : tmp6759;
  assign tmp6757 = ~(s3 ? tmp6758 : tmp6604);
  assign tmp6750 = s4 ? tmp6751 : tmp6757;
  assign tmp6724 = s5 ? tmp6725 : tmp6750;
  assign tmp6700 = s6 ? tmp6701 : tmp6724;
  assign tmp6699 = s8 ? tmp6612 : tmp6700;
  assign tmp6520 = s9 ? tmp6521 : tmp6699;
  assign tmp6765 = s0 ? tmp6343 : tmp6704;
  assign tmp6766 = s0 ? tmp6705 : tmp6704;
  assign tmp6764 = s1 ? tmp6765 : tmp6766;
  assign tmp6767 = s1 ? tmp6729 : tmp6704;
  assign tmp6763 = s2 ? tmp6764 : tmp6767;
  assign tmp6762 = s3 ? tmp6703 : tmp6763;
  assign tmp6761 = s4 ? tmp6762 : tmp6713;
  assign tmp6772 = s1 ? tmp6729 : tmp6342;
  assign tmp6771 = s2 ? tmp6772 : tmp6730;
  assign tmp6776 = ~(l1 ? tmp4415 : tmp3782);
  assign tmp6775 = s0 ? 1 : tmp6776;
  assign tmp6774 = s1 ? tmp6775 : tmp6564;
  assign tmp6773 = s2 ? tmp6774 : tmp6738;
  assign tmp6770 = s3 ? tmp6771 : tmp6773;
  assign tmp6769 = s4 ? tmp6770 : tmp6739;
  assign tmp6777 = s4 ? tmp6581 : tmp6595;
  assign tmp6768 = s5 ? tmp6769 : tmp6777;
  assign tmp6760 = s6 ? tmp6761 : tmp6768;
  assign tmp6519 = s10 ? tmp6520 : tmp6760;
  assign tmp6389 = s12 ? tmp6390 : tmp6519;
  assign tmp5803 = ~(s13 ? tmp5804 : tmp6389);
  assign tmp5231 = ~(s14 ? tmp5232 : tmp5803);
  assign tmp3407 = s15 ? tmp3408 : tmp5231;
  assign tmp6782 = s9 ? tmp3412 : tmp3532;
  assign tmp6781 = s10 ? tmp6782 : tmp3532;
  assign tmp6791 = l1 ? tmp3789 : tmp3530;
  assign tmp6790 = s1 ? tmp6791 : tmp4098;
  assign tmp6795 = l1 ? tmp3863 : tmp3640;
  assign tmp6794 = s0 ? tmp6795 : tmp6791;
  assign tmp6797 = l1 ? tmp3789 : tmp3640;
  assign tmp6796 = s0 ? tmp6797 : tmp6791;
  assign tmp6793 = s1 ? tmp6794 : tmp6796;
  assign tmp6799 = s0 ? tmp6797 : tmp3845;
  assign tmp6798 = s1 ? tmp6799 : tmp6791;
  assign tmp6792 = s2 ? tmp6793 : tmp6798;
  assign tmp6789 = s3 ? tmp6790 : tmp6792;
  assign tmp6802 = s1 ? tmp4111 : tmp6791;
  assign tmp6804 = s0 ? tmp6791 : 1;
  assign tmp6803 = s1 ? tmp6804 : tmp4114;
  assign tmp6801 = s2 ? tmp6802 : tmp6803;
  assign tmp6808 = ~(l1 ? tmp3789 : tmp3530);
  assign tmp6807 = ~(s0 ? 1 : tmp6808);
  assign tmp6806 = s1 ? tmp6791 : tmp6807;
  assign tmp6805 = s2 ? tmp4117 : tmp6806;
  assign tmp6800 = s3 ? tmp6801 : tmp6805;
  assign tmp6788 = s4 ? tmp6789 : tmp6800;
  assign tmp6814 = s0 ? tmp3845 : tmp6795;
  assign tmp6813 = s1 ? tmp4107 : tmp6814;
  assign tmp6817 = l1 ? tmp3822 : tmp3530;
  assign tmp6816 = s0 ? tmp6817 : tmp3845;
  assign tmp6815 = s1 ? tmp4128 : tmp6816;
  assign tmp6812 = s2 ? tmp6813 : tmp6815;
  assign tmp6821 = l1 ? tmp3822 : tmp3640;
  assign tmp6820 = s0 ? tmp3845 : tmp6821;
  assign tmp6819 = s1 ? tmp6820 : tmp4136;
  assign tmp6818 = s2 ? tmp6819 : tmp4137;
  assign tmp6811 = s3 ? tmp6812 : tmp6818;
  assign tmp6810 = s4 ? tmp6811 : tmp4140;
  assign tmp6809 = s5 ? tmp6810 : 0;
  assign tmp6787 = s6 ? tmp6788 : tmp6809;
  assign tmp6786 = ~(s8 ? tmp4154 : tmp6787);
  assign tmp6785 = s9 ? tmp4035 : tmp6786;
  assign tmp6784 = s10 ? tmp6785 : tmp4092;
  assign tmp6783 = s12 ? tmp3762 : tmp6784;
  assign tmp6780 = s13 ? tmp6781 : tmp6783;
  assign tmp6831 = l2 ? tmp4287 : tmp3548;
  assign tmp6830 = l1 ? tmp3822 : tmp6831;
  assign tmp6833 = l1 ? tmp3434 : tmp4538;
  assign tmp6834 = l1 ? tmp3822 : tmp4706;
  assign tmp6832 = s0 ? tmp6833 : tmp6834;
  assign tmp6829 = s1 ? tmp6830 : tmp6832;
  assign tmp6838 = l1 ? tmp3822 : tmp3486;
  assign tmp6839 = l1 ? tmp3822 : tmp3789;
  assign tmp6837 = s0 ? tmp6838 : tmp6839;
  assign tmp6840 = s0 ? tmp6834 : tmp6839;
  assign tmp6836 = s1 ? tmp6837 : tmp6840;
  assign tmp6842 = s0 ? tmp6834 : tmp3644;
  assign tmp6843 = s0 ? tmp6839 : tmp6830;
  assign tmp6841 = s1 ? tmp6842 : tmp6843;
  assign tmp6835 = s2 ? tmp6836 : tmp6841;
  assign tmp6828 = s3 ? tmp6829 : tmp6835;
  assign tmp6847 = s0 ? tmp6830 : tmp6839;
  assign tmp6846 = s1 ? tmp6842 : tmp6847;
  assign tmp6849 = s0 ? tmp6830 : tmp3644;
  assign tmp6851 = l1 ? tmp3434 : tmp4287;
  assign tmp6850 = s0 ? tmp6851 : tmp3644;
  assign tmp6848 = s1 ? tmp6849 : tmp6850;
  assign tmp6845 = s2 ? tmp6846 : tmp6848;
  assign tmp6853 = s1 ? tmp6833 : tmp5400;
  assign tmp6855 = s0 ? tmp6839 : tmp3789;
  assign tmp6856 = s0 ? tmp3420 : tmp6839;
  assign tmp6854 = s1 ? tmp6855 : tmp6856;
  assign tmp6852 = s2 ? tmp6853 : tmp6854;
  assign tmp6844 = s3 ? tmp6845 : tmp6852;
  assign tmp6827 = s4 ? tmp6828 : tmp6844;
  assign tmp6862 = s0 ? tmp6834 : tmp3457;
  assign tmp6864 = ~(l1 ? tmp3822 : tmp3486);
  assign tmp6863 = ~(s0 ? tmp3460 : tmp6864);
  assign tmp6861 = s1 ? tmp6862 : tmp6863;
  assign tmp6868 = l2 ? tmp4287 : 0;
  assign tmp6867 = ~(l1 ? tmp3822 : tmp6868);
  assign tmp6866 = s0 ? tmp3460 : tmp6867;
  assign tmp6865 = ~(s1 ? tmp6866 : tmp4270);
  assign tmp6860 = s2 ? tmp6861 : tmp6865;
  assign tmp6871 = s0 ? 1 : tmp6834;
  assign tmp6870 = s1 ? tmp6871 : tmp3821;
  assign tmp6872 = s1 ? tmp3509 : tmp3822;
  assign tmp6869 = s2 ? tmp6870 : tmp6872;
  assign tmp6859 = s3 ? tmp6860 : tmp6869;
  assign tmp6876 = s0 ? 1 : tmp6867;
  assign tmp6877 = ~(s0 ? tmp3644 : tmp4783);
  assign tmp6875 = s1 ? tmp6876 : tmp6877;
  assign tmp6879 = s0 ? tmp3644 : tmp4783;
  assign tmp6881 = l1 ? tmp3822 : tmp6868;
  assign tmp6880 = s0 ? tmp6881 : tmp3644;
  assign tmp6878 = ~(s1 ? tmp6879 : tmp6880);
  assign tmp6874 = s2 ? tmp6875 : tmp6878;
  assign tmp6884 = s0 ? tmp4319 : tmp4275;
  assign tmp6885 = ~(s0 ? tmp4783 : 0);
  assign tmp6883 = s1 ? tmp6884 : tmp6885;
  assign tmp6882 = s2 ? tmp6883 : 1;
  assign tmp6873 = ~(s3 ? tmp6874 : tmp6882);
  assign tmp6858 = s4 ? tmp6859 : tmp6873;
  assign tmp6886 = s4 ? tmp4341 : tmp4347;
  assign tmp6857 = s5 ? tmp6858 : tmp6886;
  assign tmp6826 = s6 ? tmp6827 : tmp6857;
  assign tmp6892 = l1 ? tmp3822 : tmp6154;
  assign tmp6894 = l1 ? tmp3822 : tmp4287;
  assign tmp6893 = s0 ? tmp6833 : tmp6894;
  assign tmp6891 = s1 ? tmp6892 : tmp6893;
  assign tmp6898 = l1 ? tmp3822 : 1;
  assign tmp6899 = l1 ? tmp3822 : tmp3420;
  assign tmp6897 = s0 ? tmp6898 : tmp6899;
  assign tmp6901 = l1 ? tmp3822 : tmp4538;
  assign tmp6900 = s0 ? tmp6901 : tmp6899;
  assign tmp6896 = s1 ? tmp6897 : tmp6900;
  assign tmp6903 = s0 ? tmp6901 : tmp3644;
  assign tmp6904 = s0 ? tmp6899 : tmp6892;
  assign tmp6902 = s1 ? tmp6903 : tmp6904;
  assign tmp6895 = s2 ? tmp6896 : tmp6902;
  assign tmp6890 = s3 ? tmp6891 : tmp6895;
  assign tmp6908 = s0 ? tmp6894 : tmp3644;
  assign tmp6909 = s0 ? tmp6892 : tmp6899;
  assign tmp6907 = s1 ? tmp6908 : tmp6909;
  assign tmp6911 = s0 ? tmp6892 : tmp3644;
  assign tmp6910 = s1 ? tmp6911 : tmp6850;
  assign tmp6906 = s2 ? tmp6907 : tmp6910;
  assign tmp6914 = s0 ? tmp3420 : tmp6899;
  assign tmp6913 = s1 ? tmp6899 : tmp6914;
  assign tmp6912 = s2 ? tmp6853 : tmp6913;
  assign tmp6905 = s3 ? tmp6906 : tmp6912;
  assign tmp6889 = s4 ? tmp6890 : tmp6905;
  assign tmp6920 = s0 ? tmp6894 : tmp3457;
  assign tmp6922 = ~(l1 ? tmp3822 : 1);
  assign tmp6921 = ~(s0 ? tmp3460 : tmp6922);
  assign tmp6919 = s1 ? tmp6920 : tmp6921;
  assign tmp6925 = ~(l1 ? tmp3822 : tmp4287);
  assign tmp6924 = s0 ? tmp3460 : tmp6925;
  assign tmp6926 = ~(s0 ? tmp6899 : 1);
  assign tmp6923 = ~(s1 ? tmp6924 : tmp6926);
  assign tmp6918 = s2 ? tmp6919 : tmp6923;
  assign tmp6929 = s0 ? 1 : tmp6901;
  assign tmp6930 = s0 ? 1 : tmp4377;
  assign tmp6928 = s1 ? tmp6929 : tmp6930;
  assign tmp6931 = s1 ? tmp3509 : tmp6899;
  assign tmp6927 = s2 ? tmp6928 : tmp6931;
  assign tmp6917 = s3 ? tmp6918 : tmp6927;
  assign tmp6934 = ~(s1 ? tmp6879 : tmp6908);
  assign tmp6933 = s2 ? tmp6875 : tmp6934;
  assign tmp6937 = s0 ? tmp4306 : tmp4275;
  assign tmp6936 = s1 ? tmp6937 : tmp6885;
  assign tmp6935 = s2 ? tmp6936 : 1;
  assign tmp6932 = ~(s3 ? tmp6933 : tmp6935);
  assign tmp6916 = s4 ? tmp6917 : tmp6932;
  assign tmp6938 = ~(s4 ? tmp4397 : tmp4402);
  assign tmp6915 = s5 ? tmp6916 : tmp6938;
  assign tmp6888 = s6 ? tmp6889 : tmp6915;
  assign tmp6887 = s8 ? tmp6826 : tmp6888;
  assign tmp6825 = s9 ? tmp6826 : tmp6887;
  assign tmp6824 = s10 ? tmp6825 : tmp6826;
  assign tmp6943 = l1 ? tmp3582 : tmp4435;
  assign tmp6945 = l1 ? tmp3438 : tmp4435;
  assign tmp6944 = s0 ? tmp3795 : tmp6945;
  assign tmp6942 = s1 ? tmp6943 : tmp6944;
  assign tmp6948 = l1 ? tmp3582 : tmp3436;
  assign tmp6947 = s0 ? tmp6948 : tmp6945;
  assign tmp6950 = s0 ? tmp6948 : tmp3646;
  assign tmp6949 = s1 ? tmp6950 : tmp6945;
  assign tmp6946 = s2 ? tmp6947 : tmp6949;
  assign tmp6941 = s3 ? tmp6942 : tmp6946;
  assign tmp6955 = l1 ? tmp3781 : 0;
  assign tmp6954 = s0 ? tmp6943 : tmp6955;
  assign tmp6953 = s1 ? tmp6954 : tmp6945;
  assign tmp6957 = s0 ? tmp6943 : tmp3434;
  assign tmp6958 = s0 ? tmp3795 : tmp3434;
  assign tmp6956 = s1 ? tmp6957 : tmp6958;
  assign tmp6952 = s2 ? tmp6953 : tmp6956;
  assign tmp6961 = s0 ? tmp3434 : tmp3607;
  assign tmp6960 = s1 ? tmp3795 : tmp6961;
  assign tmp6963 = s0 ? tmp6945 : tmp4449;
  assign tmp6965 = ~(l1 ? tmp3438 : tmp4435);
  assign tmp6964 = ~(s0 ? tmp3868 : tmp6965);
  assign tmp6962 = s1 ? tmp6963 : tmp6964;
  assign tmp6959 = s2 ? tmp6960 : tmp6962;
  assign tmp6951 = s3 ? tmp6952 : tmp6959;
  assign tmp6940 = s4 ? tmp6941 : tmp6951;
  assign tmp6971 = s0 ? tmp6945 : 0;
  assign tmp6973 = ~(l1 ? tmp3582 : tmp3436);
  assign tmp6972 = ~(s0 ? 1 : tmp6973);
  assign tmp6970 = s1 ? tmp6971 : tmp6972;
  assign tmp6976 = ~(l1 ? tmp3438 : tmp4454);
  assign tmp6975 = s0 ? 1 : tmp6976;
  assign tmp6977 = ~(s0 ? tmp4449 : tmp3913);
  assign tmp6974 = ~(s1 ? tmp6975 : tmp6977);
  assign tmp6969 = s2 ? tmp6970 : tmp6974;
  assign tmp6980 = s0 ? tmp3913 : tmp6948;
  assign tmp6981 = s0 ? tmp3913 : tmp4472;
  assign tmp6979 = s1 ? tmp6980 : tmp6981;
  assign tmp6984 = l1 ? tmp3438 : tmp4454;
  assign tmp6983 = ~(s0 ? tmp6984 : tmp4472);
  assign tmp6982 = ~(s1 ? tmp4456 : tmp6983);
  assign tmp6978 = s2 ? tmp6979 : tmp6982;
  assign tmp6968 = s3 ? tmp6969 : tmp6978;
  assign tmp6988 = s0 ? tmp3868 : tmp6976;
  assign tmp6989 = ~(s0 ? tmp6955 : 1);
  assign tmp6987 = s1 ? tmp6988 : tmp6989;
  assign tmp6991 = s0 ? tmp6955 : 1;
  assign tmp6993 = l1 ? tmp3582 : tmp4454;
  assign tmp6992 = s0 ? tmp6993 : tmp6955;
  assign tmp6990 = ~(s1 ? tmp6991 : tmp6992);
  assign tmp6986 = s2 ? tmp6987 : tmp6990;
  assign tmp6997 = ~(l1 ? tmp3582 : tmp4500);
  assign tmp6996 = s0 ? tmp4468 : tmp6997;
  assign tmp6995 = s1 ? tmp6996 : tmp4471;
  assign tmp6994 = s2 ? tmp6995 : tmp4473;
  assign tmp6985 = ~(s3 ? tmp6986 : tmp6994);
  assign tmp6967 = s4 ? tmp6968 : tmp6985;
  assign tmp7003 = l1 ? tmp3434 : tmp3427;
  assign tmp7002 = s0 ? tmp3460 : tmp7003;
  assign tmp7004 = s0 ? tmp3512 : tmp7003;
  assign tmp7001 = ~(s1 ? tmp7002 : tmp7004);
  assign tmp7000 = s2 ? tmp4478 : tmp7001;
  assign tmp6999 = s3 ? tmp7000 : tmp4483;
  assign tmp7008 = s0 ? tmp7003 : tmp3512;
  assign tmp7007 = s1 ? tmp4493 : tmp7008;
  assign tmp7006 = s2 ? tmp4489 : tmp7007;
  assign tmp7005 = ~(s3 ? tmp7006 : tmp4496);
  assign tmp6998 = s4 ? tmp6999 : tmp7005;
  assign tmp6966 = s5 ? tmp6967 : tmp6998;
  assign tmp6939 = s6 ? tmp6940 : tmp6966;
  assign tmp6823 = s12 ? tmp6824 : tmp6939;
  assign tmp7011 = s9 ? tmp4599 : tmp4701;
  assign tmp7010 = s10 ? tmp7011 : tmp4701;
  assign tmp7009 = ~(s12 ? tmp7010 : tmp4960);
  assign tmp6822 = ~(s13 ? tmp6823 : tmp7009);
  assign tmp6779 = s14 ? tmp6780 : tmp6822;
  assign tmp7016 = s9 ? tmp6048 : tmp6149;
  assign tmp7015 = s10 ? tmp7016 : tmp6149;
  assign tmp7014 = s12 ? tmp5805 : tmp7015;
  assign tmp7013 = ~(s13 ? tmp7014 : tmp6389);
  assign tmp7012 = ~(s14 ? tmp5232 : tmp7013);
  assign tmp6778 = s15 ? tmp6779 : tmp7012;
  assign tmp3406 = s16 ? tmp3407 : tmp6778;
  assign tmp7025 = ~(s6 ? tmp4356 : tmp4378);
  assign tmp7024 = s8 ? tmp6826 : tmp7025;
  assign tmp7023 = s9 ? tmp6826 : tmp7024;
  assign tmp7026 = ~(s6 ? tmp4282 : tmp4312);
  assign tmp7022 = s10 ? tmp7023 : tmp7026;
  assign tmp7035 = l1 ? tmp4418 : tmp3544;
  assign tmp7034 = s0 ? tmp4509 : tmp7035;
  assign tmp7033 = s1 ? tmp4509 : tmp7034;
  assign tmp7039 = l1 ? tmp4418 : tmp4538;
  assign tmp7038 = s0 ? tmp3685 : tmp7039;
  assign tmp7040 = s0 ? tmp4509 : tmp7039;
  assign tmp7037 = s1 ? tmp7038 : tmp7040;
  assign tmp7042 = s0 ? tmp4509 : 1;
  assign tmp7043 = s0 ? tmp7039 : tmp7035;
  assign tmp7041 = s1 ? tmp7042 : tmp7043;
  assign tmp7036 = s2 ? tmp7037 : tmp7041;
  assign tmp7032 = s3 ? tmp7033 : tmp7036;
  assign tmp7047 = s0 ? tmp4509 : tmp3685;
  assign tmp7048 = s0 ? tmp7035 : tmp7039;
  assign tmp7046 = s1 ? tmp7047 : tmp7048;
  assign tmp7049 = s1 ? tmp7042 : tmp4528;
  assign tmp7045 = s2 ? tmp7046 : tmp7049;
  assign tmp7053 = l1 ? tmp3429 : tmp4538;
  assign tmp7052 = s0 ? tmp7039 : tmp7053;
  assign tmp7054 = s0 ? tmp4537 : tmp7039;
  assign tmp7051 = s1 ? tmp7052 : tmp7054;
  assign tmp7050 = s2 ? tmp4531 : tmp7051;
  assign tmp7044 = s3 ? tmp7045 : tmp7050;
  assign tmp7031 = s4 ? tmp7032 : tmp7044;
  assign tmp7060 = s0 ? tmp7035 : 1;
  assign tmp7061 = s0 ? 1 : tmp3685;
  assign tmp7059 = s1 ? tmp7060 : tmp7061;
  assign tmp7063 = s0 ? 1 : tmp7035;
  assign tmp7064 = s0 ? tmp7053 : 1;
  assign tmp7062 = s1 ? tmp7063 : tmp7064;
  assign tmp7058 = s2 ? tmp7059 : tmp7062;
  assign tmp7067 = s0 ? 1 : tmp4509;
  assign tmp7069 = ~(l1 ? tmp3420 : tmp4290);
  assign tmp7068 = s0 ? 1 : tmp7069;
  assign tmp7066 = s1 ? tmp7067 : tmp7068;
  assign tmp7070 = s1 ? tmp4558 : tmp7052;
  assign tmp7065 = s2 ? tmp7066 : tmp7070;
  assign tmp7057 = s3 ? tmp7058 : tmp7065;
  assign tmp7074 = s0 ? tmp3868 : tmp7035;
  assign tmp7073 = s1 ? tmp7074 : tmp4567;
  assign tmp7075 = s1 ? tmp4567 : tmp7047;
  assign tmp7072 = s2 ? tmp7073 : tmp7075;
  assign tmp7079 = l1 ? tmp3434 : tmp3544;
  assign tmp7078 = s0 ? tmp7079 : tmp4509;
  assign tmp7081 = ~(l1 ? tmp3420 : tmp3607);
  assign tmp7080 = s0 ? tmp3822 : tmp7081;
  assign tmp7077 = s1 ? tmp7078 : tmp7080;
  assign tmp7076 = s2 ? tmp7077 : tmp4473;
  assign tmp7071 = s3 ? tmp7072 : tmp7076;
  assign tmp7056 = s4 ? tmp7057 : tmp7071;
  assign tmp7087 = l1 ? tmp3420 : tmp4290;
  assign tmp7086 = s0 ? tmp7087 : 0;
  assign tmp7085 = s1 ? tmp7086 : tmp4582;
  assign tmp7089 = s0 ? tmp4583 : tmp3644;
  assign tmp7090 = s0 ? tmp3434 : tmp3644;
  assign tmp7088 = ~(s1 ? tmp7089 : tmp7090);
  assign tmp7084 = s2 ? tmp7085 : tmp7088;
  assign tmp7093 = s0 ? tmp3845 : tmp3639;
  assign tmp7092 = s1 ? tmp3844 : tmp7093;
  assign tmp7091 = ~(s2 ? tmp3697 : tmp7092);
  assign tmp7083 = s3 ? tmp7084 : tmp7091;
  assign tmp7096 = s1 ? tmp6598 : tmp4589;
  assign tmp7099 = l1 ? tmp3429 : tmp3544;
  assign tmp7098 = s0 ? 1 : tmp7099;
  assign tmp7100 = s0 ? tmp3644 : tmp3434;
  assign tmp7097 = s1 ? tmp7098 : tmp7100;
  assign tmp7095 = s2 ? tmp7096 : tmp7097;
  assign tmp7104 = ~(l1 ? tmp3420 : tmp3434);
  assign tmp7103 = s0 ? 1 : tmp7104;
  assign tmp7102 = s1 ? tmp4595 : tmp7103;
  assign tmp7105 = s1 ? tmp7093 : 1;
  assign tmp7101 = s2 ? tmp7102 : tmp7105;
  assign tmp7094 = ~(s3 ? tmp7095 : tmp7101);
  assign tmp7082 = ~(s4 ? tmp7083 : tmp7094);
  assign tmp7055 = s5 ? tmp7056 : tmp7082;
  assign tmp7030 = ~(s6 ? tmp7031 : tmp7055);
  assign tmp7029 = s8 ? tmp6939 : tmp7030;
  assign tmp7028 = s9 ? tmp6939 : tmp7029;
  assign tmp7106 = ~(s6 ? tmp4503 : tmp4539);
  assign tmp7027 = s10 ? tmp7028 : tmp7106;
  assign tmp7021 = s12 ? tmp7022 : tmp7027;
  assign tmp7107 = ~(s12 ? tmp4597 : tmp4960);
  assign tmp7020 = ~(s13 ? tmp7021 : tmp7107);
  assign tmp7019 = s14 ? tmp3409 : tmp7020;
  assign tmp7018 = s15 ? tmp7019 : tmp5231;
  assign tmp7017 = s16 ? tmp7018 : tmp6778;
  assign tmp3405 = s17 ? tmp3406 : tmp7017;
  assign recovery__2 = tmp3405;

  assign tmp7123 = ~(l2 ? 1 : 0);
  assign tmp7122 = l1 ? 1 : tmp7123;
  assign tmp7125 = l1 ? 1 : 0;
  assign tmp7124 = s0 ? tmp7125 : tmp7122;
  assign tmp7121 = s1 ? tmp7122 : tmp7124;
  assign tmp7128 = s0 ? tmp7122 : tmp7125;
  assign tmp7127 = s1 ? tmp7128 : tmp7122;
  assign tmp7126 = s2 ? tmp7122 : tmp7127;
  assign tmp7120 = s3 ? tmp7121 : tmp7126;
  assign tmp7132 = s0 ? tmp7122 : 1;
  assign tmp7133 = s0 ? tmp7125 : 1;
  assign tmp7131 = s1 ? tmp7132 : tmp7133;
  assign tmp7130 = s2 ? tmp7127 : tmp7131;
  assign tmp7135 = s1 ? tmp7125 : 1;
  assign tmp7137 = s0 ? tmp7122 : tmp7123;
  assign tmp7138 = s0 ? 1 : tmp7122;
  assign tmp7136 = s1 ? tmp7137 : tmp7138;
  assign tmp7134 = s2 ? tmp7135 : tmp7136;
  assign tmp7129 = s3 ? tmp7130 : tmp7134;
  assign tmp7119 = s4 ? tmp7120 : tmp7129;
  assign tmp7143 = s1 ? tmp7128 : tmp7124;
  assign tmp7146 = l2 ? 1 : 0;
  assign tmp7145 = ~(s0 ? tmp7146 : 1);
  assign tmp7144 = s1 ? tmp7124 : tmp7145;
  assign tmp7142 = s2 ? tmp7143 : tmp7144;
  assign tmp7148 = s0 ? 1 : tmp7146;
  assign tmp7149 = ~(s1 ? 1 : tmp7132);
  assign tmp7147 = ~(s2 ? tmp7148 : tmp7149);
  assign tmp7141 = s3 ? tmp7142 : tmp7147;
  assign tmp7152 = s1 ? tmp7138 : tmp7133;
  assign tmp7153 = s1 ? tmp7133 : tmp7128;
  assign tmp7151 = s2 ? tmp7152 : tmp7153;
  assign tmp7155 = s1 ? tmp7146 : 0;
  assign tmp7154 = ~(s2 ? tmp7155 : 0);
  assign tmp7150 = s3 ? tmp7151 : tmp7154;
  assign tmp7140 = s4 ? tmp7141 : tmp7150;
  assign tmp7160 = s0 ? tmp7146 : 0;
  assign tmp7159 = s1 ? tmp7160 : 0;
  assign tmp7162 = s0 ? 1 : tmp7123;
  assign tmp7161 = ~(s1 ? tmp7162 : tmp7123);
  assign tmp7158 = s2 ? tmp7159 : tmp7161;
  assign tmp7157 = s3 ? tmp7158 : 0;
  assign tmp7165 = s1 ? tmp7162 : tmp7123;
  assign tmp7164 = s2 ? 1 : tmp7165;
  assign tmp7163 = ~(s3 ? tmp7164 : 1);
  assign tmp7156 = ~(s4 ? tmp7157 : tmp7163);
  assign tmp7139 = s5 ? tmp7140 : tmp7156;
  assign tmp7118 = s6 ? tmp7119 : tmp7139;
  assign tmp7170 = s1 ? tmp7132 : tmp7125;
  assign tmp7169 = s2 ? tmp7127 : tmp7170;
  assign tmp7168 = s3 ? tmp7169 : tmp7134;
  assign tmp7167 = s4 ? tmp7120 : tmp7168;
  assign tmp7175 = s1 ? tmp7122 : tmp7145;
  assign tmp7174 = s2 ? tmp7127 : tmp7175;
  assign tmp7176 = ~(s2 ? tmp7146 : tmp7149);
  assign tmp7173 = s3 ? tmp7174 : tmp7176;
  assign tmp7179 = s1 ? tmp7125 : tmp7128;
  assign tmp7178 = s2 ? tmp7152 : tmp7179;
  assign tmp7177 = s3 ? tmp7178 : tmp7154;
  assign tmp7172 = s4 ? tmp7173 : tmp7177;
  assign tmp7182 = s2 ? tmp7159 : tmp7155;
  assign tmp7181 = s3 ? tmp7182 : 0;
  assign tmp7184 = s2 ? 1 : tmp7123;
  assign tmp7183 = ~(s3 ? tmp7184 : 1);
  assign tmp7180 = ~(s4 ? tmp7181 : tmp7183);
  assign tmp7171 = s5 ? tmp7172 : tmp7180;
  assign tmp7166 = s6 ? tmp7167 : tmp7171;
  assign tmp7117 = s7 ? tmp7118 : tmp7166;
  assign tmp7190 = s1 ? tmp7122 : tmp7138;
  assign tmp7189 = s2 ? tmp7135 : tmp7190;
  assign tmp7188 = s3 ? tmp7130 : tmp7189;
  assign tmp7187 = s4 ? tmp7120 : tmp7188;
  assign tmp7195 = s1 ? tmp7124 : tmp7128;
  assign tmp7194 = s2 ? tmp7143 : tmp7195;
  assign tmp7198 = s0 ? tmp7125 : tmp7123;
  assign tmp7197 = s1 ? tmp7124 : tmp7198;
  assign tmp7199 = s1 ? 1 : tmp7132;
  assign tmp7196 = s2 ? tmp7197 : tmp7199;
  assign tmp7193 = s3 ? tmp7194 : tmp7196;
  assign tmp7201 = ~(s2 ? tmp7159 : 0);
  assign tmp7200 = s3 ? tmp7151 : tmp7201;
  assign tmp7192 = s4 ? tmp7193 : tmp7200;
  assign tmp7191 = s5 ? tmp7192 : tmp7156;
  assign tmp7186 = s6 ? tmp7187 : tmp7191;
  assign tmp7204 = s3 ? tmp7169 : tmp7189;
  assign tmp7203 = s4 ? tmp7120 : tmp7204;
  assign tmp7209 = s1 ? tmp7122 : tmp7128;
  assign tmp7208 = s2 ? tmp7127 : tmp7209;
  assign tmp7211 = s1 ? tmp7122 : tmp7123;
  assign tmp7210 = s2 ? tmp7211 : tmp7199;
  assign tmp7207 = s3 ? tmp7208 : tmp7210;
  assign tmp7213 = s2 ? tmp7152 : tmp7122;
  assign tmp7212 = s3 ? tmp7213 : tmp7201;
  assign tmp7206 = s4 ? tmp7207 : tmp7212;
  assign tmp7205 = s5 ? tmp7206 : tmp7180;
  assign tmp7202 = s6 ? tmp7203 : tmp7205;
  assign tmp7185 = s7 ? tmp7186 : tmp7202;
  assign tmp7116 = s8 ? tmp7117 : tmp7185;
  assign tmp7219 = s2 ? tmp7125 : tmp7133;
  assign tmp7222 = s0 ? 1 : tmp7125;
  assign tmp7221 = s1 ? tmp7125 : tmp7222;
  assign tmp7220 = s2 ? tmp7135 : tmp7221;
  assign tmp7218 = s3 ? tmp7219 : tmp7220;
  assign tmp7217 = s4 ? tmp7125 : tmp7218;
  assign tmp7228 = s0 ? tmp7125 : 0;
  assign tmp7227 = s1 ? tmp7125 : tmp7228;
  assign tmp7226 = s2 ? tmp7125 : tmp7227;
  assign tmp7231 = ~(l1 ? 1 : 0);
  assign tmp7230 = s0 ? 1 : tmp7231;
  assign tmp7232 = ~(s1 ? 1 : tmp7133);
  assign tmp7229 = ~(s2 ? tmp7230 : tmp7232);
  assign tmp7225 = s3 ? tmp7226 : tmp7229;
  assign tmp7235 = s1 ? tmp7222 : tmp7133;
  assign tmp7236 = s1 ? tmp7133 : tmp7125;
  assign tmp7234 = s2 ? tmp7235 : tmp7236;
  assign tmp7237 = s2 ? tmp7125 : 1;
  assign tmp7233 = s3 ? tmp7234 : tmp7237;
  assign tmp7224 = s4 ? tmp7225 : tmp7233;
  assign tmp7241 = s1 ? tmp7133 : 1;
  assign tmp7242 = s1 ? tmp7222 : tmp7125;
  assign tmp7240 = s2 ? tmp7241 : tmp7242;
  assign tmp7239 = s3 ? tmp7240 : 1;
  assign tmp7244 = s2 ? 1 : tmp7242;
  assign tmp7243 = s3 ? tmp7244 : 1;
  assign tmp7238 = s4 ? tmp7239 : tmp7243;
  assign tmp7223 = s5 ? tmp7224 : tmp7238;
  assign tmp7216 = s6 ? tmp7217 : tmp7223;
  assign tmp7248 = s2 ? tmp7125 : tmp7236;
  assign tmp7247 = s3 ? tmp7248 : tmp7220;
  assign tmp7246 = s4 ? tmp7125 : tmp7247;
  assign tmp7253 = s1 ? 1 : tmp7133;
  assign tmp7252 = s2 ? tmp7125 : tmp7253;
  assign tmp7251 = s3 ? tmp7226 : tmp7252;
  assign tmp7255 = s2 ? tmp7235 : tmp7125;
  assign tmp7256 = s2 ? tmp7135 : 1;
  assign tmp7254 = s3 ? tmp7255 : tmp7256;
  assign tmp7250 = s4 ? tmp7251 : tmp7254;
  assign tmp7259 = s2 ? tmp7241 : tmp7135;
  assign tmp7258 = s3 ? tmp7259 : 1;
  assign tmp7261 = s2 ? 1 : tmp7125;
  assign tmp7260 = s3 ? tmp7261 : 1;
  assign tmp7257 = s4 ? tmp7258 : tmp7260;
  assign tmp7249 = s5 ? tmp7250 : tmp7257;
  assign tmp7245 = s6 ? tmp7246 : tmp7249;
  assign tmp7215 = s7 ? tmp7216 : tmp7245;
  assign tmp7214 = s8 ? tmp7185 : tmp7215;
  assign tmp7115 = s9 ? tmp7116 : tmp7214;
  assign tmp7268 = s3 ? tmp7213 : tmp7154;
  assign tmp7267 = s4 ? tmp7173 : tmp7268;
  assign tmp7266 = s5 ? tmp7267 : tmp7180;
  assign tmp7265 = s6 ? tmp7167 : tmp7266;
  assign tmp7264 = s7 ? tmp7118 : tmp7265;
  assign tmp7263 = s8 ? tmp7264 : tmp7118;
  assign tmp7276 = s1 ? tmp7125 : tmp7122;
  assign tmp7275 = s2 ? tmp7152 : tmp7276;
  assign tmp7274 = s3 ? tmp7275 : tmp7154;
  assign tmp7273 = s4 ? tmp7173 : tmp7274;
  assign tmp7272 = s5 ? tmp7273 : tmp7180;
  assign tmp7271 = s6 ? tmp7167 : tmp7272;
  assign tmp7270 = s7 ? tmp7271 : tmp7245;
  assign tmp7277 = s7 ? tmp7202 : tmp7265;
  assign tmp7269 = s8 ? tmp7270 : tmp7277;
  assign tmp7262 = s9 ? tmp7263 : tmp7269;
  assign tmp7114 = s10 ? tmp7115 : tmp7262;
  assign tmp7281 = s7 ? tmp7166 : tmp7245;
  assign tmp7280 = s8 ? tmp7281 : tmp7277;
  assign tmp7279 = s9 ? tmp7263 : tmp7280;
  assign tmp7278 = s10 ? tmp7115 : tmp7279;
  assign tmp7113 = s11 ? tmp7114 : tmp7278;
  assign tmp7293 = ~(s0 ? 1 : tmp7231);
  assign tmp7292 = s1 ? tmp7228 : tmp7293;
  assign tmp7291 = s2 ? tmp7227 : tmp7292;
  assign tmp7290 = s3 ? tmp7125 : tmp7291;
  assign tmp7289 = s4 ? tmp7125 : tmp7290;
  assign tmp7298 = s1 ? tmp7125 : 0;
  assign tmp7297 = s2 ? tmp7125 : tmp7298;
  assign tmp7301 = ~(s0 ? tmp7125 : 0);
  assign tmp7300 = s1 ? 1 : tmp7301;
  assign tmp7299 = ~(s2 ? 1 : tmp7300);
  assign tmp7296 = s3 ? tmp7297 : tmp7299;
  assign tmp7304 = s1 ? tmp7230 : tmp7301;
  assign tmp7305 = ~(s1 ? tmp7228 : tmp7125);
  assign tmp7303 = s2 ? tmp7304 : tmp7305;
  assign tmp7302 = ~(s3 ? tmp7303 : 1);
  assign tmp7295 = s4 ? tmp7296 : tmp7302;
  assign tmp7294 = s5 ? tmp7295 : 0;
  assign tmp7288 = s6 ? tmp7289 : tmp7294;
  assign tmp7310 = s2 ? tmp7304 : tmp7231;
  assign tmp7309 = ~(s3 ? tmp7310 : 1);
  assign tmp7308 = s4 ? tmp7296 : tmp7309;
  assign tmp7307 = s5 ? tmp7308 : 0;
  assign tmp7306 = s6 ? tmp7289 : tmp7307;
  assign tmp7287 = s7 ? tmp7288 : tmp7306;
  assign tmp7316 = s1 ? tmp7125 : tmp7293;
  assign tmp7315 = s2 ? tmp7227 : tmp7316;
  assign tmp7314 = s3 ? tmp7125 : tmp7315;
  assign tmp7313 = s4 ? tmp7125 : tmp7314;
  assign tmp7322 = ~(s0 ? tmp7125 : 1);
  assign tmp7321 = ~(s1 ? 1 : tmp7322);
  assign tmp7320 = s2 ? tmp7227 : tmp7321;
  assign tmp7319 = s3 ? tmp7125 : tmp7320;
  assign tmp7325 = s1 ? tmp7230 : tmp7322;
  assign tmp7326 = ~(s1 ? tmp7133 : tmp7125);
  assign tmp7324 = s2 ? tmp7325 : tmp7326;
  assign tmp7329 = s0 ? 1 : 0;
  assign tmp7330 = ~(s0 ? 1 : 0);
  assign tmp7328 = s1 ? tmp7329 : tmp7330;
  assign tmp7327 = s2 ? tmp7328 : 1;
  assign tmp7323 = ~(s3 ? tmp7324 : tmp7327);
  assign tmp7318 = s4 ? tmp7319 : tmp7323;
  assign tmp7317 = s5 ? tmp7318 : 0;
  assign tmp7312 = s6 ? tmp7313 : tmp7317;
  assign tmp7334 = s2 ? tmp7298 : tmp7316;
  assign tmp7333 = s3 ? tmp7125 : tmp7334;
  assign tmp7332 = s4 ? tmp7125 : tmp7333;
  assign tmp7338 = s2 ? tmp7298 : tmp7321;
  assign tmp7337 = s3 ? tmp7125 : tmp7338;
  assign tmp7340 = s2 ? tmp7325 : tmp7231;
  assign tmp7342 = s1 ? tmp7329 : 1;
  assign tmp7341 = s2 ? tmp7342 : 1;
  assign tmp7339 = ~(s3 ? tmp7340 : tmp7341);
  assign tmp7336 = s4 ? tmp7337 : tmp7339;
  assign tmp7335 = s5 ? tmp7336 : 0;
  assign tmp7331 = s6 ? tmp7332 : tmp7335;
  assign tmp7311 = s7 ? tmp7312 : tmp7331;
  assign tmp7286 = s8 ? tmp7287 : tmp7311;
  assign tmp7350 = s1 ? tmp7230 : tmp7231;
  assign tmp7349 = s2 ? tmp7350 : tmp7231;
  assign tmp7348 = ~(s3 ? tmp7349 : 1);
  assign tmp7347 = s4 ? tmp7296 : tmp7348;
  assign tmp7346 = s5 ? tmp7347 : 0;
  assign tmp7345 = s6 ? tmp7289 : tmp7346;
  assign tmp7354 = s2 ? tmp7298 : tmp7292;
  assign tmp7353 = s3 ? tmp7125 : tmp7354;
  assign tmp7352 = s4 ? tmp7125 : tmp7353;
  assign tmp7351 = s6 ? tmp7352 : tmp7346;
  assign tmp7344 = s7 ? tmp7345 : tmp7351;
  assign tmp7343 = s8 ? tmp7311 : tmp7344;
  assign tmp7285 = s9 ? tmp7286 : tmp7343;
  assign tmp7356 = s8 ? tmp7344 : tmp7345;
  assign tmp7359 = s6 ? tmp7352 : tmp7307;
  assign tmp7358 = s7 ? tmp7359 : tmp7351;
  assign tmp7360 = s7 ? tmp7331 : tmp7351;
  assign tmp7357 = s8 ? tmp7358 : tmp7360;
  assign tmp7355 = s9 ? tmp7356 : tmp7357;
  assign tmp7284 = s10 ? tmp7285 : tmp7355;
  assign tmp7364 = s7 ? tmp7306 : tmp7351;
  assign tmp7363 = s8 ? tmp7364 : tmp7360;
  assign tmp7362 = s9 ? tmp7356 : tmp7363;
  assign tmp7361 = s10 ? tmp7285 : tmp7362;
  assign tmp7283 = s11 ? tmp7284 : tmp7361;
  assign tmp7375 = s0 ? tmp7125 : tmp7231;
  assign tmp7374 = s1 ? tmp7125 : tmp7375;
  assign tmp7373 = s2 ? tmp7374 : tmp7292;
  assign tmp7372 = s3 ? tmp7125 : tmp7373;
  assign tmp7371 = s4 ? tmp7125 : tmp7372;
  assign tmp7380 = s1 ? 1 : tmp7230;
  assign tmp7382 = ~(s0 ? 1 : tmp7125);
  assign tmp7381 = s1 ? 1 : tmp7382;
  assign tmp7379 = ~(s2 ? tmp7380 : tmp7381);
  assign tmp7378 = s3 ? tmp7297 : tmp7379;
  assign tmp7385 = s1 ? tmp7228 : tmp7382;
  assign tmp7386 = ~(s1 ? tmp7222 : 1);
  assign tmp7384 = s2 ? tmp7385 : tmp7386;
  assign tmp7388 = s1 ? tmp7125 : tmp7133;
  assign tmp7387 = ~(s2 ? tmp7388 : tmp7232);
  assign tmp7383 = ~(s3 ? tmp7384 : tmp7387);
  assign tmp7377 = s4 ? tmp7378 : tmp7383;
  assign tmp7392 = s1 ? tmp7228 : 0;
  assign tmp7393 = ~(s1 ? tmp7230 : tmp7382);
  assign tmp7391 = s2 ? tmp7392 : tmp7393;
  assign tmp7395 = s1 ? 1 : tmp7329;
  assign tmp7396 = ~(s1 ? tmp7222 : tmp7228);
  assign tmp7394 = s2 ? tmp7395 : tmp7396;
  assign tmp7390 = s3 ? tmp7391 : tmp7394;
  assign tmp7399 = ~(s1 ? tmp7230 : tmp7322);
  assign tmp7398 = s2 ? tmp7325 : tmp7399;
  assign tmp7401 = s1 ? tmp7222 : tmp7329;
  assign tmp7400 = ~(s2 ? tmp7401 : tmp7292);
  assign tmp7397 = s3 ? tmp7398 : tmp7400;
  assign tmp7389 = s4 ? tmp7390 : tmp7397;
  assign tmp7376 = s5 ? tmp7377 : tmp7389;
  assign tmp7370 = s6 ? tmp7371 : tmp7376;
  assign tmp7407 = s1 ? 1 : 0;
  assign tmp7406 = s2 ? tmp7125 : tmp7407;
  assign tmp7409 = s1 ? 1 : tmp7231;
  assign tmp7408 = ~(s2 ? tmp7409 : tmp7381);
  assign tmp7405 = s3 ? tmp7406 : tmp7408;
  assign tmp7411 = s2 ? tmp7385 : 0;
  assign tmp7413 = ~(s1 ? 1 : tmp7125);
  assign tmp7412 = ~(s2 ? tmp7135 : tmp7413);
  assign tmp7410 = ~(s3 ? tmp7411 : tmp7412);
  assign tmp7404 = s4 ? tmp7405 : tmp7410;
  assign tmp7416 = s2 ? tmp7392 : tmp7135;
  assign tmp7418 = ~(s1 ? tmp7125 : 0);
  assign tmp7417 = s2 ? tmp7407 : tmp7418;
  assign tmp7415 = s3 ? tmp7416 : tmp7417;
  assign tmp7420 = s2 ? tmp7135 : tmp7231;
  assign tmp7419 = ~(s3 ? tmp7420 : tmp7298);
  assign tmp7414 = s4 ? tmp7415 : tmp7419;
  assign tmp7403 = s5 ? tmp7404 : tmp7414;
  assign tmp7402 = s6 ? tmp7371 : tmp7403;
  assign tmp7369 = s7 ? tmp7370 : tmp7402;
  assign tmp7425 = s2 ? tmp7374 : tmp7316;
  assign tmp7424 = s3 ? tmp7125 : tmp7425;
  assign tmp7423 = s4 ? tmp7125 : tmp7424;
  assign tmp7430 = ~(s1 ? 1 : 0);
  assign tmp7429 = s2 ? tmp7388 : tmp7430;
  assign tmp7428 = s3 ? tmp7248 : tmp7429;
  assign tmp7432 = s2 ? tmp7392 : 0;
  assign tmp7433 = ~(s2 ? 1 : tmp7232);
  assign tmp7431 = ~(s3 ? tmp7432 : tmp7433);
  assign tmp7427 = s4 ? tmp7428 : tmp7431;
  assign tmp7437 = s1 ? tmp7329 : 0;
  assign tmp7438 = ~(s1 ? tmp7329 : 0);
  assign tmp7436 = s2 ? tmp7437 : tmp7438;
  assign tmp7435 = s3 ? tmp7436 : tmp7394;
  assign tmp7440 = s2 ? tmp7325 : tmp7438;
  assign tmp7439 = s3 ? tmp7440 : tmp7400;
  assign tmp7434 = s4 ? tmp7435 : tmp7439;
  assign tmp7426 = s5 ? tmp7427 : tmp7434;
  assign tmp7422 = s6 ? tmp7423 : tmp7426;
  assign tmp7444 = s2 ? tmp7125 : tmp7135;
  assign tmp7446 = s1 ? tmp7125 : tmp7231;
  assign tmp7445 = s2 ? tmp7446 : tmp7316;
  assign tmp7443 = s3 ? tmp7444 : tmp7445;
  assign tmp7442 = s4 ? tmp7125 : tmp7443;
  assign tmp7451 = s1 ? 1 : tmp7125;
  assign tmp7450 = s2 ? tmp7125 : tmp7451;
  assign tmp7452 = s2 ? tmp7135 : tmp7430;
  assign tmp7449 = s3 ? tmp7450 : tmp7452;
  assign tmp7454 = ~(s2 ? 1 : tmp7413);
  assign tmp7453 = ~(s3 ? tmp7432 : tmp7454);
  assign tmp7448 = s4 ? tmp7449 : tmp7453;
  assign tmp7457 = s2 ? tmp7437 : 1;
  assign tmp7456 = s3 ? tmp7457 : tmp7417;
  assign tmp7459 = s2 ? tmp7135 : 0;
  assign tmp7458 = ~(s3 ? tmp7459 : tmp7298);
  assign tmp7455 = s4 ? tmp7456 : tmp7458;
  assign tmp7447 = s5 ? tmp7448 : tmp7455;
  assign tmp7441 = s6 ? tmp7442 : tmp7447;
  assign tmp7421 = s7 ? tmp7422 : tmp7441;
  assign tmp7368 = s8 ? tmp7369 : tmp7421;
  assign tmp7466 = ~(s2 ? tmp7395 : tmp7407);
  assign tmp7465 = s3 ? tmp7297 : tmp7466;
  assign tmp7464 = s4 ? tmp7465 : tmp7431;
  assign tmp7463 = s5 ? tmp7464 : tmp7434;
  assign tmp7462 = s6 ? tmp7371 : tmp7463;
  assign tmp7470 = s2 ? tmp7446 : tmp7292;
  assign tmp7469 = s3 ? tmp7444 : tmp7470;
  assign tmp7468 = s4 ? tmp7125 : tmp7469;
  assign tmp7473 = s3 ? tmp7406 : tmp7430;
  assign tmp7472 = s4 ? tmp7473 : tmp7453;
  assign tmp7471 = s5 ? tmp7472 : tmp7455;
  assign tmp7467 = s6 ? tmp7468 : tmp7471;
  assign tmp7461 = s7 ? tmp7462 : tmp7467;
  assign tmp7460 = s8 ? tmp7421 : tmp7461;
  assign tmp7367 = s9 ? tmp7368 : tmp7460;
  assign tmp7475 = s8 ? tmp7461 : tmp7462;
  assign tmp7480 = s3 ? tmp7125 : tmp7470;
  assign tmp7479 = s4 ? tmp7125 : tmp7480;
  assign tmp7478 = s6 ? tmp7479 : tmp7403;
  assign tmp7477 = s7 ? tmp7478 : tmp7467;
  assign tmp7481 = s7 ? tmp7441 : tmp7467;
  assign tmp7476 = s8 ? tmp7477 : tmp7481;
  assign tmp7474 = s9 ? tmp7475 : tmp7476;
  assign tmp7366 = s10 ? tmp7367 : tmp7474;
  assign tmp7485 = s7 ? tmp7402 : tmp7467;
  assign tmp7484 = s8 ? tmp7485 : tmp7481;
  assign tmp7483 = s9 ? tmp7475 : tmp7484;
  assign tmp7482 = s10 ? tmp7367 : tmp7483;
  assign tmp7365 = s11 ? tmp7366 : tmp7482;
  assign tmp7282 = s12 ? tmp7283 : tmp7365;
  assign tmp7112 = s13 ? tmp7113 : tmp7282;
  assign tmp7497 = ~(s0 ? tmp7125 : tmp7123);
  assign tmp7496 = s1 ? tmp7146 : tmp7497;
  assign tmp7499 = s1 ? tmp7160 : tmp7146;
  assign tmp7498 = s2 ? tmp7146 : tmp7499;
  assign tmp7495 = s3 ? tmp7496 : tmp7498;
  assign tmp7502 = s1 ? tmp7160 : tmp7322;
  assign tmp7501 = s2 ? tmp7499 : tmp7502;
  assign tmp7504 = s1 ? tmp7125 : tmp7329;
  assign tmp7505 = ~(s1 ? tmp7146 : tmp7148);
  assign tmp7503 = ~(s2 ? tmp7504 : tmp7505);
  assign tmp7500 = s3 ? tmp7501 : tmp7503;
  assign tmp7494 = s4 ? tmp7495 : tmp7500;
  assign tmp7510 = s1 ? 1 : tmp7146;
  assign tmp7509 = s2 ? tmp7146 : tmp7510;
  assign tmp7508 = s3 ? tmp7158 : tmp7509;
  assign tmp7513 = s1 ? tmp7148 : tmp7231;
  assign tmp7515 = ~(s0 ? tmp7146 : 0);
  assign tmp7514 = ~(s1 ? tmp7125 : tmp7515);
  assign tmp7512 = s2 ? tmp7513 : tmp7514;
  assign tmp7516 = s2 ? tmp7496 : 1;
  assign tmp7511 = s3 ? tmp7512 : tmp7516;
  assign tmp7507 = s4 ? tmp7508 : tmp7511;
  assign tmp7521 = s0 ? tmp7146 : 1;
  assign tmp7520 = s1 ? tmp7521 : 1;
  assign tmp7519 = s2 ? tmp7520 : tmp7437;
  assign tmp7523 = ~(s1 ? 1 : tmp7148);
  assign tmp7522 = ~(s2 ? tmp7437 : tmp7523);
  assign tmp7518 = s3 ? tmp7519 : tmp7522;
  assign tmp7526 = s1 ? tmp7148 : 0;
  assign tmp7525 = s2 ? tmp7520 : tmp7526;
  assign tmp7528 = s1 ? 1 : tmp7148;
  assign tmp7529 = s1 ? tmp7148 : 1;
  assign tmp7527 = s2 ? tmp7528 : tmp7529;
  assign tmp7524 = s3 ? tmp7525 : tmp7527;
  assign tmp7517 = s4 ? tmp7518 : tmp7524;
  assign tmp7506 = s5 ? tmp7507 : tmp7517;
  assign tmp7493 = s6 ? tmp7494 : tmp7506;
  assign tmp7534 = s1 ? tmp7160 : tmp7231;
  assign tmp7533 = s2 ? tmp7499 : tmp7534;
  assign tmp7535 = ~(s2 ? tmp7298 : tmp7505);
  assign tmp7532 = s3 ? tmp7533 : tmp7535;
  assign tmp7531 = s4 ? tmp7495 : tmp7532;
  assign tmp7539 = s2 ? tmp7159 : tmp7146;
  assign tmp7538 = s3 ? tmp7539 : tmp7509;
  assign tmp7542 = ~(s1 ? tmp7125 : tmp7123);
  assign tmp7541 = s2 ? tmp7513 : tmp7542;
  assign tmp7540 = s3 ? tmp7541 : tmp7516;
  assign tmp7537 = s4 ? tmp7538 : tmp7540;
  assign tmp7545 = s2 ? tmp7520 : 0;
  assign tmp7546 = s2 ? 1 : tmp7510;
  assign tmp7544 = s3 ? tmp7545 : tmp7546;
  assign tmp7548 = s2 ? 1 : tmp7146;
  assign tmp7547 = s3 ? tmp7548 : tmp7510;
  assign tmp7543 = s4 ? tmp7544 : tmp7547;
  assign tmp7536 = s5 ? tmp7537 : tmp7543;
  assign tmp7530 = s6 ? tmp7531 : tmp7536;
  assign tmp7492 = s7 ? tmp7493 : tmp7530;
  assign tmp7555 = ~(s1 ? tmp7162 : tmp7515);
  assign tmp7554 = s2 ? tmp7159 : tmp7555;
  assign tmp7557 = ~(s1 ? 1 : tmp7146);
  assign tmp7556 = ~(s2 ? tmp7162 : tmp7557);
  assign tmp7553 = s3 ? tmp7554 : tmp7556;
  assign tmp7552 = s4 ? tmp7553 : tmp7511;
  assign tmp7551 = s5 ? tmp7552 : tmp7517;
  assign tmp7550 = s6 ? tmp7494 : tmp7551;
  assign tmp7563 = s1 ? tmp7146 : tmp7160;
  assign tmp7562 = s2 ? tmp7159 : tmp7563;
  assign tmp7561 = s3 ? tmp7562 : tmp7509;
  assign tmp7565 = s2 ? tmp7513 : tmp7146;
  assign tmp7566 = s2 ? tmp7146 : 1;
  assign tmp7564 = s3 ? tmp7565 : tmp7566;
  assign tmp7560 = s4 ? tmp7561 : tmp7564;
  assign tmp7559 = s5 ? tmp7560 : tmp7543;
  assign tmp7558 = s6 ? tmp7531 : tmp7559;
  assign tmp7549 = s7 ? tmp7550 : tmp7558;
  assign tmp7491 = s8 ? tmp7492 : tmp7549;
  assign tmp7571 = s3 ? tmp7125 : tmp7248;
  assign tmp7573 = s2 ? tmp7504 : tmp7316;
  assign tmp7572 = s3 ? tmp7219 : tmp7573;
  assign tmp7570 = s4 ? tmp7571 : tmp7572;
  assign tmp7578 = ~(s1 ? 1 : tmp7231);
  assign tmp7577 = s2 ? tmp7125 : tmp7578;
  assign tmp7576 = s3 ? tmp7240 : tmp7577;
  assign tmp7580 = ~(s2 ? tmp7125 : 0);
  assign tmp7579 = ~(s3 ? tmp7349 : tmp7580);
  assign tmp7575 = s4 ? tmp7576 : tmp7579;
  assign tmp7583 = s2 ? tmp7392 : tmp7438;
  assign tmp7585 = ~(s1 ? 1 : tmp7230);
  assign tmp7584 = s2 ? tmp7437 : tmp7585;
  assign tmp7582 = s3 ? tmp7583 : tmp7584;
  assign tmp7588 = ~(s1 ? tmp7230 : 0);
  assign tmp7587 = s2 ? tmp7392 : tmp7588;
  assign tmp7590 = s1 ? tmp7230 : 1;
  assign tmp7589 = ~(s2 ? tmp7380 : tmp7590);
  assign tmp7586 = s3 ? tmp7587 : tmp7589;
  assign tmp7581 = s4 ? tmp7582 : tmp7586;
  assign tmp7574 = s5 ? tmp7575 : tmp7581;
  assign tmp7569 = s6 ? tmp7570 : tmp7574;
  assign tmp7593 = s3 ? tmp7248 : tmp7334;
  assign tmp7592 = s4 ? tmp7571 : tmp7593;
  assign tmp7597 = s2 ? tmp7241 : tmp7125;
  assign tmp7596 = s3 ? tmp7597 : tmp7577;
  assign tmp7595 = s4 ? tmp7596 : tmp7579;
  assign tmp7600 = s2 ? tmp7392 : 1;
  assign tmp7601 = ~(s2 ? 1 : tmp7409);
  assign tmp7599 = s3 ? tmp7600 : tmp7601;
  assign tmp7603 = s2 ? 1 : tmp7231;
  assign tmp7602 = ~(s3 ? tmp7603 : tmp7409);
  assign tmp7598 = s4 ? tmp7599 : tmp7602;
  assign tmp7594 = s5 ? tmp7595 : tmp7598;
  assign tmp7591 = s6 ? tmp7592 : tmp7594;
  assign tmp7568 = ~(s7 ? tmp7569 : tmp7591);
  assign tmp7567 = s8 ? tmp7549 : tmp7568;
  assign tmp7490 = s9 ? tmp7491 : tmp7567;
  assign tmp7609 = s4 ? tmp7538 : tmp7564;
  assign tmp7608 = s5 ? tmp7609 : tmp7543;
  assign tmp7607 = s6 ? tmp7531 : tmp7608;
  assign tmp7606 = s7 ? tmp7493 : tmp7607;
  assign tmp7605 = s8 ? tmp7606 : tmp7493;
  assign tmp7615 = s3 ? tmp7541 : tmp7566;
  assign tmp7614 = s4 ? tmp7538 : tmp7615;
  assign tmp7613 = s5 ? tmp7614 : tmp7543;
  assign tmp7612 = s6 ? tmp7531 : tmp7613;
  assign tmp7616 = ~(s6 ? tmp7592 : tmp7594);
  assign tmp7611 = s7 ? tmp7612 : tmp7616;
  assign tmp7617 = s7 ? tmp7558 : tmp7607;
  assign tmp7610 = s8 ? tmp7611 : tmp7617;
  assign tmp7604 = s9 ? tmp7605 : tmp7610;
  assign tmp7489 = s10 ? tmp7490 : tmp7604;
  assign tmp7621 = s7 ? tmp7530 : tmp7616;
  assign tmp7620 = s8 ? tmp7621 : tmp7617;
  assign tmp7619 = s9 ? tmp7605 : tmp7620;
  assign tmp7618 = s10 ? tmp7490 : tmp7619;
  assign tmp7488 = s11 ? tmp7489 : tmp7618;
  assign tmp7487 = s12 ? 1 : tmp7488;
  assign tmp7632 = s1 ? tmp7228 : tmp7125;
  assign tmp7631 = s2 ? tmp7125 : tmp7632;
  assign tmp7630 = s3 ? tmp7125 : tmp7631;
  assign tmp7634 = s2 ? tmp7125 : tmp7228;
  assign tmp7636 = s1 ? tmp7125 : tmp7330;
  assign tmp7635 = s2 ? tmp7636 : tmp7221;
  assign tmp7633 = s3 ? tmp7634 : tmp7635;
  assign tmp7629 = s4 ? tmp7630 : tmp7633;
  assign tmp7641 = ~(s1 ? tmp7230 : tmp7301);
  assign tmp7640 = s2 ? tmp7292 : tmp7641;
  assign tmp7642 = ~(s2 ? tmp7230 : tmp7413);
  assign tmp7639 = s3 ? tmp7640 : tmp7642;
  assign tmp7644 = s2 ? tmp7242 : tmp7125;
  assign tmp7643 = s3 ? tmp7644 : tmp7256;
  assign tmp7638 = s4 ? tmp7639 : tmp7643;
  assign tmp7637 = s5 ? tmp7638 : tmp7238;
  assign tmp7628 = s6 ? tmp7629 : tmp7637;
  assign tmp7647 = s3 ? tmp7631 : tmp7220;
  assign tmp7646 = s4 ? tmp7630 : tmp7647;
  assign tmp7651 = s2 ? tmp7632 : tmp7227;
  assign tmp7650 = s3 ? tmp7651 : tmp7450;
  assign tmp7649 = s4 ? tmp7650 : tmp7643;
  assign tmp7654 = s2 ? tmp7241 : 1;
  assign tmp7653 = s3 ? tmp7597 : tmp7654;
  assign tmp7652 = s4 ? tmp7653 : tmp7260;
  assign tmp7648 = s5 ? tmp7649 : tmp7652;
  assign tmp7645 = s6 ? tmp7646 : tmp7648;
  assign tmp7627 = s7 ? tmp7628 : tmp7645;
  assign tmp7660 = ~(l3 ? 1 : 0);
  assign tmp7659 = l1 ? 1 : tmp7660;
  assign tmp7663 = s0 ? tmp7659 : tmp7660;
  assign tmp7662 = s1 ? tmp7663 : tmp7659;
  assign tmp7661 = s2 ? tmp7659 : tmp7662;
  assign tmp7658 = s3 ? tmp7659 : tmp7661;
  assign tmp7667 = s0 ? tmp7659 : tmp7125;
  assign tmp7666 = s1 ? tmp7667 : tmp7659;
  assign tmp7668 = s0 ? tmp7659 : 0;
  assign tmp7665 = s2 ? tmp7666 : tmp7668;
  assign tmp7670 = s1 ? tmp7659 : tmp7330;
  assign tmp7672 = s0 ? 1 : tmp7659;
  assign tmp7671 = s1 ? tmp7659 : tmp7672;
  assign tmp7669 = s2 ? tmp7670 : tmp7671;
  assign tmp7664 = s3 ? tmp7665 : tmp7669;
  assign tmp7657 = s4 ? tmp7658 : tmp7664;
  assign tmp7679 = ~(l1 ? 1 : tmp7660);
  assign tmp7678 = ~(s0 ? 1 : tmp7679);
  assign tmp7677 = s1 ? tmp7668 : tmp7678;
  assign tmp7681 = s0 ? 1 : tmp7679;
  assign tmp7682 = ~(s0 ? tmp7659 : tmp7660);
  assign tmp7680 = ~(s1 ? tmp7681 : tmp7682);
  assign tmp7676 = s2 ? tmp7677 : tmp7680;
  assign tmp7685 = l3 ? 1 : 0;
  assign tmp7684 = s0 ? tmp7685 : tmp7679;
  assign tmp7686 = ~(s1 ? 1 : tmp7659);
  assign tmp7683 = ~(s2 ? tmp7684 : tmp7686);
  assign tmp7675 = s3 ? tmp7676 : tmp7683;
  assign tmp7689 = s1 ? tmp7672 : tmp7133;
  assign tmp7690 = s1 ? tmp7133 : tmp7667;
  assign tmp7688 = s2 ? tmp7689 : tmp7690;
  assign tmp7692 = s1 ? tmp7659 : 1;
  assign tmp7691 = s2 ? tmp7692 : 1;
  assign tmp7687 = s3 ? tmp7688 : tmp7691;
  assign tmp7674 = s4 ? tmp7675 : tmp7687;
  assign tmp7697 = s0 ? tmp7659 : 1;
  assign tmp7696 = s1 ? tmp7697 : 1;
  assign tmp7695 = s2 ? tmp7696 : tmp7672;
  assign tmp7694 = s3 ? tmp7695 : 1;
  assign tmp7700 = s1 ? tmp7672 : tmp7697;
  assign tmp7699 = s2 ? 1 : tmp7700;
  assign tmp7698 = s3 ? tmp7699 : 1;
  assign tmp7693 = s4 ? tmp7694 : tmp7698;
  assign tmp7673 = s5 ? tmp7674 : tmp7693;
  assign tmp7656 = s6 ? tmp7657 : tmp7673;
  assign tmp7705 = s1 ? tmp7668 : tmp7659;
  assign tmp7704 = s2 ? tmp7666 : tmp7705;
  assign tmp7706 = s2 ? tmp7692 : tmp7671;
  assign tmp7703 = s3 ? tmp7704 : tmp7706;
  assign tmp7702 = s4 ? tmp7658 : tmp7703;
  assign tmp7711 = s1 ? tmp7659 : tmp7663;
  assign tmp7710 = s2 ? tmp7705 : tmp7711;
  assign tmp7713 = s1 ? 1 : tmp7659;
  assign tmp7712 = s2 ? tmp7659 : tmp7713;
  assign tmp7709 = s3 ? tmp7710 : tmp7712;
  assign tmp7715 = s2 ? tmp7689 : tmp7659;
  assign tmp7714 = s3 ? tmp7715 : tmp7691;
  assign tmp7708 = s4 ? tmp7709 : tmp7714;
  assign tmp7718 = s2 ? tmp7696 : tmp7692;
  assign tmp7717 = s3 ? tmp7718 : tmp7654;
  assign tmp7721 = s1 ? tmp7659 : tmp7125;
  assign tmp7720 = s2 ? 1 : tmp7721;
  assign tmp7719 = s3 ? tmp7720 : 1;
  assign tmp7716 = s4 ? tmp7717 : tmp7719;
  assign tmp7707 = s5 ? tmp7708 : tmp7716;
  assign tmp7701 = s6 ? tmp7702 : tmp7707;
  assign tmp7655 = s7 ? tmp7656 : tmp7701;
  assign tmp7626 = s8 ? tmp7627 : tmp7655;
  assign tmp7725 = s5 ? tmp7649 : tmp7257;
  assign tmp7724 = s6 ? tmp7646 : tmp7725;
  assign tmp7723 = s7 ? tmp7628 : tmp7724;
  assign tmp7722 = s8 ? tmp7655 : tmp7723;
  assign tmp7625 = s9 ? tmp7626 : tmp7722;
  assign tmp7732 = s3 ? tmp7259 : tmp7654;
  assign tmp7731 = s4 ? tmp7732 : tmp7260;
  assign tmp7730 = s5 ? tmp7649 : tmp7731;
  assign tmp7729 = s6 ? tmp7646 : tmp7730;
  assign tmp7728 = s7 ? tmp7628 : tmp7729;
  assign tmp7727 = s8 ? tmp7728 : tmp7628;
  assign tmp7734 = s7 ? tmp7645 : tmp7724;
  assign tmp7740 = s2 ? 1 : tmp7659;
  assign tmp7739 = s3 ? tmp7740 : 1;
  assign tmp7738 = s4 ? tmp7717 : tmp7739;
  assign tmp7737 = s5 ? tmp7708 : tmp7738;
  assign tmp7736 = s6 ? tmp7702 : tmp7737;
  assign tmp7735 = s7 ? tmp7736 : tmp7729;
  assign tmp7733 = s8 ? tmp7734 : tmp7735;
  assign tmp7726 = s9 ? tmp7727 : tmp7733;
  assign tmp7624 = s10 ? tmp7625 : tmp7726;
  assign tmp7744 = s7 ? tmp7701 : tmp7729;
  assign tmp7743 = s8 ? tmp7734 : tmp7744;
  assign tmp7742 = s9 ? tmp7727 : tmp7743;
  assign tmp7741 = s10 ? tmp7625 : tmp7742;
  assign tmp7623 = s11 ? tmp7624 : tmp7741;
  assign tmp7753 = s3 ? 1 : tmp7654;
  assign tmp7752 = s4 ? tmp7753 : tmp7260;
  assign tmp7751 = s5 ? 1 : tmp7752;
  assign tmp7750 = s6 ? 1 : tmp7751;
  assign tmp7749 = s7 ? 1 : tmp7750;
  assign tmp7759 = s2 ? 1 : tmp7451;
  assign tmp7758 = s3 ? tmp7759 : 1;
  assign tmp7757 = s4 ? tmp7753 : tmp7758;
  assign tmp7756 = s5 ? 1 : tmp7757;
  assign tmp7755 = s6 ? 1 : tmp7756;
  assign tmp7754 = s7 ? 1 : tmp7755;
  assign tmp7748 = s8 ? tmp7749 : tmp7754;
  assign tmp7760 = s8 ? tmp7754 : 1;
  assign tmp7747 = s9 ? tmp7748 : tmp7760;
  assign tmp7762 = s8 ? tmp7749 : 1;
  assign tmp7767 = s4 ? tmp7753 : 1;
  assign tmp7766 = s5 ? 1 : tmp7767;
  assign tmp7765 = s6 ? 1 : tmp7766;
  assign tmp7764 = s7 ? tmp7765 : 1;
  assign tmp7763 = s8 ? tmp7764 : tmp7765;
  assign tmp7761 = s9 ? tmp7762 : tmp7763;
  assign tmp7746 = s10 ? tmp7747 : tmp7761;
  assign tmp7771 = s7 ? tmp7750 : 1;
  assign tmp7772 = s7 ? tmp7755 : tmp7750;
  assign tmp7770 = s8 ? tmp7771 : tmp7772;
  assign tmp7769 = s9 ? tmp7762 : tmp7770;
  assign tmp7768 = s10 ? tmp7747 : tmp7769;
  assign tmp7745 = s11 ? tmp7746 : tmp7768;
  assign tmp7622 = ~(s12 ? tmp7623 : tmp7745);
  assign tmp7486 = ~(s13 ? tmp7487 : tmp7622);
  assign tmp7111 = s14 ? tmp7112 : tmp7486;
  assign tmp7782 = s2 ? tmp7222 : tmp7451;
  assign tmp7781 = s3 ? 1 : tmp7782;
  assign tmp7784 = s2 ? tmp7451 : 1;
  assign tmp7786 = s1 ? 1 : tmp7222;
  assign tmp7785 = s2 ? tmp7786 : tmp7125;
  assign tmp7783 = s3 ? tmp7784 : tmp7785;
  assign tmp7780 = s4 ? tmp7781 : tmp7783;
  assign tmp7790 = s2 ? 1 : tmp7253;
  assign tmp7789 = s3 ? tmp7790 : tmp7785;
  assign tmp7791 = s3 ? tmp7256 : tmp7785;
  assign tmp7788 = s4 ? tmp7789 : tmp7791;
  assign tmp7794 = s2 ? tmp7388 : 1;
  assign tmp7795 = s2 ? tmp7786 : tmp7241;
  assign tmp7793 = s3 ? tmp7794 : tmp7795;
  assign tmp7796 = s3 ? tmp7795 : tmp7794;
  assign tmp7792 = s4 ? tmp7793 : tmp7796;
  assign tmp7787 = s5 ? tmp7788 : tmp7792;
  assign tmp7779 = s6 ? tmp7780 : tmp7787;
  assign tmp7800 = s2 ? tmp7451 : tmp7125;
  assign tmp7799 = s3 ? tmp7784 : tmp7800;
  assign tmp7798 = s4 ? tmp7781 : tmp7799;
  assign tmp7803 = s3 ? tmp7790 : tmp7800;
  assign tmp7804 = s3 ? tmp7256 : tmp7800;
  assign tmp7802 = s4 ? tmp7803 : tmp7804;
  assign tmp7806 = s3 ? tmp7794 : tmp7784;
  assign tmp7808 = s2 ? tmp7451 : tmp7133;
  assign tmp7807 = s3 ? tmp7808 : tmp7135;
  assign tmp7805 = s4 ? tmp7806 : tmp7807;
  assign tmp7801 = s5 ? tmp7802 : tmp7805;
  assign tmp7797 = s6 ? tmp7798 : tmp7801;
  assign tmp7778 = s7 ? tmp7779 : tmp7797;
  assign tmp7810 = s8 ? tmp7778 : tmp7779;
  assign tmp7814 = s3 ? tmp7784 : tmp7135;
  assign tmp7813 = s4 ? tmp7806 : tmp7814;
  assign tmp7812 = s5 ? tmp7802 : tmp7813;
  assign tmp7811 = s6 ? tmp7798 : tmp7812;
  assign tmp7809 = s9 ? tmp7810 : tmp7811;
  assign tmp7777 = s10 ? tmp7778 : tmp7809;
  assign tmp7816 = s9 ? tmp7810 : tmp7797;
  assign tmp7815 = s10 ? tmp7778 : tmp7816;
  assign tmp7776 = s11 ? tmp7777 : tmp7815;
  assign tmp7821 = s3 ? tmp7298 : tmp7125;
  assign tmp7820 = s4 ? tmp7821 : tmp7125;
  assign tmp7825 = s2 ? 1 : tmp7409;
  assign tmp7824 = s3 ? tmp7825 : tmp7231;
  assign tmp7823 = s4 ? tmp7824 : tmp7231;
  assign tmp7828 = ~(s2 ? 1 : tmp7350);
  assign tmp7827 = s3 ? tmp7125 : tmp7828;
  assign tmp7830 = ~(s1 ? tmp7228 : 0);
  assign tmp7829 = ~(s2 ? tmp7380 : tmp7830);
  assign tmp7826 = ~(s4 ? tmp7827 : tmp7829);
  assign tmp7822 = ~(s5 ? tmp7823 : tmp7826);
  assign tmp7819 = s6 ? tmp7820 : tmp7822;
  assign tmp7835 = ~(s2 ? 1 : tmp7231);
  assign tmp7834 = s3 ? tmp7125 : tmp7835;
  assign tmp7836 = ~(s2 ? tmp7409 : 1);
  assign tmp7833 = ~(s4 ? tmp7834 : tmp7836);
  assign tmp7832 = ~(s5 ? tmp7823 : tmp7833);
  assign tmp7831 = s6 ? tmp7820 : tmp7832;
  assign tmp7818 = s7 ? tmp7819 : tmp7831;
  assign tmp7838 = s8 ? tmp7818 : tmp7819;
  assign tmp7837 = s9 ? tmp7838 : tmp7831;
  assign tmp7817 = s10 ? tmp7818 : tmp7837;
  assign tmp7775 = s12 ? tmp7776 : tmp7817;
  assign tmp7845 = ~(s2 ? tmp7350 : tmp7305);
  assign tmp7844 = s3 ? tmp7316 : tmp7845;
  assign tmp7847 = s2 ? tmp7409 : tmp7830;
  assign tmp7848 = s2 ? tmp7380 : tmp7231;
  assign tmp7846 = ~(s3 ? tmp7847 : tmp7848);
  assign tmp7843 = s4 ? tmp7844 : tmp7846;
  assign tmp7852 = s2 ? tmp7392 : tmp7641;
  assign tmp7853 = ~(s2 ? tmp7230 : tmp7231);
  assign tmp7851 = s3 ? tmp7852 : tmp7853;
  assign tmp7855 = s2 ? tmp7298 : 0;
  assign tmp7854 = s3 ? tmp7855 : tmp7853;
  assign tmp7850 = s4 ? tmp7851 : tmp7854;
  assign tmp7858 = s2 ? tmp7221 : tmp7392;
  assign tmp7860 = ~(s1 ? tmp7125 : tmp7228);
  assign tmp7859 = ~(s2 ? tmp7380 : tmp7860);
  assign tmp7857 = s3 ? tmp7858 : tmp7859;
  assign tmp7863 = ~(s1 ? tmp7222 : 0);
  assign tmp7862 = s2 ? tmp7350 : tmp7863;
  assign tmp7864 = ~(s2 ? tmp7125 : tmp7292);
  assign tmp7861 = ~(s3 ? tmp7862 : tmp7864);
  assign tmp7856 = s4 ? tmp7857 : tmp7861;
  assign tmp7849 = s5 ? tmp7850 : tmp7856;
  assign tmp7842 = s6 ? tmp7843 : tmp7849;
  assign tmp7868 = s2 ? tmp7409 : tmp7231;
  assign tmp7867 = ~(s3 ? tmp7847 : tmp7868);
  assign tmp7866 = s4 ? tmp7844 : tmp7867;
  assign tmp7872 = s2 ? tmp7392 : tmp7227;
  assign tmp7871 = s3 ? tmp7872 : tmp7125;
  assign tmp7870 = s4 ? tmp7871 : tmp7854;
  assign tmp7875 = s2 ? tmp7125 : 0;
  assign tmp7876 = ~(s2 ? tmp7409 : tmp7860);
  assign tmp7874 = s3 ? tmp7875 : tmp7876;
  assign tmp7873 = s4 ? tmp7874 : tmp7125;
  assign tmp7869 = s5 ? tmp7870 : tmp7873;
  assign tmp7865 = s6 ? tmp7866 : tmp7869;
  assign tmp7841 = s7 ? tmp7842 : tmp7865;
  assign tmp7878 = s8 ? tmp7841 : tmp7842;
  assign tmp7877 = s9 ? tmp7878 : tmp7865;
  assign tmp7840 = s10 ? tmp7841 : tmp7877;
  assign tmp7883 = s3 ? tmp7135 : tmp7782;
  assign tmp7885 = s2 ? tmp7451 : tmp7241;
  assign tmp7884 = s3 ? tmp7885 : tmp7785;
  assign tmp7882 = s4 ? tmp7883 : tmp7884;
  assign tmp7890 = ~(s1 ? 1 : tmp7301);
  assign tmp7889 = s2 ? tmp7222 : tmp7890;
  assign tmp7888 = s3 ? tmp7256 : tmp7889;
  assign tmp7887 = s4 ? tmp7789 : tmp7888;
  assign tmp7893 = s2 ? tmp7242 : tmp7388;
  assign tmp7892 = s3 ? tmp7237 : tmp7893;
  assign tmp7895 = s2 ? tmp7242 : tmp7133;
  assign tmp7894 = s3 ? tmp7885 : tmp7895;
  assign tmp7891 = s4 ? tmp7892 : tmp7894;
  assign tmp7886 = s5 ? tmp7887 : tmp7891;
  assign tmp7881 = s6 ? tmp7882 : tmp7886;
  assign tmp7898 = s3 ? tmp7885 : tmp7800;
  assign tmp7897 = s4 ? tmp7883 : tmp7898;
  assign tmp7902 = s2 ? tmp7242 : tmp7578;
  assign tmp7901 = s3 ? tmp7256 : tmp7902;
  assign tmp7900 = s4 ? tmp7803 : tmp7901;
  assign tmp7904 = s3 ? tmp7256 : tmp7444;
  assign tmp7905 = s3 ? tmp7237 : tmp7125;
  assign tmp7903 = s4 ? tmp7904 : tmp7905;
  assign tmp7899 = s5 ? tmp7900 : tmp7903;
  assign tmp7896 = s6 ? tmp7897 : tmp7899;
  assign tmp7880 = s7 ? tmp7881 : tmp7896;
  assign tmp7907 = s8 ? tmp7880 : tmp7881;
  assign tmp7906 = s9 ? tmp7907 : tmp7896;
  assign tmp7879 = s10 ? tmp7880 : tmp7906;
  assign tmp7839 = s12 ? tmp7840 : tmp7879;
  assign tmp7774 = s13 ? tmp7775 : tmp7839;
  assign tmp7918 = s2 ? tmp7236 : tmp7133;
  assign tmp7919 = s2 ? tmp7504 : tmp7125;
  assign tmp7917 = s3 ? tmp7918 : tmp7919;
  assign tmp7916 = s4 ? tmp7571 : tmp7917;
  assign tmp7922 = s3 ? tmp7240 : tmp7631;
  assign tmp7925 = ~(s1 ? tmp7125 : tmp7133);
  assign tmp7924 = s2 ? tmp7350 : tmp7925;
  assign tmp7923 = ~(s3 ? tmp7924 : tmp7580);
  assign tmp7921 = s4 ? tmp7922 : tmp7923;
  assign tmp7928 = s2 ? tmp7292 : tmp7241;
  assign tmp7927 = s3 ? tmp7928 : tmp7584;
  assign tmp7930 = s2 ? tmp7125 : tmp7588;
  assign tmp7931 = s2 ? tmp7316 : tmp7293;
  assign tmp7929 = s3 ? tmp7930 : tmp7931;
  assign tmp7926 = s4 ? tmp7927 : tmp7929;
  assign tmp7920 = s5 ? tmp7921 : tmp7926;
  assign tmp7915 = s6 ? tmp7916 : tmp7920;
  assign tmp7935 = s2 ? tmp7298 : tmp7125;
  assign tmp7934 = s3 ? tmp7236 : tmp7935;
  assign tmp7933 = s4 ? tmp7571 : tmp7934;
  assign tmp7938 = s3 ? tmp7597 : tmp7631;
  assign tmp7937 = s4 ? tmp7938 : tmp7579;
  assign tmp7941 = s2 ? tmp7632 : 1;
  assign tmp7942 = s2 ? tmp7392 : tmp7578;
  assign tmp7940 = s3 ? tmp7941 : tmp7942;
  assign tmp7939 = s4 ? tmp7940 : tmp7125;
  assign tmp7936 = s5 ? tmp7937 : tmp7939;
  assign tmp7932 = s6 ? tmp7933 : tmp7936;
  assign tmp7914 = s7 ? tmp7915 : tmp7932;
  assign tmp7950 = l4 ? 1 : 0;
  assign tmp7949 = l2 ? tmp7950 : 0;
  assign tmp7948 = l1 ? 1 : tmp7949;
  assign tmp7952 = l1 ? 1 : tmp7950;
  assign tmp7951 = s0 ? tmp7952 : tmp7948;
  assign tmp7947 = s1 ? tmp7948 : tmp7951;
  assign tmp7955 = s0 ? tmp7952 : 1;
  assign tmp7954 = s1 ? tmp7955 : tmp7948;
  assign tmp7953 = s2 ? tmp7948 : tmp7954;
  assign tmp7946 = s3 ? tmp7947 : tmp7953;
  assign tmp7959 = s0 ? tmp7948 : 1;
  assign tmp7958 = s1 ? tmp7959 : tmp7948;
  assign tmp7960 = s1 ? tmp7959 : tmp7955;
  assign tmp7957 = s2 ? tmp7958 : tmp7960;
  assign tmp7962 = s1 ? tmp7952 : tmp7329;
  assign tmp7961 = s2 ? tmp7962 : tmp7948;
  assign tmp7956 = s3 ? tmp7957 : tmp7961;
  assign tmp7945 = s4 ? tmp7946 : tmp7956;
  assign tmp7967 = s1 ? tmp7959 : 1;
  assign tmp7969 = s0 ? 1 : tmp7948;
  assign tmp7968 = s1 ? tmp7969 : tmp7959;
  assign tmp7966 = s2 ? tmp7967 : tmp7968;
  assign tmp7972 = s0 ? tmp7948 : 0;
  assign tmp7971 = s1 ? tmp7972 : tmp7948;
  assign tmp7970 = s2 ? tmp7969 : tmp7971;
  assign tmp7965 = s3 ? tmp7966 : tmp7970;
  assign tmp7977 = ~(l1 ? 1 : tmp7949);
  assign tmp7976 = s0 ? 1 : tmp7977;
  assign tmp7978 = ~(s0 ? 1 : tmp7952);
  assign tmp7975 = s1 ? tmp7976 : tmp7978;
  assign tmp7980 = s0 ? 1 : tmp7952;
  assign tmp7979 = ~(s1 ? tmp7980 : tmp7959);
  assign tmp7974 = s2 ? tmp7975 : tmp7979;
  assign tmp7983 = s0 ? tmp7952 : tmp7125;
  assign tmp7982 = s1 ? tmp7948 : tmp7983;
  assign tmp7981 = ~(s2 ? tmp7982 : 0);
  assign tmp7973 = ~(s3 ? tmp7974 : tmp7981);
  assign tmp7964 = s4 ? tmp7965 : tmp7973;
  assign tmp7989 = ~(l1 ? 1 : tmp7950);
  assign tmp7988 = ~(s0 ? 1 : tmp7989);
  assign tmp7987 = s1 ? tmp7972 : tmp7988;
  assign tmp7990 = s1 ? tmp7955 : 1;
  assign tmp7986 = s2 ? tmp7987 : tmp7990;
  assign tmp7985 = s3 ? tmp7986 : tmp7584;
  assign tmp7994 = s0 ? tmp7125 : tmp7948;
  assign tmp7993 = s1 ? tmp7125 : tmp7994;
  assign tmp7995 = ~(s1 ? tmp7976 : 0);
  assign tmp7992 = s2 ? tmp7993 : tmp7995;
  assign tmp7997 = s1 ? tmp7983 : tmp7293;
  assign tmp7996 = s2 ? tmp7997 : tmp7293;
  assign tmp7991 = s3 ? tmp7992 : tmp7996;
  assign tmp7984 = s4 ? tmp7985 : tmp7991;
  assign tmp7963 = s5 ? tmp7964 : tmp7984;
  assign tmp7944 = s6 ? tmp7945 : tmp7963;
  assign tmp8002 = s1 ? tmp7959 : tmp7952;
  assign tmp8001 = s2 ? tmp7958 : tmp8002;
  assign tmp8004 = s1 ? tmp7952 : 0;
  assign tmp8003 = s2 ? tmp8004 : tmp7948;
  assign tmp8000 = s3 ? tmp8001 : tmp8003;
  assign tmp7999 = s4 ? tmp7946 : tmp8000;
  assign tmp8009 = s1 ? tmp7948 : tmp7959;
  assign tmp8008 = s2 ? tmp7967 : tmp8009;
  assign tmp8010 = s2 ? tmp7948 : tmp7971;
  assign tmp8007 = s3 ? tmp8008 : tmp8010;
  assign tmp8012 = s2 ? tmp7975 : tmp7977;
  assign tmp8014 = s1 ? tmp7948 : tmp7125;
  assign tmp8013 = ~(s2 ? tmp8014 : 0);
  assign tmp8011 = ~(s3 ? tmp8012 : tmp8013);
  assign tmp8006 = s4 ? tmp8007 : tmp8011;
  assign tmp8018 = s1 ? tmp7972 : tmp7952;
  assign tmp8017 = s2 ? tmp8018 : 1;
  assign tmp8016 = s3 ? tmp8017 : tmp7942;
  assign tmp8021 = s1 ? tmp7125 : tmp7948;
  assign tmp8020 = s2 ? tmp8021 : tmp8014;
  assign tmp8019 = s3 ? tmp8020 : tmp7125;
  assign tmp8015 = s4 ? tmp8016 : tmp8019;
  assign tmp8005 = s5 ? tmp8006 : tmp8015;
  assign tmp7998 = s6 ? tmp7999 : tmp8005;
  assign tmp7943 = s7 ? tmp7944 : tmp7998;
  assign tmp7913 = s8 ? tmp7914 : tmp7943;
  assign tmp8028 = s2 ? tmp7437 : tmp7578;
  assign tmp8027 = s3 ? tmp7941 : tmp8028;
  assign tmp8026 = s4 ? tmp8027 : tmp7125;
  assign tmp8025 = s5 ? tmp7937 : tmp8026;
  assign tmp8024 = s6 ? tmp7933 : tmp8025;
  assign tmp8023 = s7 ? tmp7915 : tmp8024;
  assign tmp8022 = s8 ? tmp7943 : tmp8023;
  assign tmp7912 = s9 ? tmp7913 : tmp8022;
  assign tmp8030 = s8 ? tmp7914 : tmp7915;
  assign tmp8032 = s7 ? tmp7932 : tmp8024;
  assign tmp8038 = s2 ? tmp8021 : tmp7948;
  assign tmp8037 = s3 ? tmp8038 : tmp7125;
  assign tmp8036 = s4 ? tmp8016 : tmp8037;
  assign tmp8035 = s5 ? tmp8006 : tmp8036;
  assign tmp8034 = s6 ? tmp7999 : tmp8035;
  assign tmp8033 = s7 ? tmp8034 : tmp7932;
  assign tmp8031 = s8 ? tmp8032 : tmp8033;
  assign tmp8029 = s9 ? tmp8030 : tmp8031;
  assign tmp7911 = s10 ? tmp7912 : tmp8029;
  assign tmp8042 = s7 ? tmp7998 : tmp7932;
  assign tmp8041 = s8 ? tmp8032 : tmp8042;
  assign tmp8040 = s9 ? tmp8030 : tmp8041;
  assign tmp8039 = s10 ? tmp7912 : tmp8040;
  assign tmp7910 = s11 ? tmp7911 : tmp8039;
  assign tmp8052 = ~(l1 ? 1 : tmp7123);
  assign tmp8051 = s0 ? 1 : tmp8052;
  assign tmp8054 = s1 ? tmp7138 : tmp7122;
  assign tmp8056 = s0 ? tmp7122 : 0;
  assign tmp8055 = s1 ? tmp8056 : tmp7122;
  assign tmp8053 = ~(s2 ? tmp8054 : tmp8055);
  assign tmp8050 = s3 ? tmp8051 : tmp8053;
  assign tmp8060 = s0 ? tmp7122 : tmp7231;
  assign tmp8059 = s1 ? tmp8060 : tmp7122;
  assign tmp8061 = s1 ? tmp8056 : 0;
  assign tmp8058 = s2 ? tmp8059 : tmp8061;
  assign tmp8063 = ~(s1 ? tmp7122 : tmp7124);
  assign tmp8062 = ~(s2 ? tmp7380 : tmp8063);
  assign tmp8057 = ~(s3 ? tmp8058 : tmp8062);
  assign tmp8049 = s4 ? tmp8050 : tmp8057;
  assign tmp8068 = s1 ? tmp7132 : 1;
  assign tmp8069 = s1 ? tmp7138 : tmp8056;
  assign tmp8067 = s2 ? tmp8068 : tmp8069;
  assign tmp8071 = ~(s1 ? tmp7133 : tmp7122);
  assign tmp8070 = ~(s2 ? tmp8051 : tmp8071);
  assign tmp8066 = s3 ? tmp8067 : tmp8070;
  assign tmp8074 = s1 ? tmp7124 : tmp7322;
  assign tmp8076 = ~(s0 ? tmp7122 : tmp7231);
  assign tmp8075 = ~(s1 ? tmp7133 : tmp8076);
  assign tmp8073 = s2 ? tmp8074 : tmp8075;
  assign tmp8079 = ~(s0 ? 1 : tmp8052);
  assign tmp8078 = s1 ? tmp7122 : tmp8079;
  assign tmp8077 = s2 ? tmp8078 : tmp7253;
  assign tmp8072 = s3 ? tmp8073 : tmp8077;
  assign tmp8065 = s4 ? tmp8066 : tmp8072;
  assign tmp8083 = s1 ? tmp7132 : tmp7222;
  assign tmp8082 = s2 ? tmp8083 : tmp7241;
  assign tmp8085 = s1 ? tmp7125 : tmp7124;
  assign tmp8084 = s2 ? 1 : tmp8085;
  assign tmp8081 = s3 ? tmp8082 : tmp8084;
  assign tmp8088 = s1 ? tmp7138 : 1;
  assign tmp8087 = s2 ? tmp7170 : tmp8088;
  assign tmp8090 = s1 ? tmp7125 : tmp7138;
  assign tmp8091 = s1 ? tmp7124 : 1;
  assign tmp8089 = s2 ? tmp8090 : tmp8091;
  assign tmp8086 = s3 ? tmp8087 : tmp8089;
  assign tmp8080 = s4 ? tmp8081 : tmp8086;
  assign tmp8064 = ~(s5 ? tmp8065 : tmp8080);
  assign tmp8048 = s6 ? tmp8049 : tmp8064;
  assign tmp8095 = ~(s2 ? tmp7409 : tmp8063);
  assign tmp8094 = ~(s3 ? tmp8058 : tmp8095);
  assign tmp8093 = s4 ? tmp8050 : tmp8094;
  assign tmp8100 = s1 ? tmp7122 : tmp8056;
  assign tmp8099 = s2 ? tmp8068 : tmp8100;
  assign tmp8102 = s1 ? tmp7133 : tmp7122;
  assign tmp8101 = s2 ? tmp7122 : tmp8102;
  assign tmp8098 = s3 ? tmp8099 : tmp8101;
  assign tmp8104 = s2 ? tmp8074 : tmp7122;
  assign tmp8105 = s2 ? tmp7122 : tmp7451;
  assign tmp8103 = s3 ? tmp8104 : tmp8105;
  assign tmp8097 = s4 ? tmp8098 : tmp8103;
  assign tmp8108 = s2 ? tmp7170 : tmp7241;
  assign tmp8109 = s2 ? 1 : tmp7276;
  assign tmp8107 = s3 ? tmp8108 : tmp8109;
  assign tmp8111 = s2 ? tmp7125 : tmp7122;
  assign tmp8110 = s3 ? tmp8111 : tmp7276;
  assign tmp8106 = s4 ? tmp8107 : tmp8110;
  assign tmp8096 = ~(s5 ? tmp8097 : tmp8106);
  assign tmp8092 = s6 ? tmp8093 : tmp8096;
  assign tmp8047 = s7 ? tmp8048 : tmp8092;
  assign tmp8117 = s0 ? tmp7950 : tmp7952;
  assign tmp8116 = s1 ? tmp7952 : tmp8117;
  assign tmp8119 = s1 ? tmp7980 : tmp7952;
  assign tmp8120 = s1 ? tmp7955 : tmp7952;
  assign tmp8118 = s2 ? tmp8119 : tmp8120;
  assign tmp8115 = s3 ? tmp8116 : tmp8118;
  assign tmp8124 = s0 ? tmp7952 : 0;
  assign tmp8125 = s0 ? tmp7950 : 0;
  assign tmp8123 = s1 ? tmp8124 : tmp8125;
  assign tmp8122 = s2 ? tmp8120 : tmp8123;
  assign tmp8127 = s1 ? tmp7950 : tmp7293;
  assign tmp8126 = s2 ? tmp8127 : tmp7952;
  assign tmp8121 = s3 ? tmp8122 : tmp8126;
  assign tmp8114 = s4 ? tmp8115 : tmp8121;
  assign tmp8132 = s1 ? tmp7980 : tmp7955;
  assign tmp8131 = s2 ? tmp7990 : tmp8132;
  assign tmp8133 = s2 ? tmp7980 : tmp8120;
  assign tmp8130 = s3 ? tmp8131 : tmp8133;
  assign tmp8137 = s0 ? tmp7125 : tmp7952;
  assign tmp8138 = s0 ? 1 : tmp7950;
  assign tmp8136 = s1 ? tmp8137 : tmp8138;
  assign tmp8139 = s1 ? tmp8138 : tmp7955;
  assign tmp8135 = s2 ? tmp8136 : tmp8139;
  assign tmp8142 = s0 ? tmp7950 : tmp7122;
  assign tmp8141 = s1 ? tmp7952 : tmp8142;
  assign tmp8140 = s2 ? tmp8141 : tmp7253;
  assign tmp8134 = s3 ? tmp8135 : tmp8140;
  assign tmp8129 = s4 ? tmp8130 : tmp8134;
  assign tmp8146 = s1 ? tmp7955 : tmp7980;
  assign tmp8145 = s2 ? tmp8146 : tmp7990;
  assign tmp8144 = s3 ? tmp8145 : tmp8084;
  assign tmp8149 = s1 ? tmp7132 : tmp7980;
  assign tmp8150 = s1 ? tmp7980 : 1;
  assign tmp8148 = s2 ? tmp8149 : tmp8150;
  assign tmp8152 = s1 ? tmp7955 : tmp7138;
  assign tmp8151 = s2 ? tmp8152 : tmp8091;
  assign tmp8147 = s3 ? tmp8148 : tmp8151;
  assign tmp8143 = s4 ? tmp8144 : tmp8147;
  assign tmp8128 = s5 ? tmp8129 : tmp8143;
  assign tmp8113 = s6 ? tmp8114 : tmp8128;
  assign tmp8157 = s1 ? tmp8124 : tmp7950;
  assign tmp8156 = s2 ? tmp8120 : tmp8157;
  assign tmp8159 = s1 ? tmp7950 : tmp7125;
  assign tmp8158 = s2 ? tmp8159 : tmp7952;
  assign tmp8155 = s3 ? tmp8156 : tmp8158;
  assign tmp8154 = s4 ? tmp8115 : tmp8155;
  assign tmp8164 = s1 ? tmp7952 : tmp7955;
  assign tmp8163 = s2 ? tmp7990 : tmp8164;
  assign tmp8165 = s2 ? tmp7952 : tmp8120;
  assign tmp8162 = s3 ? tmp8163 : tmp8165;
  assign tmp8167 = s2 ? tmp8136 : tmp7952;
  assign tmp8169 = s1 ? tmp7952 : tmp7122;
  assign tmp8168 = s2 ? tmp8169 : tmp7451;
  assign tmp8166 = s3 ? tmp8167 : tmp8168;
  assign tmp8161 = s4 ? tmp8162 : tmp8166;
  assign tmp8172 = s2 ? tmp8120 : 1;
  assign tmp8171 = s3 ? tmp8172 : tmp8109;
  assign tmp8175 = s1 ? 1 : tmp7952;
  assign tmp8174 = s2 ? tmp8175 : tmp7952;
  assign tmp8176 = s1 ? 1 : tmp7122;
  assign tmp8173 = s3 ? tmp8174 : tmp8176;
  assign tmp8170 = s4 ? tmp8171 : tmp8173;
  assign tmp8160 = s5 ? tmp8161 : tmp8170;
  assign tmp8153 = s6 ? tmp8154 : tmp8160;
  assign tmp8112 = ~(s7 ? tmp8113 : tmp8153);
  assign tmp8046 = s8 ? tmp8047 : tmp8112;
  assign tmp8178 = s7 ? tmp8113 : tmp8153;
  assign tmp8183 = ~(s2 ? tmp7242 : tmp7125);
  assign tmp8182 = s3 ? tmp7230 : tmp8183;
  assign tmp8185 = s2 ? tmp7236 : tmp7392;
  assign tmp8186 = ~(s2 ? tmp7380 : tmp7231);
  assign tmp8184 = ~(s3 ? tmp8185 : tmp8186);
  assign tmp8181 = s4 ? tmp8182 : tmp8184;
  assign tmp8189 = s3 ? tmp7240 : tmp7248;
  assign tmp8192 = s1 ? tmp7329 : tmp7133;
  assign tmp8191 = s2 ? tmp7504 : tmp8192;
  assign tmp8193 = s2 ? tmp7316 : tmp7253;
  assign tmp8190 = s3 ? tmp8191 : tmp8193;
  assign tmp8188 = s4 ? tmp8189 : tmp8190;
  assign tmp8197 = s1 ? tmp7133 : tmp7222;
  assign tmp8196 = s2 ? tmp8197 : tmp7241;
  assign tmp8195 = s3 ? tmp8196 : tmp7261;
  assign tmp8200 = s1 ? tmp7222 : 1;
  assign tmp8199 = s2 ? tmp7236 : tmp8200;
  assign tmp8201 = s2 ? tmp7221 : tmp7135;
  assign tmp8198 = s3 ? tmp8199 : tmp8201;
  assign tmp8194 = s4 ? tmp8195 : tmp8198;
  assign tmp8187 = ~(s5 ? tmp8188 : tmp8194);
  assign tmp8180 = s6 ? tmp8181 : tmp8187;
  assign tmp8205 = ~(s2 ? tmp7409 : tmp7231);
  assign tmp8204 = ~(s3 ? tmp8185 : tmp8205);
  assign tmp8203 = s4 ? tmp8182 : tmp8204;
  assign tmp8208 = s3 ? tmp7597 : tmp7248;
  assign tmp8209 = s3 ? tmp7919 : tmp7450;
  assign tmp8207 = s4 ? tmp8208 : tmp8209;
  assign tmp8212 = s2 ? tmp7236 : 1;
  assign tmp8211 = s3 ? tmp8212 : tmp7261;
  assign tmp8210 = s4 ? tmp8211 : tmp7125;
  assign tmp8206 = ~(s5 ? tmp8207 : tmp8210);
  assign tmp8202 = s6 ? tmp8203 : tmp8206;
  assign tmp8179 = ~(s7 ? tmp8180 : tmp8202);
  assign tmp8177 = ~(s8 ? tmp8178 : tmp8179);
  assign tmp8045 = s9 ? tmp8046 : tmp8177;
  assign tmp8219 = ~(s2 ? tmp8054 : tmp7122);
  assign tmp8218 = s3 ? tmp8051 : tmp8219;
  assign tmp8222 = s1 ? tmp7132 : tmp7122;
  assign tmp8221 = s2 ? tmp8222 : tmp8061;
  assign tmp8220 = ~(s3 ? tmp8221 : tmp8062);
  assign tmp8217 = s4 ? tmp8218 : tmp8220;
  assign tmp8226 = s2 ? tmp8068 : tmp8054;
  assign tmp8225 = s3 ? tmp8226 : tmp8101;
  assign tmp8229 = s1 ? tmp7124 : tmp7329;
  assign tmp8230 = s1 ? tmp7329 : tmp7132;
  assign tmp8228 = s2 ? tmp8229 : tmp8230;
  assign tmp8227 = s3 ? tmp8228 : tmp8077;
  assign tmp8224 = s4 ? tmp8225 : tmp8227;
  assign tmp8223 = ~(s5 ? tmp8224 : tmp8080);
  assign tmp8216 = s6 ? tmp8217 : tmp8223;
  assign tmp8233 = ~(s3 ? tmp8221 : tmp8095);
  assign tmp8232 = s4 ? tmp8218 : tmp8233;
  assign tmp8237 = s2 ? tmp8068 : tmp7122;
  assign tmp8236 = s3 ? tmp8237 : tmp8101;
  assign tmp8239 = s2 ? tmp8229 : tmp7122;
  assign tmp8238 = s3 ? tmp8239 : tmp8105;
  assign tmp8235 = s4 ? tmp8236 : tmp8238;
  assign tmp8242 = s2 ? tmp7170 : 1;
  assign tmp8241 = s3 ? tmp8242 : tmp8109;
  assign tmp8243 = s3 ? tmp8111 : tmp8176;
  assign tmp8240 = s4 ? tmp8241 : tmp8243;
  assign tmp8234 = ~(s5 ? tmp8235 : tmp8240);
  assign tmp8231 = s6 ? tmp8232 : tmp8234;
  assign tmp8215 = s7 ? tmp8216 : tmp8231;
  assign tmp8214 = s8 ? tmp8215 : tmp8216;
  assign tmp8248 = s4 ? tmp8107 : tmp8243;
  assign tmp8247 = ~(s5 ? tmp8097 : tmp8248);
  assign tmp8246 = s6 ? tmp8093 : tmp8247;
  assign tmp8245 = s7 ? tmp8246 : tmp8202;
  assign tmp8250 = ~(s6 ? tmp8232 : tmp8234);
  assign tmp8249 = ~(s7 ? tmp8153 : tmp8250);
  assign tmp8244 = s8 ? tmp8245 : tmp8249;
  assign tmp8213 = s9 ? tmp8214 : tmp8244;
  assign tmp8044 = s10 ? tmp8045 : tmp8213;
  assign tmp8254 = s7 ? tmp8092 : tmp8202;
  assign tmp8253 = s8 ? tmp8254 : tmp8249;
  assign tmp8252 = s9 ? tmp8214 : tmp8253;
  assign tmp8251 = s10 ? tmp8045 : tmp8252;
  assign tmp8043 = ~(s11 ? tmp8044 : tmp8251);
  assign tmp7909 = s12 ? tmp7910 : tmp8043;
  assign tmp8261 = s2 ? tmp7230 : tmp7409;
  assign tmp8260 = s3 ? tmp7380 : tmp8261;
  assign tmp8263 = s2 ? tmp7409 : 1;
  assign tmp8262 = s3 ? tmp8263 : tmp7848;
  assign tmp8259 = s4 ? tmp8260 : tmp8262;
  assign tmp8266 = s3 ? tmp7852 : tmp8186;
  assign tmp8268 = s2 ? tmp7590 : 1;
  assign tmp8269 = s2 ? tmp7380 : tmp7300;
  assign tmp8267 = ~(s3 ? tmp8268 : tmp8269);
  assign tmp8265 = s4 ? tmp8266 : tmp8267;
  assign tmp8272 = ~(s2 ? tmp7350 : tmp7830);
  assign tmp8271 = s3 ? tmp7432 : tmp8272;
  assign tmp8274 = s2 ? tmp7350 : tmp7590;
  assign tmp8275 = s2 ? tmp7350 : tmp7409;
  assign tmp8273 = ~(s3 ? tmp8274 : tmp8275);
  assign tmp8270 = s4 ? tmp8271 : tmp8273;
  assign tmp8264 = ~(s5 ? tmp8265 : tmp8270);
  assign tmp8258 = s6 ? tmp8259 : tmp8264;
  assign tmp8278 = s3 ? tmp8263 : tmp7868;
  assign tmp8277 = s4 ? tmp8260 : tmp8278;
  assign tmp8281 = s3 ? tmp7872 : tmp8205;
  assign tmp8282 = ~(s3 ? tmp8268 : tmp7409);
  assign tmp8280 = s4 ? tmp8281 : tmp8282;
  assign tmp8284 = s3 ? tmp7432 : tmp7875;
  assign tmp8283 = s4 ? tmp8284 : tmp7125;
  assign tmp8279 = ~(s5 ? tmp8280 : tmp8283);
  assign tmp8276 = s6 ? tmp8277 : tmp8279;
  assign tmp8257 = s7 ? tmp8258 : tmp8276;
  assign tmp8286 = s8 ? tmp8257 : tmp8258;
  assign tmp8285 = s9 ? tmp8286 : tmp8276;
  assign tmp8256 = s10 ? tmp8257 : tmp8285;
  assign tmp8295 = s1 ? tmp7952 : tmp7980;
  assign tmp8296 = s2 ? tmp7980 : tmp8175;
  assign tmp8294 = s3 ? tmp8295 : tmp8296;
  assign tmp8299 = s1 ? tmp7952 : 1;
  assign tmp8298 = s2 ? tmp8120 : tmp8299;
  assign tmp8301 = s1 ? tmp7952 : tmp8137;
  assign tmp8300 = s2 ? tmp7451 : tmp8301;
  assign tmp8297 = s3 ? tmp8298 : tmp8300;
  assign tmp8293 = s4 ? tmp8294 : tmp8297;
  assign tmp8306 = s1 ? 1 : tmp7980;
  assign tmp8307 = s1 ? tmp7133 : tmp7952;
  assign tmp8305 = s2 ? tmp8306 : tmp8307;
  assign tmp8304 = s3 ? tmp8131 : tmp8305;
  assign tmp8310 = s1 ? tmp8137 : 1;
  assign tmp8311 = s1 ? 1 : tmp7955;
  assign tmp8309 = s2 ? tmp8310 : tmp8311;
  assign tmp8312 = s2 ? tmp8295 : tmp7253;
  assign tmp8308 = s3 ? tmp8309 : tmp8312;
  assign tmp8303 = s4 ? tmp8304 : tmp8308;
  assign tmp8315 = s2 ? tmp7990 : 1;
  assign tmp8317 = s1 ? tmp7222 : tmp8137;
  assign tmp8316 = s2 ? tmp7235 : tmp8317;
  assign tmp8314 = s3 ? tmp8315 : tmp8316;
  assign tmp8320 = s1 ? tmp7983 : tmp7125;
  assign tmp8319 = s2 ? tmp8320 : tmp8150;
  assign tmp8322 = s1 ? tmp7222 : tmp7980;
  assign tmp8323 = s1 ? tmp8137 : tmp7125;
  assign tmp8321 = s2 ? tmp8322 : tmp8323;
  assign tmp8318 = s3 ? tmp8319 : tmp8321;
  assign tmp8313 = s4 ? tmp8314 : tmp8318;
  assign tmp8302 = s5 ? tmp8303 : tmp8313;
  assign tmp8292 = s6 ? tmp8293 : tmp8302;
  assign tmp8328 = s2 ? tmp8175 : tmp8307;
  assign tmp8327 = s3 ? tmp8163 : tmp8328;
  assign tmp8330 = s2 ? tmp8310 : tmp7952;
  assign tmp8331 = s2 ? tmp7952 : tmp7451;
  assign tmp8329 = s3 ? tmp8330 : tmp8331;
  assign tmp8326 = s4 ? tmp8327 : tmp8329;
  assign tmp8335 = s1 ? tmp7125 : tmp7952;
  assign tmp8334 = s2 ? tmp7135 : tmp8335;
  assign tmp8333 = s3 ? tmp8315 : tmp8334;
  assign tmp8337 = s2 ? tmp7125 : tmp7952;
  assign tmp8338 = s2 ? tmp8335 : tmp7125;
  assign tmp8336 = s3 ? tmp8337 : tmp8338;
  assign tmp8332 = s4 ? tmp8333 : tmp8336;
  assign tmp8325 = s5 ? tmp8326 : tmp8332;
  assign tmp8324 = s6 ? tmp8293 : tmp8325;
  assign tmp8291 = s7 ? tmp8292 : tmp8324;
  assign tmp8346 = l1 ? 1 : tmp7146;
  assign tmp8345 = s0 ? tmp8346 : tmp7952;
  assign tmp8344 = s1 ? tmp7952 : tmp8345;
  assign tmp8343 = s2 ? tmp7451 : tmp8344;
  assign tmp8342 = s3 ? tmp8298 : tmp8343;
  assign tmp8341 = s4 ? tmp8294 : tmp8342;
  assign tmp8352 = s0 ? tmp8346 : 1;
  assign tmp8351 = s1 ? tmp8352 : tmp7952;
  assign tmp8350 = s2 ? tmp8306 : tmp8351;
  assign tmp8349 = s3 ? tmp8131 : tmp8350;
  assign tmp8348 = s4 ? tmp8349 : tmp8308;
  assign tmp8357 = s0 ? tmp7125 : tmp8346;
  assign tmp8356 = s1 ? tmp7983 : tmp8357;
  assign tmp8355 = s2 ? tmp8356 : tmp8150;
  assign tmp8354 = s3 ? tmp8355 : tmp8321;
  assign tmp8353 = s4 ? tmp8314 : tmp8354;
  assign tmp8347 = s5 ? tmp8348 : tmp8353;
  assign tmp8340 = s6 ? tmp8341 : tmp8347;
  assign tmp8362 = s2 ? tmp8175 : tmp8351;
  assign tmp8361 = s3 ? tmp8163 : tmp8362;
  assign tmp8360 = s4 ? tmp8361 : tmp8329;
  assign tmp8366 = s1 ? tmp7125 : tmp8357;
  assign tmp8365 = s2 ? tmp8366 : tmp7952;
  assign tmp8364 = s3 ? tmp8365 : tmp8338;
  assign tmp8363 = s4 ? tmp8333 : tmp8364;
  assign tmp8359 = s5 ? tmp8360 : tmp8363;
  assign tmp8358 = s6 ? tmp8341 : tmp8359;
  assign tmp8339 = s7 ? tmp8340 : tmp8358;
  assign tmp8290 = s8 ? tmp8291 : tmp8339;
  assign tmp8371 = s3 ? tmp7221 : tmp7782;
  assign tmp8373 = s2 ? tmp7236 : tmp7135;
  assign tmp8372 = s3 ? tmp8373 : tmp7800;
  assign tmp8370 = s4 ? tmp8371 : tmp8372;
  assign tmp8377 = s2 ? tmp7241 : tmp7235;
  assign tmp8378 = s2 ? tmp7786 : tmp7236;
  assign tmp8376 = s3 ? tmp8377 : tmp8378;
  assign tmp8380 = s2 ? tmp7135 : tmp7253;
  assign tmp8379 = s3 ? tmp8380 : tmp7252;
  assign tmp8375 = s4 ? tmp8376 : tmp8379;
  assign tmp8383 = s2 ? tmp7235 : tmp7242;
  assign tmp8382 = s3 ? tmp7654 : tmp8383;
  assign tmp8385 = s2 ? tmp7125 : tmp8200;
  assign tmp8386 = s2 ? tmp7222 : tmp7125;
  assign tmp8384 = s3 ? tmp8385 : tmp8386;
  assign tmp8381 = s4 ? tmp8382 : tmp8384;
  assign tmp8374 = s5 ? tmp8375 : tmp8381;
  assign tmp8369 = s6 ? tmp8370 : tmp8374;
  assign tmp8391 = s2 ? tmp7241 : tmp7388;
  assign tmp8392 = s2 ? tmp7451 : tmp7236;
  assign tmp8390 = s3 ? tmp8391 : tmp8392;
  assign tmp8394 = s2 ? tmp7135 : tmp7125;
  assign tmp8393 = s3 ? tmp8394 : tmp7450;
  assign tmp8389 = s4 ? tmp8390 : tmp8393;
  assign tmp8396 = s3 ? tmp7654 : tmp8394;
  assign tmp8395 = s4 ? tmp8396 : tmp7125;
  assign tmp8388 = s5 ? tmp8389 : tmp8395;
  assign tmp8387 = s6 ? tmp8370 : tmp8388;
  assign tmp8368 = s7 ? tmp8369 : tmp8387;
  assign tmp8367 = s8 ? tmp8339 : tmp8368;
  assign tmp8289 = s9 ? tmp8290 : tmp8367;
  assign tmp8404 = s2 ? tmp7952 : tmp7253;
  assign tmp8403 = s3 ? tmp8309 : tmp8404;
  assign tmp8402 = s4 ? tmp8304 : tmp8403;
  assign tmp8401 = s5 ? tmp8402 : tmp8313;
  assign tmp8400 = s6 ? tmp8293 : tmp8401;
  assign tmp8399 = s7 ? tmp8400 : tmp8324;
  assign tmp8398 = s8 ? tmp8399 : tmp8400;
  assign tmp8410 = s3 ? tmp8337 : tmp8335;
  assign tmp8409 = s4 ? tmp8333 : tmp8410;
  assign tmp8408 = s5 ? tmp8326 : tmp8409;
  assign tmp8407 = s6 ? tmp8293 : tmp8408;
  assign tmp8406 = s7 ? tmp8407 : tmp8387;
  assign tmp8415 = s3 ? tmp8365 : tmp8335;
  assign tmp8414 = s4 ? tmp8333 : tmp8415;
  assign tmp8413 = s5 ? tmp8360 : tmp8414;
  assign tmp8412 = s6 ? tmp8341 : tmp8413;
  assign tmp8411 = s7 ? tmp8412 : tmp8407;
  assign tmp8405 = s8 ? tmp8406 : tmp8411;
  assign tmp8397 = s9 ? tmp8398 : tmp8405;
  assign tmp8288 = s10 ? tmp8289 : tmp8397;
  assign tmp8419 = s7 ? tmp8324 : tmp8387;
  assign tmp8420 = s7 ? tmp8358 : tmp8324;
  assign tmp8418 = s8 ? tmp8419 : tmp8420;
  assign tmp8417 = s9 ? tmp8398 : tmp8418;
  assign tmp8416 = s10 ? tmp8289 : tmp8417;
  assign tmp8287 = ~(s11 ? tmp8288 : tmp8416);
  assign tmp8255 = ~(s12 ? tmp8256 : tmp8287);
  assign tmp7908 = s13 ? tmp7909 : tmp8255;
  assign tmp7773 = s14 ? tmp7774 : tmp7908;
  assign tmp7110 = s15 ? tmp7111 : tmp7773;
  assign tmp8432 = s3 ? tmp7178 : tmp7201;
  assign tmp8431 = s4 ? tmp7207 : tmp8432;
  assign tmp8430 = s5 ? tmp8431 : tmp7180;
  assign tmp8429 = s6 ? tmp7203 : tmp8430;
  assign tmp8428 = s7 ? tmp7186 : tmp8429;
  assign tmp8427 = s8 ? tmp7117 : tmp8428;
  assign tmp8438 = s3 ? tmp7125 : tmp7252;
  assign tmp8439 = s3 ? tmp7234 : tmp7654;
  assign tmp8437 = s4 ? tmp8438 : tmp8439;
  assign tmp8436 = s5 ? tmp8437 : tmp7238;
  assign tmp8435 = s6 ? tmp7217 : tmp8436;
  assign tmp8443 = s3 ? tmp7255 : tmp7654;
  assign tmp8442 = s4 ? tmp8438 : tmp8443;
  assign tmp8441 = s5 ? tmp8442 : tmp7257;
  assign tmp8440 = s6 ? tmp7246 : tmp8441;
  assign tmp8434 = s7 ? tmp8435 : tmp8440;
  assign tmp8433 = s8 ? tmp8428 : tmp8434;
  assign tmp8426 = s9 ? tmp8427 : tmp8433;
  assign tmp8445 = s8 ? tmp8428 : tmp7186;
  assign tmp8447 = s7 ? tmp7271 : tmp8440;
  assign tmp8451 = s3 ? tmp7275 : tmp7201;
  assign tmp8450 = s4 ? tmp7207 : tmp8451;
  assign tmp8449 = s5 ? tmp8450 : tmp7180;
  assign tmp8448 = s6 ? tmp7203 : tmp8449;
  assign tmp8446 = s8 ? tmp8447 : tmp8448;
  assign tmp8444 = s9 ? tmp8445 : tmp8446;
  assign tmp8425 = s10 ? tmp8426 : tmp8444;
  assign tmp8455 = s7 ? tmp7166 : tmp8440;
  assign tmp8454 = s8 ? tmp8455 : tmp8429;
  assign tmp8453 = s9 ? tmp8445 : tmp8454;
  assign tmp8452 = s10 ? tmp8426 : tmp8453;
  assign tmp8424 = s11 ? tmp8425 : tmp8452;
  assign tmp8466 = s1 ? tmp7228 : tmp7222;
  assign tmp8465 = s2 ? tmp7388 : tmp8466;
  assign tmp8464 = s3 ? tmp7125 : tmp8465;
  assign tmp8463 = s4 ? tmp7125 : tmp8464;
  assign tmp8470 = ~(s2 ? tmp7395 : 0);
  assign tmp8469 = s3 ? tmp7297 : tmp8470;
  assign tmp8468 = s4 ? tmp8469 : 1;
  assign tmp8467 = s5 ? tmp8468 : 1;
  assign tmp8462 = s6 ? tmp8463 : tmp8467;
  assign tmp8475 = ~(s2 ? tmp7407 : 0);
  assign tmp8474 = s3 ? tmp7406 : tmp8475;
  assign tmp8473 = s4 ? tmp8474 : 1;
  assign tmp8472 = s5 ? tmp8473 : 1;
  assign tmp8471 = s6 ? tmp8463 : tmp8472;
  assign tmp8461 = s7 ? tmp8462 : tmp8471;
  assign tmp8480 = s2 ? tmp7388 : tmp7221;
  assign tmp8479 = s3 ? tmp7125 : tmp8480;
  assign tmp8478 = s4 ? tmp7125 : tmp8479;
  assign tmp8483 = s3 ? tmp7248 : tmp7794;
  assign tmp8482 = s4 ? tmp8483 : 1;
  assign tmp8481 = s5 ? tmp8482 : 1;
  assign tmp8477 = s6 ? tmp8478 : tmp8481;
  assign tmp8487 = s3 ? tmp7450 : tmp7256;
  assign tmp8486 = s4 ? tmp8487 : 1;
  assign tmp8485 = s5 ? tmp8486 : 1;
  assign tmp8484 = s6 ? tmp8478 : tmp8485;
  assign tmp8476 = s7 ? tmp8477 : tmp8484;
  assign tmp8460 = s8 ? tmp8461 : tmp8476;
  assign tmp8459 = s9 ? tmp8460 : tmp8476;
  assign tmp8489 = s8 ? tmp8476 : tmp8477;
  assign tmp8495 = s2 ? tmp7135 : tmp8466;
  assign tmp8494 = s3 ? tmp7125 : tmp8495;
  assign tmp8493 = s4 ? tmp7125 : tmp8494;
  assign tmp8492 = s6 ? tmp8493 : tmp8472;
  assign tmp8498 = s3 ? tmp7125 : tmp7220;
  assign tmp8497 = s4 ? tmp7125 : tmp8498;
  assign tmp8496 = s6 ? tmp8497 : tmp8485;
  assign tmp8491 = s7 ? tmp8492 : tmp8496;
  assign tmp8490 = s8 ? tmp8491 : tmp8496;
  assign tmp8488 = s9 ? tmp8489 : tmp8490;
  assign tmp8458 = s10 ? tmp8459 : tmp8488;
  assign tmp8502 = s7 ? tmp8471 : tmp8484;
  assign tmp8501 = s8 ? tmp8502 : tmp8484;
  assign tmp8500 = s9 ? tmp8489 : tmp8501;
  assign tmp8499 = s10 ? tmp8459 : tmp8500;
  assign tmp8457 = s11 ? tmp8458 : tmp8499;
  assign tmp8456 = s12 ? tmp7283 : tmp8457;
  assign tmp8423 = s13 ? tmp8424 : tmp8456;
  assign tmp8515 = ~(s1 ? tmp7230 : tmp7231);
  assign tmp8514 = s2 ? tmp7292 : tmp8515;
  assign tmp8516 = s2 ? tmp7227 : tmp7578;
  assign tmp8513 = s3 ? tmp8514 : tmp8516;
  assign tmp8518 = s2 ? tmp7304 : 1;
  assign tmp8517 = ~(s3 ? tmp7349 : tmp8518);
  assign tmp8512 = s4 ? tmp8513 : tmp8517;
  assign tmp8511 = s5 ? tmp8512 : 0;
  assign tmp8510 = s6 ? tmp7313 : tmp8511;
  assign tmp8523 = s2 ? tmp7632 : tmp7125;
  assign tmp8522 = s3 ? tmp8523 : tmp8516;
  assign tmp8524 = ~(s3 ? tmp7349 : tmp8268);
  assign tmp8521 = s4 ? tmp8522 : tmp8524;
  assign tmp8520 = s5 ? tmp8521 : 0;
  assign tmp8519 = s6 ? tmp7332 : tmp8520;
  assign tmp8509 = ~(s7 ? tmp8510 : tmp8519);
  assign tmp8508 = s8 ? 1 : tmp8509;
  assign tmp8507 = s9 ? tmp8508 : tmp8509;
  assign tmp8527 = s7 ? tmp8510 : tmp8519;
  assign tmp8526 = s8 ? tmp8527 : tmp8510;
  assign tmp8534 = s2 ? tmp7298 : tmp7578;
  assign tmp8533 = s3 ? tmp8523 : tmp8534;
  assign tmp8532 = s4 ? tmp8533 : tmp8524;
  assign tmp8531 = s5 ? tmp8532 : 0;
  assign tmp8530 = ~(s6 ? tmp7332 : tmp8531);
  assign tmp8529 = s7 ? 1 : tmp8530;
  assign tmp8528 = ~(s8 ? tmp8529 : tmp8530);
  assign tmp8525 = ~(s9 ? tmp8526 : tmp8528);
  assign tmp8506 = s10 ? tmp8507 : tmp8525;
  assign tmp8539 = ~(s6 ? tmp7332 : tmp8520);
  assign tmp8538 = s7 ? 1 : tmp8539;
  assign tmp8537 = ~(s8 ? tmp8538 : tmp8539);
  assign tmp8536 = ~(s9 ? tmp8526 : tmp8537);
  assign tmp8535 = s10 ? tmp8507 : tmp8536;
  assign tmp8505 = s11 ? tmp8506 : tmp8535;
  assign tmp8547 = s4 ? tmp7561 : tmp7540;
  assign tmp8546 = s5 ? tmp8547 : tmp7543;
  assign tmp8545 = s6 ? tmp7531 : tmp8546;
  assign tmp8544 = s7 ? tmp7550 : tmp8545;
  assign tmp8552 = s2 ? tmp8222 : tmp7131;
  assign tmp8553 = s2 ? tmp7504 : tmp8078;
  assign tmp8551 = s3 ? tmp8552 : tmp8553;
  assign tmp8550 = s4 ? tmp7120 : tmp8551;
  assign tmp8558 = s1 ? tmp7132 : tmp7138;
  assign tmp8559 = s1 ? tmp7138 : tmp7128;
  assign tmp8557 = s2 ? tmp8558 : tmp8559;
  assign tmp8561 = ~(s1 ? 1 : tmp8052);
  assign tmp8560 = s2 ? tmp7197 : tmp8561;
  assign tmp8556 = s3 ? tmp8557 : tmp8560;
  assign tmp8564 = s1 ? tmp8051 : tmp7231;
  assign tmp8565 = ~(s1 ? tmp7125 : tmp7132);
  assign tmp8563 = s2 ? tmp8564 : tmp8565;
  assign tmp8568 = s0 ? tmp7146 : tmp8052;
  assign tmp8567 = s1 ? tmp8568 : tmp7497;
  assign tmp8566 = s2 ? tmp8567 : 1;
  assign tmp8562 = ~(s3 ? tmp8563 : tmp8566);
  assign tmp8555 = s4 ? tmp8556 : tmp8562;
  assign tmp8572 = s1 ? tmp7148 : tmp7146;
  assign tmp8571 = s2 ? tmp7520 : tmp8572;
  assign tmp8570 = s3 ? tmp8571 : tmp7522;
  assign tmp8573 = s3 ? tmp8571 : tmp7527;
  assign tmp8569 = ~(s4 ? tmp8570 : tmp8573);
  assign tmp8554 = s5 ? tmp8555 : tmp8569;
  assign tmp8549 = s6 ? tmp8550 : tmp8554;
  assign tmp8577 = s2 ? tmp8222 : tmp7170;
  assign tmp8578 = s2 ? tmp7298 : tmp8078;
  assign tmp8576 = s3 ? tmp8577 : tmp8578;
  assign tmp8575 = s4 ? tmp7120 : tmp8576;
  assign tmp8582 = s2 ? tmp8222 : tmp7209;
  assign tmp8583 = s2 ? tmp7211 : tmp8561;
  assign tmp8581 = s3 ? tmp8582 : tmp8583;
  assign tmp8586 = ~(s1 ? tmp7125 : tmp7122);
  assign tmp8585 = s2 ? tmp8564 : tmp8586;
  assign tmp8584 = ~(s3 ? tmp8585 : tmp8566);
  assign tmp8580 = s4 ? tmp8581 : tmp8584;
  assign tmp8589 = s2 ? tmp7520 : tmp7155;
  assign tmp8588 = s3 ? tmp8589 : tmp7546;
  assign tmp8587 = ~(s4 ? tmp8588 : tmp7547);
  assign tmp8579 = s5 ? tmp8580 : tmp8587;
  assign tmp8574 = s6 ? tmp8575 : tmp8579;
  assign tmp8548 = ~(s7 ? tmp8549 : tmp8574);
  assign tmp8543 = s8 ? tmp8544 : tmp8548;
  assign tmp8591 = s7 ? tmp8549 : tmp8574;
  assign tmp8594 = s4 ? tmp7125 : tmp7572;
  assign tmp8598 = s2 ? tmp8197 : tmp7242;
  assign tmp8597 = s3 ? tmp8598 : tmp7577;
  assign tmp8596 = s4 ? tmp8597 : tmp7579;
  assign tmp8601 = s2 ? tmp7392 : tmp8515;
  assign tmp8600 = s3 ? tmp8601 : tmp7584;
  assign tmp8602 = s3 ? tmp8601 : tmp7589;
  assign tmp8599 = s4 ? tmp8600 : tmp8602;
  assign tmp8595 = s5 ? tmp8596 : tmp8599;
  assign tmp8593 = s6 ? tmp8594 : tmp8595;
  assign tmp8604 = s4 ? tmp7125 : tmp7593;
  assign tmp8608 = s2 ? tmp7236 : tmp7125;
  assign tmp8607 = s3 ? tmp8608 : tmp7577;
  assign tmp8606 = s4 ? tmp8607 : tmp7579;
  assign tmp8610 = s3 ? tmp7416 : tmp7601;
  assign tmp8609 = s4 ? tmp8610 : tmp7602;
  assign tmp8605 = s5 ? tmp8606 : tmp8609;
  assign tmp8603 = s6 ? tmp8604 : tmp8605;
  assign tmp8592 = s7 ? tmp8593 : tmp8603;
  assign tmp8590 = ~(s8 ? tmp8591 : tmp8592);
  assign tmp8542 = s9 ? tmp8543 : tmp8590;
  assign tmp8612 = s8 ? tmp8591 : tmp8549;
  assign tmp8617 = s4 ? tmp7561 : tmp7615;
  assign tmp8616 = s5 ? tmp8617 : tmp7543;
  assign tmp8615 = s6 ? tmp7531 : tmp8616;
  assign tmp8618 = ~(s6 ? tmp8604 : tmp8605);
  assign tmp8614 = s7 ? tmp8615 : tmp8618;
  assign tmp8624 = s1 ? tmp8568 : tmp7146;
  assign tmp8623 = s2 ? tmp8624 : 1;
  assign tmp8622 = ~(s3 ? tmp8585 : tmp8623);
  assign tmp8621 = s4 ? tmp8581 : tmp8622;
  assign tmp8620 = s5 ? tmp8621 : tmp8587;
  assign tmp8619 = ~(s6 ? tmp8575 : tmp8620);
  assign tmp8613 = ~(s8 ? tmp8614 : tmp8619);
  assign tmp8611 = ~(s9 ? tmp8612 : tmp8613);
  assign tmp8541 = s10 ? tmp8542 : tmp8611;
  assign tmp8628 = s7 ? tmp8545 : tmp8618;
  assign tmp8629 = ~(s6 ? tmp8575 : tmp8579);
  assign tmp8627 = ~(s8 ? tmp8628 : tmp8629);
  assign tmp8626 = ~(s9 ? tmp8612 : tmp8627);
  assign tmp8625 = s10 ? tmp8542 : tmp8626;
  assign tmp8540 = s11 ? tmp8541 : tmp8625;
  assign tmp8504 = s12 ? tmp8505 : tmp8540;
  assign tmp8637 = s2 ? tmp7122 : tmp8055;
  assign tmp8636 = s3 ? tmp7121 : tmp8637;
  assign tmp8640 = s1 ? tmp8056 : tmp7228;
  assign tmp8639 = s2 ? tmp7127 : tmp8640;
  assign tmp8641 = s2 ? tmp7636 : tmp7190;
  assign tmp8638 = s3 ? tmp8639 : tmp8641;
  assign tmp8635 = s4 ? tmp8636 : tmp8638;
  assign tmp8646 = s1 ? tmp8056 : tmp8079;
  assign tmp8648 = ~(s0 ? tmp7122 : 0);
  assign tmp8647 = ~(s1 ? tmp8051 : tmp8648);
  assign tmp8645 = s2 ? tmp8646 : tmp8647;
  assign tmp8650 = ~(s1 ? 1 : tmp7122);
  assign tmp8649 = ~(s2 ? tmp8051 : tmp8650);
  assign tmp8644 = s3 ? tmp8645 : tmp8649;
  assign tmp8653 = s1 ? tmp7138 : tmp7125;
  assign tmp8652 = s2 ? tmp8653 : tmp7179;
  assign tmp8655 = s1 ? tmp7122 : 1;
  assign tmp8654 = s2 ? tmp8655 : 1;
  assign tmp8651 = s3 ? tmp8652 : tmp8654;
  assign tmp8643 = s4 ? tmp8644 : tmp8651;
  assign tmp8658 = s2 ? tmp8655 : tmp8054;
  assign tmp8657 = s3 ? tmp8658 : 1;
  assign tmp8660 = s2 ? 1 : tmp7122;
  assign tmp8659 = s3 ? tmp8660 : 1;
  assign tmp8656 = s4 ? tmp8657 : tmp8659;
  assign tmp8642 = s5 ? tmp8643 : tmp8656;
  assign tmp8634 = s6 ? tmp8635 : tmp8642;
  assign tmp8665 = s1 ? tmp8056 : tmp7125;
  assign tmp8664 = s2 ? tmp7127 : tmp8665;
  assign tmp8663 = s3 ? tmp8664 : tmp7189;
  assign tmp8662 = s4 ? tmp8636 : tmp8663;
  assign tmp8669 = s2 ? tmp8055 : tmp8100;
  assign tmp8670 = s2 ? tmp7122 : tmp8176;
  assign tmp8668 = s3 ? tmp8669 : tmp8670;
  assign tmp8672 = s2 ? tmp8653 : tmp7122;
  assign tmp8671 = s3 ? tmp8672 : tmp8654;
  assign tmp8667 = s4 ? tmp8668 : tmp8671;
  assign tmp8674 = s3 ? tmp8655 : 1;
  assign tmp8673 = s4 ? tmp8674 : tmp8659;
  assign tmp8666 = s5 ? tmp8667 : tmp8673;
  assign tmp8661 = s6 ? tmp8662 : tmp8666;
  assign tmp8633 = s7 ? tmp8634 : tmp8661;
  assign tmp8680 = s2 ? tmp7636 : tmp7125;
  assign tmp8679 = s3 ? tmp7634 : tmp8680;
  assign tmp8678 = s4 ? tmp7630 : tmp8679;
  assign tmp8684 = ~(s2 ? tmp7230 : tmp7326);
  assign tmp8683 = s3 ? tmp7640 : tmp8684;
  assign tmp8685 = s3 ? tmp7644 : tmp7794;
  assign tmp8682 = s4 ? tmp8683 : tmp8685;
  assign tmp8687 = s3 ? tmp7125 : 1;
  assign tmp8688 = s3 ? tmp7800 : tmp7256;
  assign tmp8686 = s4 ? tmp8687 : tmp8688;
  assign tmp8681 = s5 ? tmp8682 : tmp8686;
  assign tmp8677 = s6 ? tmp8678 : tmp8681;
  assign tmp8691 = s3 ? tmp7631 : tmp8394;
  assign tmp8690 = s4 ? tmp7630 : tmp8691;
  assign tmp8694 = s3 ? tmp7651 : tmp7248;
  assign tmp8693 = s4 ? tmp8694 : tmp7643;
  assign tmp8692 = s5 ? tmp8693 : tmp8687;
  assign tmp8689 = s6 ? tmp8690 : tmp8692;
  assign tmp8676 = s7 ? tmp8677 : tmp8689;
  assign tmp8675 = s8 ? tmp8633 : tmp8676;
  assign tmp8632 = s9 ? tmp8633 : tmp8675;
  assign tmp8701 = s2 ? tmp7636 : tmp7121;
  assign tmp8700 = s3 ? tmp8639 : tmp8701;
  assign tmp8699 = s4 ? tmp8636 : tmp8700;
  assign tmp8704 = s3 ? tmp8645 : tmp8070;
  assign tmp8707 = s1 ? tmp7122 : tmp7133;
  assign tmp8706 = s2 ? tmp8707 : 1;
  assign tmp8705 = s3 ? tmp8652 : tmp8706;
  assign tmp8703 = s4 ? tmp8704 : tmp8705;
  assign tmp8711 = s1 ? tmp7122 : tmp7125;
  assign tmp8712 = s1 ? tmp7124 : tmp7122;
  assign tmp8710 = s2 ? tmp8711 : tmp8712;
  assign tmp8709 = s3 ? tmp8710 : 1;
  assign tmp8714 = s2 ? tmp7451 : tmp7122;
  assign tmp8713 = s3 ? tmp8714 : tmp7256;
  assign tmp8708 = s4 ? tmp8709 : tmp8713;
  assign tmp8702 = s5 ? tmp8703 : tmp8708;
  assign tmp8698 = s6 ? tmp8699 : tmp8702;
  assign tmp8718 = s2 ? tmp7135 : tmp7121;
  assign tmp8717 = s3 ? tmp8664 : tmp8718;
  assign tmp8716 = s4 ? tmp8636 : tmp8717;
  assign tmp8721 = s3 ? tmp8669 : tmp8101;
  assign tmp8720 = s4 ? tmp8721 : tmp8671;
  assign tmp8724 = s2 ? tmp8711 : tmp8655;
  assign tmp8723 = s3 ? tmp8724 : 1;
  assign tmp8725 = s3 ? tmp8111 : 1;
  assign tmp8722 = s4 ? tmp8723 : tmp8725;
  assign tmp8719 = s5 ? tmp8720 : tmp8722;
  assign tmp8715 = s6 ? tmp8716 : tmp8719;
  assign tmp8697 = s7 ? tmp8698 : tmp8715;
  assign tmp8696 = s8 ? tmp8697 : tmp8698;
  assign tmp8727 = s7 ? tmp8661 : tmp8689;
  assign tmp8726 = s8 ? tmp8727 : tmp8715;
  assign tmp8695 = s9 ? tmp8696 : tmp8726;
  assign tmp8631 = s10 ? tmp8632 : tmp8695;
  assign tmp8630 = ~(s12 ? tmp8631 : 1);
  assign tmp8503 = ~(s13 ? tmp8504 : tmp8630);
  assign tmp8422 = s14 ? tmp8423 : tmp8503;
  assign tmp8742 = ~(l4 ? 1 : 0);
  assign tmp8741 = ~(l2 ? 1 : tmp8742);
  assign tmp8740 = l1 ? 1 : tmp8741;
  assign tmp8743 = s0 ? tmp7125 : tmp8740;
  assign tmp8739 = s1 ? tmp8740 : tmp8743;
  assign tmp8745 = s1 ? tmp7132 : tmp8740;
  assign tmp8744 = s2 ? tmp8740 : tmp8745;
  assign tmp8738 = s3 ? tmp8739 : tmp8744;
  assign tmp8749 = s0 ? tmp8740 : 1;
  assign tmp8748 = s1 ? tmp8749 : tmp8740;
  assign tmp8750 = s1 ? tmp8749 : tmp7133;
  assign tmp8747 = s2 ? tmp8748 : tmp8750;
  assign tmp8751 = s2 ? tmp7504 : tmp8739;
  assign tmp8746 = s3 ? tmp8747 : tmp8751;
  assign tmp8737 = s4 ? tmp8738 : tmp8746;
  assign tmp8756 = s1 ? tmp8749 : 1;
  assign tmp8758 = s0 ? 1 : tmp8740;
  assign tmp8757 = s1 ? tmp8758 : tmp8740;
  assign tmp8755 = s2 ? tmp8756 : tmp8757;
  assign tmp8760 = s1 ? tmp7228 : tmp8740;
  assign tmp8759 = s2 ? tmp8740 : tmp8760;
  assign tmp8754 = s3 ? tmp8755 : tmp8759;
  assign tmp8765 = ~(l1 ? 1 : tmp8741);
  assign tmp8764 = s0 ? 1 : tmp8765;
  assign tmp8763 = s1 ? tmp8764 : tmp7231;
  assign tmp8766 = ~(s1 ? tmp7125 : tmp8749);
  assign tmp8762 = s2 ? tmp8763 : tmp8766;
  assign tmp8767 = ~(s2 ? tmp8739 : 0);
  assign tmp8761 = ~(s3 ? tmp8762 : tmp8767);
  assign tmp8753 = s4 ? tmp8754 : tmp8761;
  assign tmp8772 = s0 ? tmp8740 : 0;
  assign tmp8771 = s1 ? tmp8772 : tmp7293;
  assign tmp8770 = s2 ? tmp8771 : tmp7241;
  assign tmp8774 = ~(s1 ? 1 : tmp8764);
  assign tmp8773 = s2 ? tmp7437 : tmp8774;
  assign tmp8769 = s3 ? tmp8770 : tmp8773;
  assign tmp8778 = s0 ? tmp8740 : tmp7125;
  assign tmp8777 = s1 ? tmp8778 : tmp7125;
  assign tmp8779 = ~(s1 ? tmp8764 : 0);
  assign tmp8776 = s2 ? tmp8777 : tmp8779;
  assign tmp8782 = ~(s0 ? 1 : tmp8765);
  assign tmp8781 = s1 ? tmp7125 : tmp8782;
  assign tmp8783 = ~(s1 ? tmp8764 : tmp7230);
  assign tmp8780 = s2 ? tmp8781 : tmp8783;
  assign tmp8775 = s3 ? tmp8776 : tmp8780;
  assign tmp8768 = s4 ? tmp8769 : tmp8775;
  assign tmp8752 = s5 ? tmp8753 : tmp8768;
  assign tmp8736 = s6 ? tmp8737 : tmp8752;
  assign tmp8788 = s1 ? tmp8749 : tmp7125;
  assign tmp8787 = s2 ? tmp8748 : tmp8788;
  assign tmp8789 = s2 ? tmp7298 : tmp8739;
  assign tmp8786 = s3 ? tmp8787 : tmp8789;
  assign tmp8785 = s4 ? tmp8738 : tmp8786;
  assign tmp8793 = s2 ? tmp8756 : tmp8740;
  assign tmp8792 = s3 ? tmp8793 : tmp8759;
  assign tmp8796 = ~(s1 ? tmp7125 : tmp8740);
  assign tmp8795 = s2 ? tmp8763 : tmp8796;
  assign tmp8794 = ~(s3 ? tmp8795 : tmp8767);
  assign tmp8791 = s4 ? tmp8792 : tmp8794;
  assign tmp8800 = s1 ? tmp8772 : tmp7125;
  assign tmp8799 = s2 ? tmp8800 : 1;
  assign tmp8802 = s1 ? 1 : tmp8765;
  assign tmp8801 = ~(s2 ? 1 : tmp8802);
  assign tmp8798 = s3 ? tmp8799 : tmp8801;
  assign tmp8804 = s2 ? tmp7125 : tmp8740;
  assign tmp8805 = s1 ? tmp7125 : tmp8740;
  assign tmp8803 = s3 ? tmp8804 : tmp8805;
  assign tmp8797 = s4 ? tmp8798 : tmp8803;
  assign tmp8790 = s5 ? tmp8791 : tmp8797;
  assign tmp8784 = s6 ? tmp8785 : tmp8790;
  assign tmp8735 = s7 ? tmp8736 : tmp8784;
  assign tmp8809 = s3 ? tmp7952 : tmp8165;
  assign tmp8811 = s2 ? tmp8120 : tmp7955;
  assign tmp8814 = s0 ? tmp7948 : tmp7952;
  assign tmp8813 = s1 ? tmp7952 : tmp8814;
  assign tmp8812 = s2 ? tmp7962 : tmp8813;
  assign tmp8810 = s3 ? tmp8811 : tmp8812;
  assign tmp8808 = s4 ? tmp8809 : tmp8810;
  assign tmp8818 = s2 ? tmp7980 : tmp8018;
  assign tmp8817 = s3 ? tmp8131 : tmp8818;
  assign tmp8822 = s0 ? 1 : tmp7989;
  assign tmp8821 = s1 ? tmp8822 : tmp7978;
  assign tmp8823 = ~(s1 ? tmp7980 : tmp7955);
  assign tmp8820 = s2 ? tmp8821 : tmp8823;
  assign tmp8826 = s0 ? tmp7952 : tmp8740;
  assign tmp8825 = s1 ? tmp7952 : tmp8826;
  assign tmp8824 = ~(s2 ? tmp8825 : 0);
  assign tmp8819 = ~(s3 ? tmp8820 : tmp8824);
  assign tmp8816 = s4 ? tmp8817 : tmp8819;
  assign tmp8830 = s1 ? tmp8124 : tmp7988;
  assign tmp8829 = s2 ? tmp8830 : tmp7990;
  assign tmp8828 = s3 ? tmp8829 : tmp8773;
  assign tmp8833 = s1 ? tmp8778 : tmp7994;
  assign tmp8834 = ~(s1 ? tmp8822 : 0);
  assign tmp8832 = s2 ? tmp8833 : tmp8834;
  assign tmp8836 = s1 ? tmp7983 : tmp8782;
  assign tmp8835 = s2 ? tmp8836 : tmp8783;
  assign tmp8831 = s3 ? tmp8832 : tmp8835;
  assign tmp8827 = s4 ? tmp8828 : tmp8831;
  assign tmp8815 = s5 ? tmp8816 : tmp8827;
  assign tmp8807 = s6 ? tmp8808 : tmp8815;
  assign tmp8840 = s2 ? tmp8004 : tmp8813;
  assign tmp8839 = s3 ? tmp8120 : tmp8840;
  assign tmp8838 = s4 ? tmp8809 : tmp8839;
  assign tmp8844 = s2 ? tmp7952 : tmp8018;
  assign tmp8843 = s3 ? tmp8163 : tmp8844;
  assign tmp8846 = s2 ? tmp8821 : tmp7989;
  assign tmp8848 = s1 ? tmp7952 : tmp8740;
  assign tmp8847 = ~(s2 ? tmp8848 : 0);
  assign tmp8845 = ~(s3 ? tmp8846 : tmp8847);
  assign tmp8842 = s4 ? tmp8843 : tmp8845;
  assign tmp8852 = s1 ? tmp8124 : tmp7952;
  assign tmp8851 = s2 ? tmp8852 : 1;
  assign tmp8850 = s3 ? tmp8851 : tmp8801;
  assign tmp8854 = s2 ? tmp8021 : tmp7952;
  assign tmp8853 = s3 ? tmp8854 : tmp8805;
  assign tmp8849 = s4 ? tmp8850 : tmp8853;
  assign tmp8841 = s5 ? tmp8842 : tmp8849;
  assign tmp8837 = s6 ? tmp8838 : tmp8841;
  assign tmp8806 = s7 ? tmp8807 : tmp8837;
  assign tmp8734 = s8 ? tmp8735 : tmp8806;
  assign tmp8855 = s8 ? tmp8806 : tmp8023;
  assign tmp8733 = s9 ? tmp8734 : tmp8855;
  assign tmp8863 = s2 ? tmp8763 : tmp8765;
  assign tmp8864 = ~(s2 ? tmp8740 : 0);
  assign tmp8862 = ~(s3 ? tmp8863 : tmp8864);
  assign tmp8861 = s4 ? tmp8792 : tmp8862;
  assign tmp8860 = s5 ? tmp8861 : tmp8797;
  assign tmp8859 = s6 ? tmp8785 : tmp8860;
  assign tmp8858 = s7 ? tmp8736 : tmp8859;
  assign tmp8857 = s8 ? tmp8858 : tmp8736;
  assign tmp8870 = ~(s3 ? tmp8795 : tmp8864);
  assign tmp8869 = s4 ? tmp8792 : tmp8870;
  assign tmp8868 = s5 ? tmp8869 : tmp8797;
  assign tmp8867 = s6 ? tmp8785 : tmp8868;
  assign tmp8866 = s7 ? tmp8867 : tmp8024;
  assign tmp8871 = s7 ? tmp8837 : tmp8859;
  assign tmp8865 = s8 ? tmp8866 : tmp8871;
  assign tmp8856 = s9 ? tmp8857 : tmp8865;
  assign tmp8732 = s10 ? tmp8733 : tmp8856;
  assign tmp8875 = s7 ? tmp8784 : tmp8024;
  assign tmp8874 = s8 ? tmp8875 : tmp8871;
  assign tmp8873 = s9 ? tmp8857 : tmp8874;
  assign tmp8872 = s10 ? tmp8733 : tmp8873;
  assign tmp8731 = s11 ? tmp8732 : tmp8872;
  assign tmp8883 = s2 ? tmp8055 : tmp8061;
  assign tmp8882 = ~(s3 ? tmp8883 : tmp8062);
  assign tmp8881 = s4 ? tmp8050 : tmp8882;
  assign tmp8887 = s2 ? tmp8655 : tmp8100;
  assign tmp8886 = s3 ? tmp8887 : tmp8070;
  assign tmp8890 = s1 ? tmp7124 : 0;
  assign tmp8891 = ~(s1 ? 1 : tmp8648);
  assign tmp8889 = s2 ? tmp8890 : tmp8891;
  assign tmp8888 = s3 ? tmp8889 : tmp8077;
  assign tmp8885 = s4 ? tmp8886 : tmp8888;
  assign tmp8884 = ~(s5 ? tmp8885 : tmp8080);
  assign tmp8880 = s6 ? tmp8881 : tmp8884;
  assign tmp8894 = ~(s3 ? tmp8883 : tmp8095);
  assign tmp8893 = s4 ? tmp8050 : tmp8894;
  assign tmp8897 = s3 ? tmp8887 : tmp8101;
  assign tmp8899 = s2 ? tmp8890 : tmp7122;
  assign tmp8898 = s3 ? tmp8899 : tmp8105;
  assign tmp8896 = s4 ? tmp8897 : tmp8898;
  assign tmp8895 = ~(s5 ? tmp8896 : tmp8106);
  assign tmp8892 = s6 ? tmp8893 : tmp8895;
  assign tmp8879 = s7 ? tmp8880 : tmp8892;
  assign tmp8905 = s2 ? tmp7122 : tmp8061;
  assign tmp8904 = ~(s3 ? tmp8905 : tmp8062);
  assign tmp8903 = s4 ? tmp8218 : tmp8904;
  assign tmp8909 = s2 ? tmp8655 : tmp7122;
  assign tmp8908 = s3 ? tmp8909 : tmp8101;
  assign tmp8911 = s2 ? tmp8890 : tmp8561;
  assign tmp8910 = s3 ? tmp8911 : tmp8077;
  assign tmp8907 = s4 ? tmp8908 : tmp8910;
  assign tmp8906 = ~(s5 ? tmp8907 : tmp8080);
  assign tmp8902 = s6 ? tmp8903 : tmp8906;
  assign tmp8914 = ~(s3 ? tmp8905 : tmp8095);
  assign tmp8913 = s4 ? tmp8218 : tmp8914;
  assign tmp8916 = s4 ? tmp8908 : tmp8898;
  assign tmp8915 = ~(s5 ? tmp8916 : tmp8106);
  assign tmp8912 = s6 ? tmp8913 : tmp8915;
  assign tmp8901 = s7 ? tmp8902 : tmp8912;
  assign tmp8921 = ~(s2 ? tmp7125 : tmp7632);
  assign tmp8920 = s3 ? tmp7230 : tmp8921;
  assign tmp8923 = s2 ? tmp7125 : tmp7392;
  assign tmp8922 = ~(s3 ? tmp8923 : tmp8186);
  assign tmp8919 = s4 ? tmp8920 : tmp8922;
  assign tmp8926 = s3 ? tmp7226 : tmp8684;
  assign tmp8927 = s3 ? tmp8534 : tmp8193;
  assign tmp8925 = s4 ? tmp8926 : tmp8927;
  assign tmp8930 = s2 ? tmp8197 : tmp7125;
  assign tmp8929 = s3 ? tmp8930 : tmp7261;
  assign tmp8932 = s2 ? tmp7236 : tmp7242;
  assign tmp8931 = s3 ? tmp8932 : tmp8201;
  assign tmp8928 = s4 ? tmp8929 : tmp8931;
  assign tmp8924 = ~(s5 ? tmp8925 : tmp8928);
  assign tmp8918 = s6 ? tmp8919 : tmp8924;
  assign tmp8935 = ~(s3 ? tmp8923 : tmp8205);
  assign tmp8934 = s4 ? tmp8920 : tmp8935;
  assign tmp8938 = s3 ? tmp7226 : tmp7248;
  assign tmp8939 = s3 ? tmp7935 : tmp7450;
  assign tmp8937 = s4 ? tmp8938 : tmp8939;
  assign tmp8941 = s3 ? tmp8373 : tmp7261;
  assign tmp8940 = s4 ? tmp8941 : tmp7125;
  assign tmp8936 = ~(s5 ? tmp8937 : tmp8940);
  assign tmp8933 = s6 ? tmp8934 : tmp8936;
  assign tmp8917 = s7 ? tmp8918 : tmp8933;
  assign tmp8900 = s8 ? tmp8901 : tmp8917;
  assign tmp8878 = s9 ? tmp8879 : tmp8900;
  assign tmp8948 = ~(s2 ? tmp7122 : tmp8055);
  assign tmp8947 = s3 ? tmp8051 : tmp8948;
  assign tmp8946 = s4 ? tmp8947 : tmp8904;
  assign tmp8952 = s2 ? tmp7122 : tmp8100;
  assign tmp8951 = s3 ? tmp8952 : tmp8070;
  assign tmp8950 = s4 ? tmp8951 : tmp8910;
  assign tmp8955 = s2 ? tmp8083 : tmp8712;
  assign tmp8954 = s3 ? tmp8955 : tmp8084;
  assign tmp8957 = s2 ? tmp7170 : tmp8054;
  assign tmp8956 = s3 ? tmp8957 : tmp8089;
  assign tmp8953 = s4 ? tmp8954 : tmp8956;
  assign tmp8949 = ~(s5 ? tmp8950 : tmp8953);
  assign tmp8945 = s6 ? tmp8946 : tmp8949;
  assign tmp8959 = s4 ? tmp8947 : tmp8914;
  assign tmp8962 = s3 ? tmp8952 : tmp8101;
  assign tmp8961 = s4 ? tmp8962 : tmp8898;
  assign tmp8965 = s2 ? tmp7170 : tmp8091;
  assign tmp8964 = s3 ? tmp8965 : tmp8109;
  assign tmp8963 = s4 ? tmp8964 : tmp8110;
  assign tmp8960 = ~(s5 ? tmp8961 : tmp8963);
  assign tmp8958 = s6 ? tmp8959 : tmp8960;
  assign tmp8944 = s7 ? tmp8945 : tmp8958;
  assign tmp8943 = s8 ? tmp8944 : tmp8945;
  assign tmp8969 = ~(s5 ? tmp8896 : tmp8248);
  assign tmp8968 = s6 ? tmp8893 : tmp8969;
  assign tmp8967 = s7 ? tmp8968 : tmp8933;
  assign tmp8972 = s4 ? tmp8964 : tmp8243;
  assign tmp8971 = ~(s5 ? tmp8961 : tmp8972);
  assign tmp8970 = s6 ? tmp8959 : tmp8971;
  assign tmp8966 = s8 ? tmp8967 : tmp8970;
  assign tmp8942 = s9 ? tmp8943 : tmp8966;
  assign tmp8877 = s10 ? tmp8878 : tmp8942;
  assign tmp8976 = s7 ? tmp8892 : tmp8933;
  assign tmp8975 = s8 ? tmp8976 : tmp8958;
  assign tmp8974 = s9 ? tmp8943 : tmp8975;
  assign tmp8973 = s10 ? tmp8878 : tmp8974;
  assign tmp8876 = ~(s11 ? tmp8877 : tmp8973);
  assign tmp8730 = s12 ? tmp8731 : tmp8876;
  assign tmp8729 = s13 ? tmp8730 : tmp8255;
  assign tmp8728 = s14 ? tmp7774 : tmp8729;
  assign tmp8421 = s15 ? tmp8422 : tmp8728;
  assign tmp7109 = s16 ? tmp7110 : tmp8421;
  assign tmp8984 = s8 ? tmp8428 : tmp7215;
  assign tmp8983 = s9 ? tmp8427 : tmp8984;
  assign tmp8987 = s7 ? tmp8448 : tmp7265;
  assign tmp8986 = s8 ? tmp7270 : tmp8987;
  assign tmp8985 = s9 ? tmp7263 : tmp8986;
  assign tmp8982 = s10 ? tmp8983 : tmp8985;
  assign tmp8991 = s7 ? tmp8429 : tmp7265;
  assign tmp8990 = s8 ? tmp7281 : tmp8991;
  assign tmp8989 = s9 ? tmp7263 : tmp8990;
  assign tmp8988 = s10 ? tmp8983 : tmp8989;
  assign tmp8981 = s11 ? tmp8982 : tmp8988;
  assign tmp9000 = s3 ? tmp7444 : tmp8495;
  assign tmp8999 = s4 ? tmp7125 : tmp9000;
  assign tmp8998 = s6 ? tmp8999 : tmp8472;
  assign tmp8997 = s7 ? tmp8462 : tmp8998;
  assign tmp8996 = s8 ? tmp8476 : tmp8997;
  assign tmp8995 = s9 ? tmp8460 : tmp8996;
  assign tmp9002 = s8 ? tmp8997 : tmp8462;
  assign tmp9004 = s7 ? tmp8492 : tmp8998;
  assign tmp9005 = s7 ? tmp8496 : tmp8998;
  assign tmp9003 = s8 ? tmp9004 : tmp9005;
  assign tmp9001 = s9 ? tmp9002 : tmp9003;
  assign tmp8994 = s10 ? tmp8995 : tmp9001;
  assign tmp9009 = s7 ? tmp8471 : tmp8998;
  assign tmp9010 = s7 ? tmp8484 : tmp8998;
  assign tmp9008 = s8 ? tmp9009 : tmp9010;
  assign tmp9007 = s9 ? tmp9002 : tmp9008;
  assign tmp9006 = s10 ? tmp8995 : tmp9007;
  assign tmp8993 = s11 ? tmp8994 : tmp9006;
  assign tmp8992 = s12 ? tmp7283 : tmp8993;
  assign tmp8980 = s13 ? tmp8981 : tmp8992;
  assign tmp9016 = ~(s8 ? tmp8527 : 0);
  assign tmp9015 = s9 ? tmp8508 : tmp9016;
  assign tmp9020 = s6 ? tmp7332 : tmp8531;
  assign tmp9019 = ~(s7 ? tmp9020 : 0);
  assign tmp9018 = s8 ? 1 : tmp9019;
  assign tmp9017 = s9 ? 1 : tmp9018;
  assign tmp9014 = s10 ? tmp9015 : tmp9017;
  assign tmp9024 = ~(s7 ? tmp8519 : 0);
  assign tmp9023 = s8 ? 1 : tmp9024;
  assign tmp9022 = s9 ? 1 : tmp9023;
  assign tmp9021 = s10 ? tmp9015 : tmp9022;
  assign tmp9013 = s11 ? tmp9014 : tmp9021;
  assign tmp9034 = s2 ? tmp7222 : tmp7578;
  assign tmp9033 = s3 ? tmp8377 : tmp9034;
  assign tmp9032 = s4 ? tmp9033 : tmp7579;
  assign tmp9031 = s5 ? tmp9032 : tmp7581;
  assign tmp9030 = s6 ? tmp7570 : tmp9031;
  assign tmp9038 = s3 ? tmp8391 : tmp7577;
  assign tmp9037 = s4 ? tmp9038 : tmp7579;
  assign tmp9036 = s5 ? tmp9037 : tmp7598;
  assign tmp9035 = s6 ? tmp7592 : tmp9036;
  assign tmp9029 = s7 ? tmp9030 : tmp9035;
  assign tmp9028 = ~(s8 ? tmp8591 : tmp9029);
  assign tmp9027 = s9 ? tmp8543 : tmp9028;
  assign tmp9040 = s8 ? tmp7549 : tmp7550;
  assign tmp9043 = ~(s6 ? tmp7592 : tmp9036);
  assign tmp9042 = s7 ? tmp8615 : tmp9043;
  assign tmp9045 = s6 ? tmp8575 : tmp8620;
  assign tmp9046 = ~(s6 ? tmp7531 : tmp7559);
  assign tmp9044 = ~(s7 ? tmp9045 : tmp9046);
  assign tmp9041 = s8 ? tmp9042 : tmp9044;
  assign tmp9039 = s9 ? tmp9040 : tmp9041;
  assign tmp9026 = s10 ? tmp9027 : tmp9039;
  assign tmp9050 = s7 ? tmp8545 : tmp9043;
  assign tmp9051 = ~(s7 ? tmp8574 : tmp9046);
  assign tmp9049 = s8 ? tmp9050 : tmp9051;
  assign tmp9048 = s9 ? tmp9040 : tmp9049;
  assign tmp9047 = s10 ? tmp9027 : tmp9048;
  assign tmp9025 = s11 ? tmp9026 : tmp9047;
  assign tmp9012 = s12 ? tmp9013 : tmp9025;
  assign tmp9059 = s3 ? tmp7125 : tmp7256;
  assign tmp9058 = s4 ? tmp7639 : tmp9059;
  assign tmp9062 = s2 ? tmp7135 : tmp7242;
  assign tmp9061 = s3 ? tmp9062 : 1;
  assign tmp9060 = s4 ? tmp9061 : tmp7260;
  assign tmp9057 = s5 ? tmp9058 : tmp9060;
  assign tmp9056 = s6 ? tmp7629 : tmp9057;
  assign tmp9065 = s4 ? tmp7650 : tmp9059;
  assign tmp9067 = s3 ? tmp8394 : tmp7654;
  assign tmp9066 = s4 ? tmp9067 : tmp7260;
  assign tmp9064 = s5 ? tmp9065 : tmp9066;
  assign tmp9063 = s6 ? tmp7646 : tmp9064;
  assign tmp9055 = s7 ? tmp9056 : tmp9063;
  assign tmp9073 = s3 ? tmp7135 : 1;
  assign tmp9072 = s4 ? tmp9073 : tmp7260;
  assign tmp9071 = s5 ? tmp9065 : tmp9072;
  assign tmp9070 = s6 ? tmp7646 : tmp9071;
  assign tmp9069 = s7 ? tmp9056 : tmp9070;
  assign tmp9068 = s8 ? tmp9055 : tmp9069;
  assign tmp9054 = s9 ? tmp9055 : tmp9068;
  assign tmp9080 = s3 ? tmp7135 : tmp7654;
  assign tmp9079 = s4 ? tmp9080 : tmp7260;
  assign tmp9078 = s5 ? tmp9065 : tmp9079;
  assign tmp9077 = s6 ? tmp7646 : tmp9078;
  assign tmp9076 = s7 ? tmp9056 : tmp9077;
  assign tmp9075 = s8 ? tmp9076 : tmp9056;
  assign tmp9081 = s7 ? tmp9063 : tmp9077;
  assign tmp9074 = s9 ? tmp9075 : tmp9081;
  assign tmp9053 = s10 ? tmp9054 : tmp9074;
  assign tmp9052 = ~(s12 ? tmp9053 : tmp7745);
  assign tmp9011 = ~(s13 ? tmp9012 : tmp9052);
  assign tmp8979 = s14 ? tmp8980 : tmp9011;
  assign tmp9091 = s4 ? tmp8182 : tmp8922;
  assign tmp9094 = s3 ? tmp8394 : tmp7248;
  assign tmp9093 = s4 ? tmp9094 : tmp8927;
  assign tmp9092 = ~(s5 ? tmp9093 : tmp8194);
  assign tmp9090 = s6 ? tmp9091 : tmp9092;
  assign tmp9096 = s4 ? tmp8182 : tmp8935;
  assign tmp9098 = s4 ? tmp9094 : tmp8939;
  assign tmp9097 = ~(s5 ? tmp9098 : tmp8210);
  assign tmp9095 = s6 ? tmp9096 : tmp9097;
  assign tmp9089 = s7 ? tmp9090 : tmp9095;
  assign tmp9088 = s8 ? tmp8901 : tmp9089;
  assign tmp9087 = s9 ? tmp8879 : tmp9088;
  assign tmp9103 = ~(s5 ? tmp8916 : tmp8240);
  assign tmp9102 = s6 ? tmp8913 : tmp9103;
  assign tmp9101 = s7 ? tmp8902 : tmp9102;
  assign tmp9100 = s8 ? tmp9101 : tmp8902;
  assign tmp9105 = s7 ? tmp8968 : tmp9095;
  assign tmp9108 = ~(s5 ? tmp8916 : tmp8248);
  assign tmp9107 = s6 ? tmp8913 : tmp9108;
  assign tmp9106 = s7 ? tmp9107 : tmp9102;
  assign tmp9104 = s8 ? tmp9105 : tmp9106;
  assign tmp9099 = s9 ? tmp9100 : tmp9104;
  assign tmp9086 = s10 ? tmp9087 : tmp9099;
  assign tmp9112 = s7 ? tmp8892 : tmp9095;
  assign tmp9113 = s7 ? tmp8912 : tmp9102;
  assign tmp9111 = s8 ? tmp9112 : tmp9113;
  assign tmp9110 = s9 ? tmp9100 : tmp9111;
  assign tmp9109 = s10 ? tmp9087 : tmp9110;
  assign tmp9085 = ~(s11 ? tmp9086 : tmp9109);
  assign tmp9084 = s12 ? tmp7910 : tmp9085;
  assign tmp9083 = s13 ? tmp9084 : tmp8255;
  assign tmp9082 = s14 ? tmp7774 : tmp9083;
  assign tmp8978 = s15 ? tmp8979 : tmp9082;
  assign tmp9123 = s3 ? tmp7125 : tmp7794;
  assign tmp9122 = s4 ? tmp8683 : tmp9123;
  assign tmp9121 = s5 ? tmp9122 : tmp8686;
  assign tmp9120 = s6 ? tmp8678 : tmp9121;
  assign tmp9126 = s4 ? tmp8694 : tmp9059;
  assign tmp9128 = s3 ? tmp7125 : tmp7654;
  assign tmp9127 = s4 ? tmp9128 : tmp8687;
  assign tmp9125 = s5 ? tmp9126 : tmp9127;
  assign tmp9124 = s6 ? tmp8690 : tmp9125;
  assign tmp9119 = s7 ? tmp9120 : tmp9124;
  assign tmp9130 = s8 ? tmp9119 : tmp9120;
  assign tmp9129 = s9 ? tmp9130 : tmp9124;
  assign tmp9118 = s10 ? tmp9119 : tmp9129;
  assign tmp9117 = ~(s12 ? tmp9118 : tmp7745);
  assign tmp9116 = ~(s13 ? tmp8504 : tmp9117);
  assign tmp9115 = s14 ? tmp8423 : tmp9116;
  assign tmp9133 = s12 ? tmp7910 : tmp8876;
  assign tmp9132 = s13 ? tmp9133 : tmp8255;
  assign tmp9131 = s14 ? tmp7774 : tmp9132;
  assign tmp9114 = s15 ? tmp9115 : tmp9131;
  assign tmp8977 = s16 ? tmp8978 : tmp9114;
  assign tmp7108 = s17 ? tmp7109 : tmp8977;
  assign l1__1 = tmp7108;

  assign tmp9149 = ~(l2 ? 1 : 0);
  assign tmp9148 = l1 ? 1 : tmp9149;
  assign tmp9151 = l1 ? 1 : 0;
  assign tmp9150 = s0 ? tmp9151 : tmp9148;
  assign tmp9147 = s1 ? tmp9148 : tmp9150;
  assign tmp9154 = s0 ? tmp9148 : tmp9151;
  assign tmp9153 = s1 ? tmp9154 : tmp9148;
  assign tmp9152 = s2 ? tmp9148 : tmp9153;
  assign tmp9146 = s3 ? tmp9147 : tmp9152;
  assign tmp9158 = s0 ? tmp9148 : 1;
  assign tmp9159 = s0 ? tmp9151 : 1;
  assign tmp9157 = s1 ? tmp9158 : tmp9159;
  assign tmp9156 = s2 ? tmp9153 : tmp9157;
  assign tmp9161 = s1 ? tmp9151 : 1;
  assign tmp9163 = s0 ? tmp9148 : tmp9149;
  assign tmp9164 = s0 ? 1 : tmp9148;
  assign tmp9162 = s1 ? tmp9163 : tmp9164;
  assign tmp9160 = s2 ? tmp9161 : tmp9162;
  assign tmp9155 = s3 ? tmp9156 : tmp9160;
  assign tmp9145 = s4 ? tmp9146 : tmp9155;
  assign tmp9169 = s1 ? tmp9154 : tmp9150;
  assign tmp9172 = l2 ? 1 : 0;
  assign tmp9171 = ~(s0 ? tmp9172 : 1);
  assign tmp9170 = s1 ? tmp9150 : tmp9171;
  assign tmp9168 = s2 ? tmp9169 : tmp9170;
  assign tmp9174 = s0 ? 1 : tmp9172;
  assign tmp9175 = ~(s1 ? 1 : tmp9158);
  assign tmp9173 = ~(s2 ? tmp9174 : tmp9175);
  assign tmp9167 = s3 ? tmp9168 : tmp9173;
  assign tmp9178 = s1 ? tmp9164 : tmp9159;
  assign tmp9179 = s1 ? tmp9159 : tmp9154;
  assign tmp9177 = s2 ? tmp9178 : tmp9179;
  assign tmp9181 = s1 ? tmp9172 : 0;
  assign tmp9180 = ~(s2 ? tmp9181 : 0);
  assign tmp9176 = s3 ? tmp9177 : tmp9180;
  assign tmp9166 = s4 ? tmp9167 : tmp9176;
  assign tmp9186 = s0 ? tmp9172 : 0;
  assign tmp9185 = s1 ? tmp9186 : 0;
  assign tmp9188 = s0 ? 1 : tmp9149;
  assign tmp9187 = ~(s1 ? tmp9188 : tmp9149);
  assign tmp9184 = s2 ? tmp9185 : tmp9187;
  assign tmp9183 = s3 ? tmp9184 : 0;
  assign tmp9191 = s1 ? tmp9188 : tmp9149;
  assign tmp9190 = s2 ? 1 : tmp9191;
  assign tmp9189 = ~(s3 ? tmp9190 : 1);
  assign tmp9182 = ~(s4 ? tmp9183 : tmp9189);
  assign tmp9165 = s5 ? tmp9166 : tmp9182;
  assign tmp9144 = s6 ? tmp9145 : tmp9165;
  assign tmp9196 = s1 ? tmp9158 : tmp9151;
  assign tmp9195 = s2 ? tmp9153 : tmp9196;
  assign tmp9194 = s3 ? tmp9195 : tmp9160;
  assign tmp9193 = s4 ? tmp9146 : tmp9194;
  assign tmp9201 = s1 ? tmp9148 : tmp9171;
  assign tmp9200 = s2 ? tmp9153 : tmp9201;
  assign tmp9202 = ~(s2 ? tmp9172 : tmp9175);
  assign tmp9199 = s3 ? tmp9200 : tmp9202;
  assign tmp9205 = s1 ? tmp9151 : tmp9154;
  assign tmp9204 = s2 ? tmp9178 : tmp9205;
  assign tmp9203 = s3 ? tmp9204 : tmp9180;
  assign tmp9198 = s4 ? tmp9199 : tmp9203;
  assign tmp9208 = s2 ? tmp9185 : tmp9181;
  assign tmp9207 = s3 ? tmp9208 : 0;
  assign tmp9210 = s2 ? 1 : tmp9149;
  assign tmp9209 = ~(s3 ? tmp9210 : 1);
  assign tmp9206 = ~(s4 ? tmp9207 : tmp9209);
  assign tmp9197 = s5 ? tmp9198 : tmp9206;
  assign tmp9192 = s6 ? tmp9193 : tmp9197;
  assign tmp9143 = s7 ? tmp9144 : tmp9192;
  assign tmp9216 = s1 ? tmp9148 : tmp9164;
  assign tmp9215 = s2 ? tmp9161 : tmp9216;
  assign tmp9214 = s3 ? tmp9156 : tmp9215;
  assign tmp9213 = s4 ? tmp9146 : tmp9214;
  assign tmp9221 = s1 ? tmp9150 : tmp9154;
  assign tmp9220 = s2 ? tmp9169 : tmp9221;
  assign tmp9224 = s0 ? tmp9151 : tmp9149;
  assign tmp9223 = s1 ? tmp9150 : tmp9224;
  assign tmp9225 = s1 ? 1 : tmp9158;
  assign tmp9222 = s2 ? tmp9223 : tmp9225;
  assign tmp9219 = s3 ? tmp9220 : tmp9222;
  assign tmp9227 = ~(s2 ? tmp9185 : 0);
  assign tmp9226 = s3 ? tmp9177 : tmp9227;
  assign tmp9218 = s4 ? tmp9219 : tmp9226;
  assign tmp9217 = s5 ? tmp9218 : tmp9182;
  assign tmp9212 = s6 ? tmp9213 : tmp9217;
  assign tmp9230 = s3 ? tmp9195 : tmp9215;
  assign tmp9229 = s4 ? tmp9146 : tmp9230;
  assign tmp9235 = s1 ? tmp9148 : tmp9154;
  assign tmp9234 = s2 ? tmp9153 : tmp9235;
  assign tmp9237 = s1 ? tmp9148 : tmp9149;
  assign tmp9236 = s2 ? tmp9237 : tmp9225;
  assign tmp9233 = s3 ? tmp9234 : tmp9236;
  assign tmp9239 = s2 ? tmp9178 : tmp9148;
  assign tmp9238 = s3 ? tmp9239 : tmp9227;
  assign tmp9232 = s4 ? tmp9233 : tmp9238;
  assign tmp9231 = s5 ? tmp9232 : tmp9206;
  assign tmp9228 = s6 ? tmp9229 : tmp9231;
  assign tmp9211 = s7 ? tmp9212 : tmp9228;
  assign tmp9142 = s8 ? tmp9143 : tmp9211;
  assign tmp9245 = s2 ? tmp9151 : tmp9159;
  assign tmp9248 = s0 ? 1 : tmp9151;
  assign tmp9247 = s1 ? tmp9151 : tmp9248;
  assign tmp9246 = s2 ? tmp9161 : tmp9247;
  assign tmp9244 = s3 ? tmp9245 : tmp9246;
  assign tmp9243 = s4 ? tmp9151 : tmp9244;
  assign tmp9254 = s0 ? tmp9151 : 0;
  assign tmp9253 = s1 ? tmp9151 : tmp9254;
  assign tmp9252 = s2 ? tmp9151 : tmp9253;
  assign tmp9257 = ~(l1 ? 1 : 0);
  assign tmp9256 = s0 ? 1 : tmp9257;
  assign tmp9258 = ~(s1 ? 1 : tmp9159);
  assign tmp9255 = ~(s2 ? tmp9256 : tmp9258);
  assign tmp9251 = s3 ? tmp9252 : tmp9255;
  assign tmp9261 = s1 ? tmp9248 : tmp9159;
  assign tmp9262 = s1 ? tmp9159 : tmp9151;
  assign tmp9260 = s2 ? tmp9261 : tmp9262;
  assign tmp9263 = s2 ? tmp9151 : 1;
  assign tmp9259 = s3 ? tmp9260 : tmp9263;
  assign tmp9250 = s4 ? tmp9251 : tmp9259;
  assign tmp9267 = s1 ? tmp9159 : 1;
  assign tmp9268 = s1 ? tmp9248 : tmp9151;
  assign tmp9266 = s2 ? tmp9267 : tmp9268;
  assign tmp9265 = s3 ? tmp9266 : 1;
  assign tmp9270 = s2 ? 1 : tmp9268;
  assign tmp9269 = s3 ? tmp9270 : 1;
  assign tmp9264 = s4 ? tmp9265 : tmp9269;
  assign tmp9249 = s5 ? tmp9250 : tmp9264;
  assign tmp9242 = s6 ? tmp9243 : tmp9249;
  assign tmp9276 = s1 ? 1 : tmp9159;
  assign tmp9275 = s2 ? tmp9151 : tmp9276;
  assign tmp9274 = s3 ? tmp9252 : tmp9275;
  assign tmp9278 = s2 ? tmp9261 : tmp9151;
  assign tmp9279 = s2 ? tmp9161 : 1;
  assign tmp9277 = s3 ? tmp9278 : tmp9279;
  assign tmp9273 = s4 ? tmp9274 : tmp9277;
  assign tmp9282 = s2 ? tmp9267 : tmp9161;
  assign tmp9281 = s3 ? tmp9282 : 1;
  assign tmp9284 = s2 ? 1 : tmp9151;
  assign tmp9283 = s3 ? tmp9284 : 1;
  assign tmp9280 = s4 ? tmp9281 : tmp9283;
  assign tmp9272 = s5 ? tmp9273 : tmp9280;
  assign tmp9271 = s6 ? tmp9243 : tmp9272;
  assign tmp9241 = s7 ? tmp9242 : tmp9271;
  assign tmp9240 = s8 ? tmp9211 : tmp9241;
  assign tmp9141 = s9 ? tmp9142 : tmp9240;
  assign tmp9291 = s3 ? tmp9239 : tmp9180;
  assign tmp9290 = s4 ? tmp9199 : tmp9291;
  assign tmp9289 = s5 ? tmp9290 : tmp9206;
  assign tmp9288 = s6 ? tmp9193 : tmp9289;
  assign tmp9287 = s7 ? tmp9144 : tmp9288;
  assign tmp9286 = s8 ? tmp9287 : tmp9144;
  assign tmp9299 = s1 ? tmp9151 : tmp9148;
  assign tmp9298 = s2 ? tmp9178 : tmp9299;
  assign tmp9297 = s3 ? tmp9298 : tmp9180;
  assign tmp9296 = s4 ? tmp9199 : tmp9297;
  assign tmp9295 = s5 ? tmp9296 : tmp9206;
  assign tmp9294 = s6 ? tmp9193 : tmp9295;
  assign tmp9293 = s7 ? tmp9294 : tmp9271;
  assign tmp9300 = s7 ? tmp9228 : tmp9288;
  assign tmp9292 = s8 ? tmp9293 : tmp9300;
  assign tmp9285 = s9 ? tmp9286 : tmp9292;
  assign tmp9140 = s10 ? tmp9141 : tmp9285;
  assign tmp9304 = s7 ? tmp9192 : tmp9271;
  assign tmp9303 = s8 ? tmp9304 : tmp9300;
  assign tmp9302 = s9 ? tmp9286 : tmp9303;
  assign tmp9301 = s10 ? tmp9141 : tmp9302;
  assign tmp9139 = s11 ? tmp9140 : tmp9301;
  assign tmp9314 = s2 ? tmp9148 : tmp9158;
  assign tmp9317 = s0 ? 1 : 0;
  assign tmp9316 = s1 ? tmp9148 : tmp9317;
  assign tmp9320 = ~(l1 ? 1 : tmp9149);
  assign tmp9319 = ~(s0 ? 1 : tmp9320);
  assign tmp9318 = s1 ? tmp9148 : tmp9319;
  assign tmp9315 = s2 ? tmp9316 : tmp9318;
  assign tmp9313 = s3 ? tmp9314 : tmp9315;
  assign tmp9312 = s4 ? tmp9148 : tmp9313;
  assign tmp9326 = ~(s0 ? tmp9151 : 0);
  assign tmp9325 = s1 ? 1 : tmp9326;
  assign tmp9324 = ~(s2 ? tmp9172 : tmp9325);
  assign tmp9323 = s3 ? tmp9148 : tmp9324;
  assign tmp9329 = s1 ? tmp9256 : tmp9326;
  assign tmp9330 = ~(s1 ? tmp9254 : tmp9151);
  assign tmp9328 = s2 ? tmp9329 : tmp9330;
  assign tmp9327 = ~(s3 ? tmp9328 : 1);
  assign tmp9322 = s4 ? tmp9323 : tmp9327;
  assign tmp9321 = s5 ? tmp9322 : 0;
  assign tmp9311 = s6 ? tmp9312 : tmp9321;
  assign tmp9335 = s2 ? tmp9329 : tmp9257;
  assign tmp9334 = ~(s3 ? tmp9335 : 1);
  assign tmp9333 = s4 ? tmp9323 : tmp9334;
  assign tmp9332 = s5 ? tmp9333 : 0;
  assign tmp9331 = s6 ? tmp9312 : tmp9332;
  assign tmp9310 = s7 ? tmp9311 : tmp9331;
  assign tmp9343 = ~(s0 ? tmp9151 : 1);
  assign tmp9342 = ~(s1 ? 1 : tmp9343);
  assign tmp9341 = s2 ? tmp9148 : tmp9342;
  assign tmp9340 = s3 ? tmp9148 : tmp9341;
  assign tmp9346 = s1 ? tmp9256 : tmp9343;
  assign tmp9347 = ~(s1 ? tmp9159 : tmp9151);
  assign tmp9345 = s2 ? tmp9346 : tmp9347;
  assign tmp9350 = ~(s0 ? 1 : 0);
  assign tmp9349 = s1 ? tmp9317 : tmp9350;
  assign tmp9348 = s2 ? tmp9349 : 1;
  assign tmp9344 = ~(s3 ? tmp9345 : tmp9348);
  assign tmp9339 = s4 ? tmp9340 : tmp9344;
  assign tmp9338 = s5 ? tmp9339 : 0;
  assign tmp9337 = s6 ? tmp9312 : tmp9338;
  assign tmp9355 = s1 ? tmp9148 : 0;
  assign tmp9354 = s2 ? tmp9355 : tmp9318;
  assign tmp9353 = s3 ? tmp9314 : tmp9354;
  assign tmp9352 = s4 ? tmp9148 : tmp9353;
  assign tmp9359 = s2 ? tmp9346 : tmp9257;
  assign tmp9361 = s1 ? tmp9317 : 1;
  assign tmp9360 = s2 ? tmp9361 : 1;
  assign tmp9358 = ~(s3 ? tmp9359 : tmp9360);
  assign tmp9357 = s4 ? tmp9340 : tmp9358;
  assign tmp9356 = s5 ? tmp9357 : 0;
  assign tmp9351 = s6 ? tmp9352 : tmp9356;
  assign tmp9336 = s7 ? tmp9337 : tmp9351;
  assign tmp9309 = s8 ? tmp9310 : tmp9336;
  assign tmp9367 = ~(s3 ? tmp9345 : 1);
  assign tmp9366 = s4 ? tmp9323 : tmp9367;
  assign tmp9365 = s5 ? tmp9366 : 0;
  assign tmp9364 = s6 ? tmp9312 : tmp9365;
  assign tmp9371 = ~(s3 ? tmp9359 : 1);
  assign tmp9370 = s4 ? tmp9323 : tmp9371;
  assign tmp9369 = s5 ? tmp9370 : 0;
  assign tmp9368 = s6 ? tmp9352 : tmp9369;
  assign tmp9363 = s7 ? tmp9364 : tmp9368;
  assign tmp9362 = s8 ? tmp9336 : tmp9363;
  assign tmp9308 = s9 ? tmp9309 : tmp9362;
  assign tmp9373 = s8 ? tmp9363 : tmp9364;
  assign tmp9381 = s1 ? tmp9151 : tmp9149;
  assign tmp9380 = s2 ? tmp9148 : tmp9381;
  assign tmp9383 = s1 ? tmp9172 : 1;
  assign tmp9382 = ~(s2 ? tmp9383 : tmp9325);
  assign tmp9379 = s3 ? tmp9380 : tmp9382;
  assign tmp9378 = s4 ? tmp9379 : tmp9334;
  assign tmp9377 = s5 ? tmp9378 : 0;
  assign tmp9376 = s6 ? tmp9352 : tmp9377;
  assign tmp9387 = s3 ? tmp9380 : tmp9324;
  assign tmp9386 = s4 ? tmp9387 : tmp9371;
  assign tmp9385 = s5 ? tmp9386 : 0;
  assign tmp9384 = s6 ? tmp9352 : tmp9385;
  assign tmp9375 = s7 ? tmp9376 : tmp9384;
  assign tmp9393 = s2 ? tmp9148 : tmp9299;
  assign tmp9392 = s3 ? tmp9393 : tmp9341;
  assign tmp9391 = s4 ? tmp9392 : tmp9358;
  assign tmp9390 = s5 ? tmp9391 : 0;
  assign tmp9389 = s6 ? tmp9352 : tmp9390;
  assign tmp9388 = s7 ? tmp9389 : tmp9384;
  assign tmp9374 = s8 ? tmp9375 : tmp9388;
  assign tmp9372 = s9 ? tmp9373 : tmp9374;
  assign tmp9307 = s10 ? tmp9308 : tmp9372;
  assign tmp9397 = s7 ? tmp9331 : tmp9368;
  assign tmp9398 = s7 ? tmp9351 : tmp9368;
  assign tmp9396 = s8 ? tmp9397 : tmp9398;
  assign tmp9395 = s9 ? tmp9373 : tmp9396;
  assign tmp9394 = s10 ? tmp9308 : tmp9395;
  assign tmp9306 = s11 ? tmp9307 : tmp9394;
  assign tmp9305 = s12 ? tmp9306 : 1;
  assign tmp9138 = s13 ? tmp9139 : tmp9305;
  assign tmp9409 = s2 ? tmp9172 : tmp9186;
  assign tmp9411 = s1 ? tmp9172 : tmp9350;
  assign tmp9412 = s1 ? tmp9172 : tmp9174;
  assign tmp9410 = s2 ? tmp9411 : tmp9412;
  assign tmp9408 = s3 ? tmp9409 : tmp9410;
  assign tmp9407 = s4 ? tmp9172 : tmp9408;
  assign tmp9416 = s2 ? tmp9172 : 1;
  assign tmp9415 = s3 ? tmp9172 : tmp9416;
  assign tmp9414 = s4 ? tmp9415 : 1;
  assign tmp9413 = s5 ? tmp9414 : 1;
  assign tmp9406 = s6 ? tmp9407 : tmp9413;
  assign tmp9420 = s2 ? tmp9383 : tmp9412;
  assign tmp9419 = s3 ? tmp9409 : tmp9420;
  assign tmp9418 = s4 ? tmp9172 : tmp9419;
  assign tmp9425 = s1 ? 1 : tmp9172;
  assign tmp9424 = s2 ? tmp9172 : tmp9425;
  assign tmp9423 = s3 ? tmp9424 : tmp9416;
  assign tmp9422 = s4 ? tmp9423 : 1;
  assign tmp9421 = s5 ? tmp9422 : 1;
  assign tmp9417 = s6 ? tmp9418 : tmp9421;
  assign tmp9405 = s7 ? tmp9406 : tmp9417;
  assign tmp9433 = s0 ? tmp9172 : 1;
  assign tmp9432 = s1 ? tmp9433 : tmp9172;
  assign tmp9431 = s2 ? tmp9172 : tmp9432;
  assign tmp9430 = s3 ? tmp9431 : tmp9416;
  assign tmp9429 = s4 ? tmp9430 : 1;
  assign tmp9428 = s5 ? tmp9429 : 1;
  assign tmp9427 = s6 ? tmp9407 : tmp9428;
  assign tmp9426 = s7 ? tmp9427 : tmp9417;
  assign tmp9404 = s8 ? tmp9405 : tmp9426;
  assign tmp9403 = s9 ? tmp9404 : tmp9426;
  assign tmp9435 = s8 ? tmp9426 : tmp9427;
  assign tmp9442 = s2 ? tmp9383 : 1;
  assign tmp9441 = s3 ? tmp9424 : tmp9442;
  assign tmp9440 = s4 ? tmp9441 : 1;
  assign tmp9439 = s5 ? tmp9440 : 1;
  assign tmp9438 = s6 ? tmp9418 : tmp9439;
  assign tmp9437 = s7 ? tmp9438 : tmp9417;
  assign tmp9436 = s8 ? tmp9437 : tmp9417;
  assign tmp9434 = s9 ? tmp9435 : tmp9436;
  assign tmp9402 = s10 ? tmp9403 : tmp9434;
  assign tmp9444 = s9 ? tmp9435 : tmp9417;
  assign tmp9443 = s10 ? tmp9403 : tmp9444;
  assign tmp9401 = s11 ? tmp9402 : tmp9443;
  assign tmp9454 = ~(s0 ? tmp9151 : tmp9149);
  assign tmp9453 = s1 ? tmp9172 : tmp9454;
  assign tmp9456 = s1 ? tmp9186 : tmp9172;
  assign tmp9455 = s2 ? tmp9172 : tmp9456;
  assign tmp9452 = s3 ? tmp9453 : tmp9455;
  assign tmp9459 = s1 ? tmp9186 : tmp9343;
  assign tmp9458 = s2 ? tmp9456 : tmp9459;
  assign tmp9461 = s1 ? tmp9151 : tmp9317;
  assign tmp9462 = ~(s1 ? tmp9172 : tmp9174);
  assign tmp9460 = ~(s2 ? tmp9461 : tmp9462);
  assign tmp9457 = s3 ? tmp9458 : tmp9460;
  assign tmp9451 = s4 ? tmp9452 : tmp9457;
  assign tmp9465 = s3 ? tmp9184 : tmp9424;
  assign tmp9468 = s1 ? tmp9174 : tmp9257;
  assign tmp9470 = ~(s0 ? tmp9172 : 0);
  assign tmp9469 = ~(s1 ? tmp9151 : tmp9470);
  assign tmp9467 = s2 ? tmp9468 : tmp9469;
  assign tmp9471 = s2 ? tmp9453 : 1;
  assign tmp9466 = s3 ? tmp9467 : tmp9471;
  assign tmp9464 = s4 ? tmp9465 : tmp9466;
  assign tmp9475 = s1 ? tmp9433 : 1;
  assign tmp9476 = s1 ? tmp9317 : 0;
  assign tmp9474 = s2 ? tmp9475 : tmp9476;
  assign tmp9478 = ~(s1 ? 1 : tmp9174);
  assign tmp9477 = ~(s2 ? tmp9476 : tmp9478);
  assign tmp9473 = s3 ? tmp9474 : tmp9477;
  assign tmp9481 = s1 ? tmp9174 : 0;
  assign tmp9480 = s2 ? tmp9475 : tmp9481;
  assign tmp9483 = s1 ? 1 : tmp9174;
  assign tmp9484 = s1 ? tmp9174 : 1;
  assign tmp9482 = s2 ? tmp9483 : tmp9484;
  assign tmp9479 = s3 ? tmp9480 : tmp9482;
  assign tmp9472 = s4 ? tmp9473 : tmp9479;
  assign tmp9463 = s5 ? tmp9464 : tmp9472;
  assign tmp9450 = s6 ? tmp9451 : tmp9463;
  assign tmp9489 = s1 ? tmp9186 : tmp9257;
  assign tmp9488 = s2 ? tmp9456 : tmp9489;
  assign tmp9491 = s1 ? tmp9151 : 0;
  assign tmp9490 = ~(s2 ? tmp9491 : tmp9462);
  assign tmp9487 = s3 ? tmp9488 : tmp9490;
  assign tmp9486 = s4 ? tmp9452 : tmp9487;
  assign tmp9495 = s2 ? tmp9185 : tmp9172;
  assign tmp9494 = s3 ? tmp9495 : tmp9424;
  assign tmp9498 = ~(s1 ? tmp9151 : tmp9149);
  assign tmp9497 = s2 ? tmp9468 : tmp9498;
  assign tmp9496 = s3 ? tmp9497 : tmp9471;
  assign tmp9493 = s4 ? tmp9494 : tmp9496;
  assign tmp9501 = s2 ? tmp9475 : 0;
  assign tmp9502 = s2 ? 1 : tmp9425;
  assign tmp9500 = s3 ? tmp9501 : tmp9502;
  assign tmp9504 = s2 ? 1 : tmp9172;
  assign tmp9503 = s3 ? tmp9504 : tmp9425;
  assign tmp9499 = s4 ? tmp9500 : tmp9503;
  assign tmp9492 = s5 ? tmp9493 : tmp9499;
  assign tmp9485 = s6 ? tmp9486 : tmp9492;
  assign tmp9449 = s7 ? tmp9450 : tmp9485;
  assign tmp9511 = ~(s1 ? tmp9188 : tmp9470);
  assign tmp9510 = s2 ? tmp9185 : tmp9511;
  assign tmp9513 = ~(s1 ? 1 : tmp9172);
  assign tmp9512 = ~(s2 ? tmp9188 : tmp9513);
  assign tmp9509 = s3 ? tmp9510 : tmp9512;
  assign tmp9508 = s4 ? tmp9509 : tmp9466;
  assign tmp9507 = s5 ? tmp9508 : tmp9472;
  assign tmp9506 = s6 ? tmp9451 : tmp9507;
  assign tmp9519 = s1 ? tmp9172 : tmp9186;
  assign tmp9518 = s2 ? tmp9185 : tmp9519;
  assign tmp9517 = s3 ? tmp9518 : tmp9424;
  assign tmp9521 = s2 ? tmp9468 : tmp9172;
  assign tmp9520 = s3 ? tmp9521 : tmp9416;
  assign tmp9516 = s4 ? tmp9517 : tmp9520;
  assign tmp9515 = s5 ? tmp9516 : tmp9499;
  assign tmp9514 = s6 ? tmp9486 : tmp9515;
  assign tmp9505 = s7 ? tmp9506 : tmp9514;
  assign tmp9448 = s8 ? tmp9449 : tmp9505;
  assign tmp9527 = s2 ? tmp9151 : tmp9262;
  assign tmp9526 = s3 ? tmp9151 : tmp9527;
  assign tmp9531 = ~(s0 ? 1 : tmp9257);
  assign tmp9530 = s1 ? tmp9151 : tmp9531;
  assign tmp9529 = s2 ? tmp9461 : tmp9530;
  assign tmp9528 = s3 ? tmp9245 : tmp9529;
  assign tmp9525 = s4 ? tmp9526 : tmp9528;
  assign tmp9536 = ~(s1 ? 1 : tmp9257);
  assign tmp9535 = s2 ? tmp9151 : tmp9536;
  assign tmp9534 = s3 ? tmp9266 : tmp9535;
  assign tmp9539 = s1 ? tmp9256 : tmp9257;
  assign tmp9538 = s2 ? tmp9539 : tmp9257;
  assign tmp9540 = ~(s2 ? tmp9151 : 0);
  assign tmp9537 = ~(s3 ? tmp9538 : tmp9540);
  assign tmp9533 = s4 ? tmp9534 : tmp9537;
  assign tmp9544 = s1 ? tmp9254 : 0;
  assign tmp9545 = ~(s1 ? tmp9317 : 0);
  assign tmp9543 = s2 ? tmp9544 : tmp9545;
  assign tmp9547 = ~(s1 ? 1 : tmp9256);
  assign tmp9546 = s2 ? tmp9476 : tmp9547;
  assign tmp9542 = s3 ? tmp9543 : tmp9546;
  assign tmp9550 = ~(s1 ? tmp9256 : 0);
  assign tmp9549 = s2 ? tmp9544 : tmp9550;
  assign tmp9552 = s1 ? 1 : tmp9256;
  assign tmp9553 = s1 ? tmp9256 : 1;
  assign tmp9551 = ~(s2 ? tmp9552 : tmp9553);
  assign tmp9548 = s3 ? tmp9549 : tmp9551;
  assign tmp9541 = s4 ? tmp9542 : tmp9548;
  assign tmp9532 = s5 ? tmp9533 : tmp9541;
  assign tmp9524 = s6 ? tmp9525 : tmp9532;
  assign tmp9557 = s2 ? tmp9491 : tmp9530;
  assign tmp9556 = s3 ? tmp9245 : tmp9557;
  assign tmp9555 = s4 ? tmp9526 : tmp9556;
  assign tmp9561 = s2 ? tmp9267 : tmp9151;
  assign tmp9560 = s3 ? tmp9561 : tmp9535;
  assign tmp9559 = s4 ? tmp9560 : tmp9537;
  assign tmp9564 = s2 ? tmp9544 : 1;
  assign tmp9566 = s1 ? 1 : tmp9257;
  assign tmp9565 = ~(s2 ? 1 : tmp9566);
  assign tmp9563 = s3 ? tmp9564 : tmp9565;
  assign tmp9568 = s2 ? 1 : tmp9257;
  assign tmp9567 = ~(s3 ? tmp9568 : tmp9566);
  assign tmp9562 = s4 ? tmp9563 : tmp9567;
  assign tmp9558 = s5 ? tmp9559 : tmp9562;
  assign tmp9554 = s6 ? tmp9555 : tmp9558;
  assign tmp9523 = ~(s7 ? tmp9524 : tmp9554);
  assign tmp9522 = s8 ? tmp9505 : tmp9523;
  assign tmp9447 = s9 ? tmp9448 : tmp9522;
  assign tmp9574 = s4 ? tmp9494 : tmp9520;
  assign tmp9573 = s5 ? tmp9574 : tmp9499;
  assign tmp9572 = s6 ? tmp9486 : tmp9573;
  assign tmp9571 = s7 ? tmp9450 : tmp9572;
  assign tmp9570 = s8 ? tmp9571 : tmp9450;
  assign tmp9580 = s3 ? tmp9497 : tmp9416;
  assign tmp9579 = s4 ? tmp9494 : tmp9580;
  assign tmp9578 = s5 ? tmp9579 : tmp9499;
  assign tmp9577 = s6 ? tmp9486 : tmp9578;
  assign tmp9581 = ~(s6 ? tmp9555 : tmp9558);
  assign tmp9576 = s7 ? tmp9577 : tmp9581;
  assign tmp9582 = s7 ? tmp9514 : tmp9572;
  assign tmp9575 = s8 ? tmp9576 : tmp9582;
  assign tmp9569 = s9 ? tmp9570 : tmp9575;
  assign tmp9446 = s10 ? tmp9447 : tmp9569;
  assign tmp9586 = s7 ? tmp9485 : tmp9581;
  assign tmp9585 = s8 ? tmp9586 : tmp9582;
  assign tmp9584 = s9 ? tmp9570 : tmp9585;
  assign tmp9583 = s10 ? tmp9447 : tmp9584;
  assign tmp9445 = s11 ? tmp9446 : tmp9583;
  assign tmp9400 = s12 ? tmp9401 : tmp9445;
  assign tmp9595 = s3 ? tmp9453 : tmp9431;
  assign tmp9599 = s0 ? tmp9172 : tmp9257;
  assign tmp9598 = s1 ? tmp9599 : tmp9172;
  assign tmp9600 = s1 ? tmp9433 : tmp9326;
  assign tmp9597 = s2 ? tmp9598 : tmp9600;
  assign tmp9596 = s3 ? tmp9597 : tmp9490;
  assign tmp9594 = s4 ? tmp9595 : tmp9596;
  assign tmp9605 = s1 ? tmp9433 : tmp9174;
  assign tmp9606 = s1 ? tmp9174 : tmp9433;
  assign tmp9604 = s2 ? tmp9605 : tmp9606;
  assign tmp9610 = l1 ? tmp9172 : 0;
  assign tmp9609 = s0 ? tmp9172 : tmp9610;
  assign tmp9608 = s1 ? 1 : tmp9609;
  assign tmp9607 = s2 ? tmp9174 : tmp9608;
  assign tmp9603 = s3 ? tmp9604 : tmp9607;
  assign tmp9613 = s1 ? tmp9174 : tmp9343;
  assign tmp9615 = ~(s0 ? tmp9172 : tmp9257);
  assign tmp9614 = ~(s1 ? tmp9159 : tmp9615);
  assign tmp9612 = s2 ? tmp9613 : tmp9614;
  assign tmp9618 = ~(s0 ? 1 : tmp9149);
  assign tmp9617 = s1 ? tmp9609 : tmp9618;
  assign tmp9616 = s2 ? tmp9617 : 1;
  assign tmp9611 = s3 ? tmp9612 : tmp9616;
  assign tmp9602 = s4 ? tmp9603 : tmp9611;
  assign tmp9622 = s0 ? tmp9610 : tmp9172;
  assign tmp9621 = s2 ? tmp9475 : tmp9622;
  assign tmp9623 = s2 ? tmp9475 : tmp9483;
  assign tmp9620 = s3 ? tmp9621 : tmp9623;
  assign tmp9626 = s1 ? tmp9174 : tmp9609;
  assign tmp9625 = s2 ? tmp9172 : tmp9626;
  assign tmp9624 = s3 ? tmp9625 : tmp9482;
  assign tmp9619 = s4 ? tmp9620 : tmp9624;
  assign tmp9601 = s5 ? tmp9602 : tmp9619;
  assign tmp9593 = s6 ? tmp9594 : tmp9601;
  assign tmp9631 = s1 ? tmp9433 : tmp9257;
  assign tmp9630 = s2 ? tmp9598 : tmp9631;
  assign tmp9629 = s3 ? tmp9630 : tmp9490;
  assign tmp9628 = s4 ? tmp9595 : tmp9629;
  assign tmp9636 = s1 ? tmp9172 : tmp9433;
  assign tmp9635 = s2 ? tmp9432 : tmp9636;
  assign tmp9637 = s2 ? tmp9172 : tmp9608;
  assign tmp9634 = s3 ? tmp9635 : tmp9637;
  assign tmp9639 = s2 ? tmp9613 : tmp9172;
  assign tmp9641 = s1 ? tmp9609 : tmp9172;
  assign tmp9640 = s2 ? tmp9641 : 1;
  assign tmp9638 = s3 ? tmp9639 : tmp9640;
  assign tmp9633 = s4 ? tmp9634 : tmp9638;
  assign tmp9645 = s1 ? tmp9172 : tmp9622;
  assign tmp9644 = s2 ? tmp9475 : tmp9645;
  assign tmp9648 = s0 ? tmp9610 : 1;
  assign tmp9647 = s1 ? tmp9648 : 1;
  assign tmp9646 = s2 ? tmp9647 : tmp9425;
  assign tmp9643 = s3 ? tmp9644 : tmp9646;
  assign tmp9651 = s1 ? tmp9172 : tmp9609;
  assign tmp9650 = s2 ? 1 : tmp9651;
  assign tmp9649 = s3 ? tmp9650 : tmp9172;
  assign tmp9642 = s4 ? tmp9643 : tmp9649;
  assign tmp9632 = s5 ? tmp9633 : tmp9642;
  assign tmp9627 = s6 ? tmp9628 : tmp9632;
  assign tmp9592 = s7 ? tmp9593 : tmp9627;
  assign tmp9657 = l1 ? tmp9172 : 1;
  assign tmp9659 = ~(l1 ? tmp9172 : 1);
  assign tmp9658 = ~(s0 ? tmp9151 : tmp9659);
  assign tmp9656 = s1 ? tmp9657 : tmp9658;
  assign tmp9662 = s0 ? tmp9657 : 1;
  assign tmp9661 = s1 ? tmp9662 : tmp9657;
  assign tmp9660 = s2 ? tmp9657 : tmp9661;
  assign tmp9655 = s3 ? tmp9656 : tmp9660;
  assign tmp9666 = s0 ? tmp9657 : tmp9257;
  assign tmp9665 = s1 ? tmp9666 : tmp9657;
  assign tmp9667 = s1 ? tmp9662 : tmp9326;
  assign tmp9664 = s2 ? tmp9665 : tmp9667;
  assign tmp9670 = s0 ? 1 : tmp9657;
  assign tmp9669 = ~(s1 ? tmp9657 : tmp9670);
  assign tmp9668 = ~(s2 ? tmp9491 : tmp9669);
  assign tmp9663 = s3 ? tmp9664 : tmp9668;
  assign tmp9654 = s4 ? tmp9655 : tmp9663;
  assign tmp9675 = s1 ? tmp9662 : tmp9670;
  assign tmp9676 = s1 ? tmp9670 : tmp9662;
  assign tmp9674 = s2 ? tmp9675 : tmp9676;
  assign tmp9678 = s1 ? 1 : tmp9657;
  assign tmp9677 = s2 ? tmp9670 : tmp9678;
  assign tmp9673 = s3 ? tmp9674 : tmp9677;
  assign tmp9681 = s1 ? tmp9670 : tmp9257;
  assign tmp9683 = ~(s0 ? tmp9657 : tmp9257);
  assign tmp9682 = ~(s1 ? tmp9151 : tmp9683);
  assign tmp9680 = s2 ? tmp9681 : tmp9682;
  assign tmp9685 = s1 ? tmp9657 : tmp9454;
  assign tmp9684 = s2 ? tmp9685 : 1;
  assign tmp9679 = s3 ? tmp9680 : tmp9684;
  assign tmp9672 = s4 ? tmp9673 : tmp9679;
  assign tmp9689 = s1 ? tmp9662 : 1;
  assign tmp9691 = s0 ? tmp9172 : tmp9657;
  assign tmp9690 = s1 ? tmp9670 : tmp9691;
  assign tmp9688 = s2 ? tmp9689 : tmp9690;
  assign tmp9687 = s3 ? tmp9688 : tmp9623;
  assign tmp9695 = s0 ? tmp9657 : tmp9172;
  assign tmp9694 = s1 ? tmp9670 : tmp9695;
  assign tmp9693 = s2 ? tmp9383 : tmp9694;
  assign tmp9692 = s3 ? tmp9693 : tmp9482;
  assign tmp9686 = s4 ? tmp9687 : tmp9692;
  assign tmp9671 = s5 ? tmp9672 : tmp9686;
  assign tmp9653 = s6 ? tmp9654 : tmp9671;
  assign tmp9700 = s1 ? tmp9662 : tmp9257;
  assign tmp9699 = s2 ? tmp9665 : tmp9700;
  assign tmp9698 = s3 ? tmp9699 : tmp9668;
  assign tmp9697 = s4 ? tmp9655 : tmp9698;
  assign tmp9705 = s1 ? tmp9657 : tmp9662;
  assign tmp9704 = s2 ? tmp9661 : tmp9705;
  assign tmp9706 = s2 ? tmp9657 : tmp9678;
  assign tmp9703 = s3 ? tmp9704 : tmp9706;
  assign tmp9708 = s2 ? tmp9681 : tmp9657;
  assign tmp9710 = s1 ? tmp9657 : tmp9172;
  assign tmp9709 = s2 ? tmp9710 : 1;
  assign tmp9707 = s3 ? tmp9708 : tmp9709;
  assign tmp9702 = s4 ? tmp9703 : tmp9707;
  assign tmp9713 = s2 ? tmp9689 : tmp9710;
  assign tmp9712 = s3 ? tmp9713 : tmp9646;
  assign tmp9716 = s1 ? tmp9657 : tmp9610;
  assign tmp9715 = s2 ? 1 : tmp9716;
  assign tmp9714 = s3 ? tmp9715 : tmp9172;
  assign tmp9711 = s4 ? tmp9712 : tmp9714;
  assign tmp9701 = s5 ? tmp9702 : tmp9711;
  assign tmp9696 = s6 ? tmp9697 : tmp9701;
  assign tmp9652 = s7 ? tmp9653 : tmp9696;
  assign tmp9591 = s8 ? tmp9592 : tmp9652;
  assign tmp9724 = s1 ? 1 : tmp9695;
  assign tmp9723 = s2 ? tmp9670 : tmp9724;
  assign tmp9722 = s3 ? tmp9674 : tmp9723;
  assign tmp9727 = s1 ? tmp9670 : tmp9343;
  assign tmp9728 = ~(s1 ? tmp9159 : tmp9683);
  assign tmp9726 = s2 ? tmp9727 : tmp9728;
  assign tmp9730 = s1 ? tmp9695 : tmp9618;
  assign tmp9729 = s2 ? tmp9730 : 1;
  assign tmp9725 = s3 ? tmp9726 : tmp9729;
  assign tmp9721 = s4 ? tmp9722 : tmp9725;
  assign tmp9733 = s2 ? tmp9689 : tmp9691;
  assign tmp9732 = s3 ? tmp9733 : tmp9623;
  assign tmp9735 = s2 ? tmp9172 : tmp9694;
  assign tmp9734 = s3 ? tmp9735 : tmp9482;
  assign tmp9731 = s4 ? tmp9732 : tmp9734;
  assign tmp9720 = s5 ? tmp9721 : tmp9731;
  assign tmp9719 = s6 ? tmp9654 : tmp9720;
  assign tmp9740 = s2 ? tmp9657 : tmp9724;
  assign tmp9739 = s3 ? tmp9704 : tmp9740;
  assign tmp9742 = s2 ? tmp9727 : tmp9657;
  assign tmp9744 = s1 ? tmp9695 : tmp9172;
  assign tmp9743 = s2 ? tmp9744 : 1;
  assign tmp9741 = s3 ? tmp9742 : tmp9743;
  assign tmp9738 = s4 ? tmp9739 : tmp9741;
  assign tmp9747 = s2 ? tmp9475 : tmp9425;
  assign tmp9746 = s3 ? tmp9713 : tmp9747;
  assign tmp9749 = s2 ? 1 : tmp9710;
  assign tmp9748 = s3 ? tmp9749 : tmp9172;
  assign tmp9745 = s4 ? tmp9746 : tmp9748;
  assign tmp9737 = s5 ? tmp9738 : tmp9745;
  assign tmp9736 = s6 ? tmp9697 : tmp9737;
  assign tmp9718 = s7 ? tmp9719 : tmp9736;
  assign tmp9717 = s8 ? tmp9652 : tmp9718;
  assign tmp9590 = s9 ? tmp9591 : tmp9717;
  assign tmp9757 = s2 ? tmp9475 : tmp9172;
  assign tmp9756 = s3 ? tmp9757 : tmp9646;
  assign tmp9760 = s1 ? tmp9172 : tmp9610;
  assign tmp9759 = s2 ? 1 : tmp9760;
  assign tmp9758 = s3 ? tmp9759 : tmp9172;
  assign tmp9755 = s4 ? tmp9756 : tmp9758;
  assign tmp9754 = s5 ? tmp9633 : tmp9755;
  assign tmp9753 = s6 ? tmp9628 : tmp9754;
  assign tmp9752 = s7 ? tmp9593 : tmp9753;
  assign tmp9751 = s8 ? tmp9752 : tmp9593;
  assign tmp9766 = s3 ? tmp9504 : tmp9172;
  assign tmp9765 = s4 ? tmp9643 : tmp9766;
  assign tmp9764 = s5 ? tmp9633 : tmp9765;
  assign tmp9763 = s6 ? tmp9628 : tmp9764;
  assign tmp9771 = s2 ? 1 : tmp9657;
  assign tmp9770 = s3 ? tmp9771 : tmp9172;
  assign tmp9769 = s4 ? tmp9746 : tmp9770;
  assign tmp9768 = s5 ? tmp9738 : tmp9769;
  assign tmp9767 = s6 ? tmp9697 : tmp9768;
  assign tmp9762 = s7 ? tmp9763 : tmp9767;
  assign tmp9775 = s4 ? tmp9712 : tmp9770;
  assign tmp9774 = s5 ? tmp9702 : tmp9775;
  assign tmp9773 = s6 ? tmp9697 : tmp9774;
  assign tmp9778 = s4 ? tmp9756 : tmp9766;
  assign tmp9777 = s5 ? tmp9633 : tmp9778;
  assign tmp9776 = s6 ? tmp9628 : tmp9777;
  assign tmp9772 = s7 ? tmp9773 : tmp9776;
  assign tmp9761 = s8 ? tmp9762 : tmp9772;
  assign tmp9750 = s9 ? tmp9751 : tmp9761;
  assign tmp9589 = s10 ? tmp9590 : tmp9750;
  assign tmp9782 = s7 ? tmp9627 : tmp9736;
  assign tmp9783 = s7 ? tmp9696 : tmp9753;
  assign tmp9781 = s8 ? tmp9782 : tmp9783;
  assign tmp9780 = s9 ? tmp9751 : tmp9781;
  assign tmp9779 = s10 ? tmp9590 : tmp9780;
  assign tmp9588 = s11 ? tmp9589 : tmp9779;
  assign tmp9792 = ~(s2 ? tmp9172 : tmp9456);
  assign tmp9791 = s3 ? tmp9188 : tmp9792;
  assign tmp9794 = s2 ? tmp9456 : tmp9185;
  assign tmp9796 = s1 ? 1 : tmp9317;
  assign tmp9795 = ~(s2 ? tmp9796 : tmp9149);
  assign tmp9793 = ~(s3 ? tmp9794 : tmp9795);
  assign tmp9790 = s4 ? tmp9791 : tmp9793;
  assign tmp9801 = s1 ? tmp9186 : tmp9618;
  assign tmp9800 = s2 ? tmp9801 : tmp9511;
  assign tmp9799 = s3 ? tmp9800 : tmp9512;
  assign tmp9804 = ~(s1 ? 1 : tmp9470);
  assign tmp9803 = s2 ? tmp9481 : tmp9804;
  assign tmp9806 = s1 ? tmp9172 : tmp9618;
  assign tmp9805 = s2 ? tmp9806 : 1;
  assign tmp9802 = s3 ? tmp9803 : tmp9805;
  assign tmp9798 = s4 ? tmp9799 : tmp9802;
  assign tmp9808 = s3 ? tmp9757 : tmp9623;
  assign tmp9811 = s1 ? tmp9174 : tmp9172;
  assign tmp9810 = s2 ? tmp9172 : tmp9811;
  assign tmp9809 = s3 ? tmp9810 : tmp9482;
  assign tmp9807 = s4 ? tmp9808 : tmp9809;
  assign tmp9797 = ~(s5 ? tmp9798 : tmp9807);
  assign tmp9789 = s6 ? tmp9790 : tmp9797;
  assign tmp9816 = s1 ? 1 : 0;
  assign tmp9815 = ~(s2 ? tmp9816 : tmp9149);
  assign tmp9814 = ~(s3 ? tmp9794 : tmp9815);
  assign tmp9813 = s4 ? tmp9791 : tmp9814;
  assign tmp9820 = s2 ? tmp9456 : tmp9519;
  assign tmp9819 = s3 ? tmp9820 : tmp9424;
  assign tmp9822 = s2 ? tmp9481 : tmp9172;
  assign tmp9821 = s3 ? tmp9822 : tmp9416;
  assign tmp9818 = s4 ? tmp9819 : tmp9821;
  assign tmp9824 = s3 ? tmp9610 : tmp9172;
  assign tmp9823 = s4 ? tmp9756 : tmp9824;
  assign tmp9817 = ~(s5 ? tmp9818 : tmp9823);
  assign tmp9812 = s6 ? tmp9813 : tmp9817;
  assign tmp9788 = s7 ? tmp9789 : tmp9812;
  assign tmp9831 = s0 ? tmp9657 : 0;
  assign tmp9830 = s1 ? tmp9831 : tmp9657;
  assign tmp9832 = s1 ? tmp9831 : tmp9343;
  assign tmp9829 = s2 ? tmp9830 : tmp9832;
  assign tmp9833 = ~(s2 ? tmp9461 : tmp9659);
  assign tmp9828 = s3 ? tmp9829 : tmp9833;
  assign tmp9827 = s4 ? tmp9655 : tmp9828;
  assign tmp9839 = ~(s0 ? 1 : tmp9659);
  assign tmp9838 = s1 ? tmp9831 : tmp9839;
  assign tmp9841 = s0 ? 1 : tmp9659;
  assign tmp9842 = ~(s0 ? tmp9657 : 1);
  assign tmp9840 = ~(s1 ? tmp9841 : tmp9842);
  assign tmp9837 = s2 ? tmp9838 : tmp9840;
  assign tmp9836 = s3 ? tmp9837 : tmp9677;
  assign tmp9846 = ~(s0 ? 1 : tmp9151);
  assign tmp9845 = s1 ? tmp9670 : tmp9846;
  assign tmp9848 = ~(s0 ? tmp9657 : 0);
  assign tmp9847 = ~(s1 ? tmp9248 : tmp9848);
  assign tmp9844 = s2 ? tmp9845 : tmp9847;
  assign tmp9843 = s3 ? tmp9844 : tmp9684;
  assign tmp9835 = s4 ? tmp9836 : tmp9843;
  assign tmp9852 = s1 ? tmp9657 : tmp9691;
  assign tmp9851 = s2 ? tmp9689 : tmp9852;
  assign tmp9850 = s3 ? tmp9851 : tmp9623;
  assign tmp9849 = s4 ? tmp9850 : tmp9692;
  assign tmp9834 = s5 ? tmp9835 : tmp9849;
  assign tmp9826 = s6 ? tmp9827 : tmp9834;
  assign tmp9857 = s1 ? tmp9831 : tmp9257;
  assign tmp9856 = s2 ? tmp9830 : tmp9857;
  assign tmp9858 = ~(s2 ? tmp9491 : tmp9659);
  assign tmp9855 = s3 ? tmp9856 : tmp9858;
  assign tmp9854 = s4 ? tmp9655 : tmp9855;
  assign tmp9862 = s2 ? tmp9830 : tmp9705;
  assign tmp9861 = s3 ? tmp9862 : tmp9706;
  assign tmp9864 = s2 ? tmp9845 : tmp9657;
  assign tmp9863 = s3 ? tmp9864 : tmp9709;
  assign tmp9860 = s4 ? tmp9861 : tmp9863;
  assign tmp9859 = s5 ? tmp9860 : tmp9711;
  assign tmp9853 = s6 ? tmp9854 : tmp9859;
  assign tmp9825 = ~(s7 ? tmp9826 : tmp9853);
  assign tmp9787 = s8 ? tmp9788 : tmp9825;
  assign tmp9866 = s7 ? tmp9826 : tmp9853;
  assign tmp9872 = s2 ? tmp9801 : tmp9187;
  assign tmp9871 = s3 ? tmp9872 : tmp9424;
  assign tmp9870 = s4 ? tmp9871 : tmp9802;
  assign tmp9869 = ~(s5 ? tmp9870 : tmp9807);
  assign tmp9868 = s6 ? tmp9790 : tmp9869;
  assign tmp9877 = s2 ? tmp9456 : tmp9172;
  assign tmp9876 = s3 ? tmp9877 : tmp9424;
  assign tmp9875 = s4 ? tmp9876 : tmp9821;
  assign tmp9879 = s3 ? tmp9757 : tmp9747;
  assign tmp9878 = s4 ? tmp9879 : tmp9172;
  assign tmp9874 = ~(s5 ? tmp9875 : tmp9878);
  assign tmp9873 = s6 ? tmp9813 : tmp9874;
  assign tmp9867 = ~(s7 ? tmp9868 : tmp9873);
  assign tmp9865 = ~(s8 ? tmp9866 : tmp9867);
  assign tmp9786 = s9 ? tmp9787 : tmp9865;
  assign tmp9884 = ~(s5 ? tmp9875 : tmp9823);
  assign tmp9883 = s6 ? tmp9813 : tmp9884;
  assign tmp9882 = s7 ? tmp9868 : tmp9883;
  assign tmp9881 = s8 ? tmp9882 : tmp9868;
  assign tmp9887 = ~(s5 ? tmp9818 : tmp9778);
  assign tmp9886 = s6 ? tmp9813 : tmp9887;
  assign tmp9890 = s5 ? tmp9860 : tmp9775;
  assign tmp9889 = s6 ? tmp9854 : tmp9890;
  assign tmp9892 = ~(s5 ? tmp9875 : tmp9778);
  assign tmp9891 = ~(s6 ? tmp9813 : tmp9892);
  assign tmp9888 = ~(s7 ? tmp9889 : tmp9891);
  assign tmp9885 = s8 ? tmp9886 : tmp9888;
  assign tmp9880 = s9 ? tmp9881 : tmp9885;
  assign tmp9785 = s10 ? tmp9786 : tmp9880;
  assign tmp9897 = ~(s6 ? tmp9813 : tmp9884);
  assign tmp9896 = ~(s7 ? tmp9853 : tmp9897);
  assign tmp9895 = s8 ? tmp9812 : tmp9896;
  assign tmp9894 = s9 ? tmp9881 : tmp9895;
  assign tmp9893 = s10 ? tmp9786 : tmp9894;
  assign tmp9784 = ~(s11 ? tmp9785 : tmp9893);
  assign tmp9587 = s12 ? tmp9588 : tmp9784;
  assign tmp9399 = ~(s13 ? tmp9400 : tmp9587);
  assign tmp9137 = s14 ? tmp9138 : tmp9399;
  assign tmp9908 = s1 ? 1 : tmp9659;
  assign tmp9907 = ~(s2 ? tmp9841 : tmp9908);
  assign tmp9906 = s3 ? tmp9181 : tmp9907;
  assign tmp9911 = ~(s1 ? tmp9186 : 0);
  assign tmp9910 = s2 ? tmp9908 : tmp9911;
  assign tmp9913 = s1 ? 1 : tmp9841;
  assign tmp9912 = s2 ? tmp9913 : tmp9659;
  assign tmp9909 = ~(s3 ? tmp9910 : tmp9912);
  assign tmp9905 = s4 ? tmp9906 : tmp9909;
  assign tmp9918 = s1 ? 1 : tmp9848;
  assign tmp9917 = s2 ? 1 : tmp9918;
  assign tmp9916 = s3 ? tmp9917 : tmp9912;
  assign tmp9921 = s1 ? tmp9657 : 0;
  assign tmp9920 = s2 ? tmp9921 : 0;
  assign tmp9923 = s1 ? tmp9188 : tmp9841;
  assign tmp9922 = ~(s2 ? tmp9923 : tmp9659);
  assign tmp9919 = ~(s3 ? tmp9920 : tmp9922);
  assign tmp9915 = s4 ? tmp9916 : tmp9919;
  assign tmp9927 = s1 ? tmp9657 : tmp9831;
  assign tmp9926 = s2 ? tmp9927 : 0;
  assign tmp9929 = s1 ? 1 : tmp9248;
  assign tmp9930 = s1 ? tmp9224 : tmp9470;
  assign tmp9928 = ~(s2 ? tmp9929 : tmp9930);
  assign tmp9925 = s3 ? tmp9926 : tmp9928;
  assign tmp9933 = ~(s1 ? tmp9831 : 0);
  assign tmp9932 = s2 ? tmp9913 : tmp9933;
  assign tmp9935 = s1 ? tmp9151 : tmp9224;
  assign tmp9934 = s2 ? tmp9935 : tmp9911;
  assign tmp9931 = ~(s3 ? tmp9932 : tmp9934);
  assign tmp9924 = ~(s4 ? tmp9925 : tmp9931);
  assign tmp9914 = ~(s5 ? tmp9915 : tmp9924);
  assign tmp9904 = s6 ? tmp9905 : tmp9914;
  assign tmp9939 = s2 ? tmp9908 : tmp9659;
  assign tmp9938 = ~(s3 ? tmp9910 : tmp9939);
  assign tmp9937 = s4 ? tmp9906 : tmp9938;
  assign tmp9942 = s3 ? tmp9917 : tmp9939;
  assign tmp9945 = s1 ? tmp9188 : tmp9659;
  assign tmp9944 = ~(s2 ? tmp9945 : tmp9659);
  assign tmp9943 = ~(s3 ? tmp9920 : tmp9944);
  assign tmp9941 = s4 ? tmp9942 : tmp9943;
  assign tmp9949 = s1 ? 1 : tmp9151;
  assign tmp9950 = ~(s1 ? tmp9172 : 0);
  assign tmp9948 = ~(s2 ? tmp9949 : tmp9950);
  assign tmp9947 = s3 ? tmp9926 : tmp9948;
  assign tmp9952 = s2 ? tmp9908 : tmp9848;
  assign tmp9951 = ~(s3 ? tmp9952 : tmp9381);
  assign tmp9946 = ~(s4 ? tmp9947 : tmp9951);
  assign tmp9940 = ~(s5 ? tmp9941 : tmp9946);
  assign tmp9936 = s6 ? tmp9937 : tmp9940;
  assign tmp9903 = s7 ? tmp9904 : tmp9936;
  assign tmp9954 = s8 ? tmp9903 : tmp9904;
  assign tmp9959 = s2 ? tmp9908 : 1;
  assign tmp9958 = ~(s3 ? tmp9959 : tmp9381);
  assign tmp9957 = ~(s4 ? tmp9947 : tmp9958);
  assign tmp9956 = ~(s5 ? tmp9941 : tmp9957);
  assign tmp9955 = s6 ? tmp9937 : tmp9956;
  assign tmp9953 = s9 ? tmp9954 : tmp9955;
  assign tmp9902 = s10 ? tmp9903 : tmp9953;
  assign tmp9961 = s9 ? tmp9954 : tmp9936;
  assign tmp9960 = s10 ? tmp9903 : tmp9961;
  assign tmp9901 = s11 ? tmp9902 : tmp9960;
  assign tmp9969 = l1 ? 1 : tmp9172;
  assign tmp9968 = s0 ? tmp9151 : tmp9969;
  assign tmp9971 = s0 ? tmp9969 : tmp9151;
  assign tmp9970 = s1 ? tmp9151 : tmp9971;
  assign tmp9967 = s2 ? tmp9968 : tmp9970;
  assign tmp9966 = s3 ? tmp9491 : tmp9967;
  assign tmp9974 = s1 ? tmp9151 : tmp9968;
  assign tmp9973 = s2 ? tmp9974 : tmp9151;
  assign tmp9975 = s2 ? tmp9974 : tmp9969;
  assign tmp9972 = s3 ? tmp9973 : tmp9975;
  assign tmp9965 = s4 ? tmp9966 : tmp9972;
  assign tmp9981 = ~(s0 ? tmp9969 : 1);
  assign tmp9980 = s1 ? 1 : tmp9981;
  assign tmp9979 = s2 ? 1 : tmp9980;
  assign tmp9984 = s0 ? 1 : tmp9969;
  assign tmp9983 = s1 ? tmp9151 : tmp9984;
  assign tmp9982 = ~(s2 ? tmp9983 : tmp9969);
  assign tmp9978 = s3 ? tmp9979 : tmp9982;
  assign tmp9987 = s1 ? tmp9971 : tmp9151;
  assign tmp9986 = s2 ? tmp9987 : tmp9151;
  assign tmp9985 = ~(s3 ? tmp9986 : tmp9975);
  assign tmp9977 = s4 ? tmp9978 : tmp9985;
  assign tmp9991 = s1 ? tmp9969 : tmp9248;
  assign tmp9990 = s2 ? tmp9991 : tmp9151;
  assign tmp9993 = s1 ? 1 : tmp9188;
  assign tmp9995 = s0 ? tmp9172 : tmp9151;
  assign tmp9994 = ~(s1 ? tmp9995 : tmp9151);
  assign tmp9992 = ~(s2 ? tmp9993 : tmp9994);
  assign tmp9989 = s3 ? tmp9990 : tmp9992;
  assign tmp10000 = ~(l1 ? 1 : tmp9172);
  assign tmp9999 = s0 ? 1 : tmp10000;
  assign tmp9998 = s1 ? 1 : tmp9999;
  assign tmp9997 = s2 ? tmp9998 : tmp9545;
  assign tmp10003 = ~(s0 ? tmp9172 : tmp9151);
  assign tmp10002 = s1 ? tmp9188 : tmp10003;
  assign tmp10004 = ~(s1 ? tmp9254 : 0);
  assign tmp10001 = s2 ? tmp10002 : tmp10004;
  assign tmp9996 = ~(s3 ? tmp9997 : tmp10001);
  assign tmp9988 = ~(s4 ? tmp9989 : tmp9996);
  assign tmp9976 = ~(s5 ? tmp9977 : tmp9988);
  assign tmp9964 = s6 ? tmp9965 : tmp9976;
  assign tmp10009 = s1 ? tmp9151 : tmp9969;
  assign tmp10008 = s2 ? tmp10009 : tmp9969;
  assign tmp10007 = s3 ? tmp9973 : tmp10008;
  assign tmp10006 = s4 ? tmp9966 : tmp10007;
  assign tmp10013 = ~(s2 ? tmp10009 : tmp9969);
  assign tmp10012 = s3 ? tmp9979 : tmp10013;
  assign tmp10014 = ~(s3 ? tmp9986 : tmp10008);
  assign tmp10011 = s4 ? tmp10012 : tmp10014;
  assign tmp10018 = s1 ? tmp9969 : tmp9151;
  assign tmp10017 = s2 ? tmp10018 : tmp9151;
  assign tmp10020 = s1 ? 1 : tmp9149;
  assign tmp10019 = ~(s2 ? tmp10020 : tmp9257);
  assign tmp10016 = s3 ? tmp10017 : tmp10019;
  assign tmp10023 = s1 ? 1 : tmp10000;
  assign tmp10022 = s2 ? tmp10023 : 1;
  assign tmp10024 = ~(s1 ? tmp9172 : tmp9151);
  assign tmp10021 = ~(s3 ? tmp10022 : tmp10024);
  assign tmp10015 = ~(s4 ? tmp10016 : tmp10021);
  assign tmp10010 = ~(s5 ? tmp10011 : tmp10015);
  assign tmp10005 = s6 ? tmp10006 : tmp10010;
  assign tmp9963 = s7 ? tmp9964 : tmp10005;
  assign tmp10026 = s8 ? tmp9963 : tmp9964;
  assign tmp10025 = s9 ? tmp10026 : tmp10005;
  assign tmp9962 = s10 ? tmp9963 : tmp10025;
  assign tmp9900 = s12 ? tmp9901 : tmp9962;
  assign tmp10036 = s1 ? tmp9172 : tmp9320;
  assign tmp10038 = s1 ? tmp9174 : tmp9454;
  assign tmp10039 = ~(s1 ? tmp9254 : tmp9149);
  assign tmp10037 = s2 ? tmp10038 : tmp10039;
  assign tmp10035 = s3 ? tmp10036 : tmp10037;
  assign tmp10041 = s2 ? tmp9432 : tmp9475;
  assign tmp10042 = s2 ? tmp9483 : tmp9172;
  assign tmp10040 = s3 ? tmp10041 : tmp10042;
  assign tmp10034 = s4 ? tmp10035 : tmp10040;
  assign tmp10046 = s2 ? tmp9355 : tmp9201;
  assign tmp10048 = s1 ? tmp9256 : tmp9174;
  assign tmp10047 = ~(s2 ? tmp10048 : tmp9641);
  assign tmp10045 = s3 ? tmp10046 : tmp10047;
  assign tmp10051 = s1 ? 1 : tmp9433;
  assign tmp10050 = s2 ? tmp9383 : tmp10051;
  assign tmp10053 = s1 ? tmp9151 : tmp9995;
  assign tmp10052 = s2 ? tmp9172 : tmp10053;
  assign tmp10049 = ~(s3 ? tmp10050 : tmp10052);
  assign tmp10044 = s4 ? tmp10045 : tmp10049;
  assign tmp10057 = s1 ? tmp9172 : tmp9599;
  assign tmp10056 = s2 ? tmp10057 : tmp10004;
  assign tmp10058 = ~(s2 ? 1 : tmp9191);
  assign tmp10055 = s3 ? tmp10056 : tmp10058;
  assign tmp10062 = s0 ? tmp9172 : tmp9320;
  assign tmp10061 = s1 ? tmp10062 : 1;
  assign tmp10060 = s2 ? tmp9801 : tmp10061;
  assign tmp10064 = s1 ? tmp9159 : tmp9188;
  assign tmp10063 = ~(s2 ? tmp10064 : tmp9950);
  assign tmp10059 = s3 ? tmp10060 : tmp10063;
  assign tmp10054 = ~(s4 ? tmp10055 : tmp10059);
  assign tmp10043 = ~(s5 ? tmp10044 : tmp10054);
  assign tmp10033 = s6 ? tmp10034 : tmp10043;
  assign tmp10068 = s2 ? tmp9425 : tmp9172;
  assign tmp10067 = s3 ? tmp10041 : tmp10068;
  assign tmp10066 = s4 ? tmp10035 : tmp10067;
  assign tmp10073 = ~(s1 ? tmp9609 : tmp9172);
  assign tmp10072 = s2 ? tmp9381 : tmp10073;
  assign tmp10071 = s3 ? tmp10046 : tmp10072;
  assign tmp10075 = s2 ? tmp9383 : tmp9172;
  assign tmp10077 = s1 ? tmp9151 : tmp9172;
  assign tmp10076 = s2 ? tmp9172 : tmp10077;
  assign tmp10074 = ~(s3 ? tmp10075 : tmp10076);
  assign tmp10070 = s4 ? tmp10071 : tmp10074;
  assign tmp10081 = s1 ? tmp9172 : tmp9257;
  assign tmp10080 = s2 ? tmp10081 : 1;
  assign tmp10082 = ~(s2 ? 1 : tmp9149);
  assign tmp10079 = s3 ? tmp10080 : tmp10082;
  assign tmp10084 = s2 ? tmp10020 : tmp9148;
  assign tmp10085 = s2 ? tmp10020 : tmp9149;
  assign tmp10083 = ~(s3 ? tmp10084 : tmp10085);
  assign tmp10078 = ~(s4 ? tmp10079 : tmp10083);
  assign tmp10069 = ~(s5 ? tmp10070 : tmp10078);
  assign tmp10065 = s6 ? tmp10066 : tmp10069;
  assign tmp10032 = s7 ? tmp10033 : tmp10065;
  assign tmp10090 = s2 ? tmp9172 : tmp9475;
  assign tmp10089 = s3 ? tmp10090 : tmp10042;
  assign tmp10088 = s4 ? tmp10035 : tmp10089;
  assign tmp10094 = s2 ? tmp9383 : tmp9425;
  assign tmp10093 = ~(s3 ? tmp10094 : tmp10052);
  assign tmp10092 = s4 ? tmp10045 : tmp10093;
  assign tmp10091 = ~(s5 ? tmp10092 : tmp10054);
  assign tmp10087 = s6 ? tmp10088 : tmp10091;
  assign tmp10097 = s3 ? tmp10090 : tmp10068;
  assign tmp10096 = s4 ? tmp10035 : tmp10097;
  assign tmp10095 = s6 ? tmp10096 : tmp10069;
  assign tmp10086 = s7 ? tmp10087 : tmp10095;
  assign tmp10031 = s8 ? tmp10032 : tmp10086;
  assign tmp10104 = s2 ? tmp10057 : tmp9257;
  assign tmp10103 = s3 ? tmp10104 : tmp10058;
  assign tmp10106 = s2 ? tmp9801 : tmp10062;
  assign tmp10105 = s3 ? tmp10106 : tmp10063;
  assign tmp10102 = ~(s4 ? tmp10103 : tmp10105);
  assign tmp10101 = ~(s5 ? tmp10092 : tmp10102);
  assign tmp10100 = s6 ? tmp10088 : tmp10101;
  assign tmp10110 = s3 ? tmp10081 : tmp10082;
  assign tmp10109 = ~(s4 ? tmp10110 : tmp10083);
  assign tmp10108 = ~(s5 ? tmp10070 : tmp10109);
  assign tmp10107 = s6 ? tmp10096 : tmp10108;
  assign tmp10099 = s7 ? tmp10100 : tmp10107;
  assign tmp10098 = s8 ? tmp10086 : tmp10099;
  assign tmp10030 = s9 ? tmp10031 : tmp10098;
  assign tmp10112 = s8 ? tmp10099 : tmp10100;
  assign tmp10118 = ~(s3 ? tmp10084 : tmp10020);
  assign tmp10117 = ~(s4 ? tmp10079 : tmp10118);
  assign tmp10116 = ~(s5 ? tmp10070 : tmp10117);
  assign tmp10115 = s6 ? tmp10066 : tmp10116;
  assign tmp10121 = ~(s4 ? tmp10110 : tmp10118);
  assign tmp10120 = ~(s5 ? tmp10070 : tmp10121);
  assign tmp10119 = s6 ? tmp10096 : tmp10120;
  assign tmp10114 = s7 ? tmp10115 : tmp10119;
  assign tmp10123 = s6 ? tmp10096 : tmp10116;
  assign tmp10122 = s7 ? tmp10123 : tmp10119;
  assign tmp10113 = s8 ? tmp10114 : tmp10122;
  assign tmp10111 = s9 ? tmp10112 : tmp10113;
  assign tmp10029 = s10 ? tmp10030 : tmp10111;
  assign tmp10127 = s7 ? tmp10065 : tmp10107;
  assign tmp10128 = s7 ? tmp10095 : tmp10107;
  assign tmp10126 = s8 ? tmp10127 : tmp10128;
  assign tmp10125 = s9 ? tmp10112 : tmp10126;
  assign tmp10124 = s10 ? tmp10030 : tmp10125;
  assign tmp10028 = s11 ? tmp10029 : tmp10124;
  assign tmp10135 = s2 ? tmp9164 : tmp9225;
  assign tmp10134 = s3 ? 1 : tmp10135;
  assign tmp10138 = s1 ? 1 : tmp9164;
  assign tmp10137 = s2 ? tmp10138 : 1;
  assign tmp10139 = s2 ? tmp10138 : tmp9148;
  assign tmp10136 = s3 ? tmp10137 : tmp10139;
  assign tmp10133 = s4 ? tmp10134 : tmp10136;
  assign tmp10143 = s2 ? 1 : tmp9225;
  assign tmp10142 = s3 ? tmp10143 : tmp10139;
  assign tmp10146 = s1 ? tmp9158 : 1;
  assign tmp10145 = s2 ? tmp10146 : 1;
  assign tmp10144 = s3 ? tmp10145 : tmp10139;
  assign tmp10141 = s4 ? tmp10142 : tmp10144;
  assign tmp10150 = s1 ? tmp9148 : tmp9159;
  assign tmp10149 = s2 ? tmp10150 : 1;
  assign tmp10151 = s2 ? tmp10138 : tmp10146;
  assign tmp10148 = s3 ? tmp10149 : tmp10151;
  assign tmp10153 = s2 ? tmp10138 : tmp9267;
  assign tmp10155 = s1 ? tmp9164 : tmp9158;
  assign tmp10154 = s2 ? tmp10155 : 1;
  assign tmp10152 = s3 ? tmp10153 : tmp10154;
  assign tmp10147 = s4 ? tmp10148 : tmp10152;
  assign tmp10140 = s5 ? tmp10141 : tmp10147;
  assign tmp10132 = s6 ? tmp10133 : tmp10140;
  assign tmp10160 = s1 ? 1 : tmp9148;
  assign tmp10159 = s2 ? tmp10160 : tmp9148;
  assign tmp10158 = s3 ? tmp10137 : tmp10159;
  assign tmp10157 = s4 ? tmp10134 : tmp10158;
  assign tmp10163 = s3 ? tmp10143 : tmp10159;
  assign tmp10164 = s3 ? tmp10145 : tmp10159;
  assign tmp10162 = s4 ? tmp10163 : tmp10164;
  assign tmp10168 = s1 ? tmp9148 : 1;
  assign tmp10167 = s2 ? tmp10168 : 1;
  assign tmp10169 = s2 ? tmp10160 : tmp10146;
  assign tmp10166 = s3 ? tmp10167 : tmp10169;
  assign tmp10171 = s2 ? tmp10160 : 1;
  assign tmp10172 = s1 ? tmp9148 : tmp9158;
  assign tmp10170 = s3 ? tmp10171 : tmp10172;
  assign tmp10165 = s4 ? tmp10166 : tmp10170;
  assign tmp10161 = s5 ? tmp10162 : tmp10165;
  assign tmp10156 = s6 ? tmp10157 : tmp10161;
  assign tmp10131 = s7 ? tmp10132 : tmp10156;
  assign tmp10174 = s8 ? tmp10131 : tmp10132;
  assign tmp10178 = s3 ? tmp10171 : tmp10168;
  assign tmp10177 = s4 ? tmp10166 : tmp10178;
  assign tmp10176 = s5 ? tmp10162 : tmp10177;
  assign tmp10175 = s6 ? tmp10157 : tmp10176;
  assign tmp10173 = s9 ? tmp10174 : tmp10175;
  assign tmp10130 = s10 ? tmp10131 : tmp10173;
  assign tmp10180 = s9 ? tmp10174 : tmp10156;
  assign tmp10179 = s10 ? tmp10131 : tmp10180;
  assign tmp10129 = ~(s11 ? tmp10130 : tmp10179);
  assign tmp10027 = s12 ? tmp10028 : tmp10129;
  assign tmp9899 = s13 ? tmp9900 : tmp10027;
  assign tmp10192 = s1 ? tmp9622 : tmp9172;
  assign tmp10191 = s2 ? tmp10192 : tmp9456;
  assign tmp10190 = s3 ? tmp9453 : tmp10191;
  assign tmp10195 = s1 ? tmp9151 : tmp9188;
  assign tmp10194 = ~(s2 ? tmp10195 : tmp9149);
  assign tmp10193 = s3 ? tmp9458 : tmp10194;
  assign tmp10189 = s4 ? tmp10190 : tmp10193;
  assign tmp10200 = ~(s1 ? tmp9186 : tmp9172);
  assign tmp10199 = ~(s2 ? tmp9188 : tmp10200);
  assign tmp10198 = s3 ? tmp9800 : tmp10199;
  assign tmp10203 = s1 ? tmp9172 : tmp9846;
  assign tmp10204 = ~(s1 ? tmp9248 : tmp9470);
  assign tmp10202 = s2 ? tmp10203 : tmp10204;
  assign tmp10205 = s2 ? tmp9453 : tmp9172;
  assign tmp10201 = s3 ? tmp10202 : tmp10205;
  assign tmp10197 = s4 ? tmp10198 : tmp10201;
  assign tmp10208 = s2 ? tmp9383 : tmp9811;
  assign tmp10207 = s3 ? tmp10208 : tmp9184;
  assign tmp10212 = s0 ? tmp9151 : tmp9172;
  assign tmp10211 = s1 ? tmp9995 : tmp10212;
  assign tmp10210 = s2 ? tmp10211 : tmp9172;
  assign tmp10214 = s1 ? tmp9248 : tmp9618;
  assign tmp10215 = s1 ? tmp9172 : tmp9531;
  assign tmp10213 = s2 ? tmp10214 : tmp10215;
  assign tmp10209 = s3 ? tmp10210 : tmp10213;
  assign tmp10206 = s4 ? tmp10207 : tmp10209;
  assign tmp10196 = s5 ? tmp10197 : tmp10206;
  assign tmp10188 = s6 ? tmp10189 : tmp10196;
  assign tmp10219 = ~(s2 ? tmp9148 : tmp9149);
  assign tmp10218 = s3 ? tmp9488 : tmp10219;
  assign tmp10217 = s4 ? tmp10190 : tmp10218;
  assign tmp10222 = s3 ? tmp9820 : tmp9455;
  assign tmp10224 = s2 ? tmp10203 : tmp9498;
  assign tmp10223 = s3 ? tmp10224 : tmp10205;
  assign tmp10221 = s4 ? tmp10222 : tmp10223;
  assign tmp10229 = s0 ? tmp9610 : 0;
  assign tmp10228 = s1 ? tmp10229 : 0;
  assign tmp10227 = s2 ? tmp10228 : tmp9172;
  assign tmp10226 = s3 ? tmp10075 : tmp10227;
  assign tmp10232 = s1 ? tmp9995 : tmp9172;
  assign tmp10231 = s2 ? tmp10232 : tmp9760;
  assign tmp10233 = s2 ? tmp10077 : tmp9172;
  assign tmp10230 = s3 ? tmp10231 : tmp10233;
  assign tmp10225 = s4 ? tmp10226 : tmp10230;
  assign tmp10220 = s5 ? tmp10221 : tmp10225;
  assign tmp10216 = s6 ? tmp10217 : tmp10220;
  assign tmp10187 = s7 ? tmp10188 : tmp10216;
  assign tmp10239 = s1 ? tmp9662 : tmp9172;
  assign tmp10238 = s2 ? tmp9172 : tmp10239;
  assign tmp10237 = s3 ? tmp9453 : tmp10238;
  assign tmp10236 = s4 ? tmp10237 : tmp10193;
  assign tmp10244 = s1 ? tmp9186 : tmp9839;
  assign tmp10245 = ~(s1 ? tmp9188 : tmp9171);
  assign tmp10243 = s2 ? tmp10244 : tmp10245;
  assign tmp10248 = s0 ? tmp9969 : 0;
  assign tmp10247 = s1 ? tmp10248 : tmp9172;
  assign tmp10246 = s2 ? tmp9174 : tmp10247;
  assign tmp10242 = s3 ? tmp10243 : tmp10246;
  assign tmp10241 = s4 ? tmp10242 : tmp10201;
  assign tmp10251 = s2 ? tmp9383 : tmp9690;
  assign tmp10250 = s3 ? tmp10251 : tmp9184;
  assign tmp10254 = s1 ? tmp9995 : tmp9968;
  assign tmp10255 = s1 ? tmp9172 : tmp9695;
  assign tmp10253 = s2 ? tmp10254 : tmp10255;
  assign tmp10252 = s3 ? tmp10253 : tmp10213;
  assign tmp10249 = s4 ? tmp10250 : tmp10252;
  assign tmp10240 = s5 ? tmp10241 : tmp10249;
  assign tmp10235 = s6 ? tmp10236 : tmp10240;
  assign tmp10259 = ~(s2 ? tmp9381 : tmp9149);
  assign tmp10258 = s3 ? tmp9488 : tmp10259;
  assign tmp10257 = s4 ? tmp10237 : tmp10258;
  assign tmp10264 = s1 ? tmp9186 : tmp9657;
  assign tmp10263 = s2 ? tmp10264 : tmp9636;
  assign tmp10265 = s2 ? tmp9172 : tmp10247;
  assign tmp10262 = s3 ? tmp10263 : tmp10265;
  assign tmp10267 = s2 ? tmp10203 : tmp9172;
  assign tmp10266 = s3 ? tmp10267 : tmp9172;
  assign tmp10261 = s4 ? tmp10262 : tmp10266;
  assign tmp10270 = s2 ? tmp9383 : tmp9710;
  assign tmp10269 = s3 ? tmp10270 : tmp10227;
  assign tmp10273 = s1 ? tmp9995 : tmp9969;
  assign tmp10272 = s2 ? tmp10273 : tmp9760;
  assign tmp10271 = s3 ? tmp10272 : tmp10233;
  assign tmp10268 = s4 ? tmp10269 : tmp10271;
  assign tmp10260 = s5 ? tmp10261 : tmp10268;
  assign tmp10256 = s6 ? tmp10257 : tmp10260;
  assign tmp10234 = s7 ? tmp10235 : tmp10256;
  assign tmp10186 = s8 ? tmp10187 : tmp10234;
  assign tmp10277 = s4 ? tmp9452 : tmp10193;
  assign tmp10280 = s3 ? tmp9872 : tmp9455;
  assign tmp10279 = s4 ? tmp10280 : tmp10201;
  assign tmp10278 = s5 ? tmp10279 : tmp10206;
  assign tmp10276 = s6 ? tmp10277 : tmp10278;
  assign tmp10282 = s4 ? tmp9452 : tmp10218;
  assign tmp10285 = s3 ? tmp9877 : tmp9455;
  assign tmp10284 = s4 ? tmp10285 : tmp10266;
  assign tmp10287 = s3 ? tmp10075 : tmp9495;
  assign tmp10289 = s2 ? tmp10232 : tmp9172;
  assign tmp10288 = s3 ? tmp10289 : tmp10233;
  assign tmp10286 = s4 ? tmp10287 : tmp10288;
  assign tmp10283 = s5 ? tmp10284 : tmp10286;
  assign tmp10281 = s6 ? tmp10282 : tmp10283;
  assign tmp10275 = s7 ? tmp10276 : tmp10281;
  assign tmp10274 = s8 ? tmp10234 : tmp10275;
  assign tmp10185 = s9 ? tmp10186 : tmp10274;
  assign tmp10293 = s6 ? tmp10189 : tmp10278;
  assign tmp10295 = s5 ? tmp10284 : tmp10225;
  assign tmp10294 = s6 ? tmp10217 : tmp10295;
  assign tmp10292 = s7 ? tmp10293 : tmp10294;
  assign tmp10291 = s8 ? tmp10292 : tmp10293;
  assign tmp10301 = s3 ? tmp10224 : tmp9172;
  assign tmp10300 = s4 ? tmp10222 : tmp10301;
  assign tmp10303 = s3 ? tmp10289 : tmp10077;
  assign tmp10302 = s4 ? tmp10226 : tmp10303;
  assign tmp10299 = s5 ? tmp10300 : tmp10302;
  assign tmp10298 = s6 ? tmp10217 : tmp10299;
  assign tmp10306 = s4 ? tmp10287 : tmp10303;
  assign tmp10305 = s5 ? tmp10284 : tmp10306;
  assign tmp10304 = s6 ? tmp10282 : tmp10305;
  assign tmp10297 = s7 ? tmp10298 : tmp10304;
  assign tmp10312 = s2 ? tmp10273 : tmp9172;
  assign tmp10311 = s3 ? tmp10312 : tmp10077;
  assign tmp10310 = s4 ? tmp10269 : tmp10311;
  assign tmp10309 = s5 ? tmp10261 : tmp10310;
  assign tmp10308 = s6 ? tmp10257 : tmp10309;
  assign tmp10314 = s5 ? tmp10284 : tmp10302;
  assign tmp10313 = s6 ? tmp10217 : tmp10314;
  assign tmp10307 = s7 ? tmp10308 : tmp10313;
  assign tmp10296 = s8 ? tmp10297 : tmp10307;
  assign tmp10290 = s9 ? tmp10291 : tmp10296;
  assign tmp10184 = s10 ? tmp10185 : tmp10290;
  assign tmp10318 = s7 ? tmp10216 : tmp10281;
  assign tmp10319 = s7 ? tmp10256 : tmp10294;
  assign tmp10317 = s8 ? tmp10318 : tmp10319;
  assign tmp10316 = s9 ? tmp10291 : tmp10317;
  assign tmp10315 = s10 ? tmp10185 : tmp10316;
  assign tmp10183 = s11 ? tmp10184 : tmp10315;
  assign tmp10328 = s1 ? tmp9657 : tmp9670;
  assign tmp10330 = s1 ? tmp9670 : tmp9657;
  assign tmp10329 = s2 ? tmp10330 : tmp9661;
  assign tmp10327 = s3 ? tmp10328 : tmp10329;
  assign tmp10332 = s2 ? tmp9678 : tmp9689;
  assign tmp10333 = s2 ? tmp9552 : tmp9657;
  assign tmp10331 = s3 ? tmp10332 : tmp10333;
  assign tmp10326 = s4 ? tmp10327 : tmp10331;
  assign tmp10337 = s2 ? tmp9689 : tmp9676;
  assign tmp10338 = s2 ? tmp9670 : tmp9830;
  assign tmp10336 = s3 ? tmp10337 : tmp10338;
  assign tmp10342 = s0 ? tmp9151 : tmp9659;
  assign tmp10341 = s1 ? tmp10342 : 0;
  assign tmp10340 = s2 ? tmp10341 : 0;
  assign tmp10343 = ~(s2 ? tmp10328 : tmp9258);
  assign tmp10339 = ~(s3 ? tmp10340 : tmp10343);
  assign tmp10335 = s4 ? tmp10336 : tmp10339;
  assign tmp10346 = s2 ? tmp9838 : tmp9689;
  assign tmp10348 = ~(s1 ? tmp9151 : tmp9254);
  assign tmp10347 = s2 ? tmp9476 : tmp10348;
  assign tmp10345 = s3 ? tmp10346 : tmp10347;
  assign tmp10351 = s1 ? tmp9174 : tmp9657;
  assign tmp10352 = ~(s1 ? tmp9841 : 0);
  assign tmp10350 = s2 ? tmp10351 : tmp10352;
  assign tmp10354 = s1 ? tmp9657 : tmp9839;
  assign tmp10355 = ~(s1 ? tmp9254 : tmp9188);
  assign tmp10353 = s2 ? tmp10354 : tmp10355;
  assign tmp10349 = s3 ? tmp10350 : tmp10353;
  assign tmp10344 = s4 ? tmp10345 : tmp10349;
  assign tmp10334 = s5 ? tmp10335 : tmp10344;
  assign tmp10325 = s6 ? tmp10326 : tmp10334;
  assign tmp10359 = s2 ? tmp9566 : tmp9657;
  assign tmp10358 = s3 ? tmp10332 : tmp10359;
  assign tmp10357 = s4 ? tmp10327 : tmp10358;
  assign tmp10363 = s2 ? tmp9689 : tmp9705;
  assign tmp10364 = s2 ? tmp9657 : tmp9830;
  assign tmp10362 = s3 ? tmp10363 : tmp10364;
  assign tmp10367 = ~(s1 ? 1 : tmp9151);
  assign tmp10366 = ~(s2 ? tmp9657 : tmp10367);
  assign tmp10365 = ~(s3 ? tmp10340 : tmp10366);
  assign tmp10361 = s4 ? tmp10362 : tmp10365;
  assign tmp10370 = s2 ? tmp9830 : tmp9689;
  assign tmp10371 = ~(s2 ? 1 : tmp9491);
  assign tmp10369 = s3 ? tmp10370 : tmp10371;
  assign tmp10368 = s4 ? tmp10369 : tmp9657;
  assign tmp10360 = s5 ? tmp10361 : tmp10368;
  assign tmp10356 = s6 ? tmp10357 : tmp10360;
  assign tmp10324 = s7 ? tmp10325 : tmp10356;
  assign tmp10378 = s1 ? tmp9174 : tmp9691;
  assign tmp10377 = s2 ? tmp10378 : tmp10352;
  assign tmp10380 = s1 ? tmp9695 : tmp9839;
  assign tmp10379 = s2 ? tmp10380 : tmp10355;
  assign tmp10376 = s3 ? tmp10377 : tmp10379;
  assign tmp10375 = s4 ? tmp10345 : tmp10376;
  assign tmp10374 = s5 ? tmp10335 : tmp10375;
  assign tmp10373 = s6 ? tmp10326 : tmp10374;
  assign tmp10385 = s2 ? tmp9830 : 1;
  assign tmp10384 = s3 ? tmp10385 : tmp10371;
  assign tmp10388 = s1 ? tmp9172 : tmp9657;
  assign tmp10387 = s2 ? tmp10388 : tmp9657;
  assign tmp10386 = s3 ? tmp10387 : tmp10388;
  assign tmp10383 = s4 ? tmp10384 : tmp10386;
  assign tmp10382 = s5 ? tmp10361 : tmp10383;
  assign tmp10381 = s6 ? tmp10357 : tmp10382;
  assign tmp10372 = s7 ? tmp10373 : tmp10381;
  assign tmp10323 = s8 ? tmp10324 : tmp10372;
  assign tmp10393 = s4 ? tmp10384 : tmp9657;
  assign tmp10392 = s5 ? tmp10361 : tmp10393;
  assign tmp10391 = s6 ? tmp10357 : tmp10392;
  assign tmp10390 = s7 ? tmp10325 : tmp10391;
  assign tmp10389 = s8 ? tmp10372 : tmp10390;
  assign tmp10322 = s9 ? tmp10323 : tmp10389;
  assign tmp10400 = s3 ? tmp9657 : tmp10388;
  assign tmp10399 = s4 ? tmp10384 : tmp10400;
  assign tmp10398 = s5 ? tmp10361 : tmp10399;
  assign tmp10397 = s6 ? tmp10357 : tmp10398;
  assign tmp10396 = s7 ? tmp10325 : tmp10397;
  assign tmp10395 = s8 ? tmp10396 : tmp10325;
  assign tmp10405 = s4 ? tmp10369 : tmp10400;
  assign tmp10404 = s5 ? tmp10361 : tmp10405;
  assign tmp10403 = s6 ? tmp10357 : tmp10404;
  assign tmp10402 = s7 ? tmp10403 : tmp10391;
  assign tmp10406 = s7 ? tmp10381 : tmp10397;
  assign tmp10401 = s8 ? tmp10402 : tmp10406;
  assign tmp10394 = s9 ? tmp10395 : tmp10401;
  assign tmp10321 = s10 ? tmp10322 : tmp10394;
  assign tmp10410 = s7 ? tmp10356 : tmp10391;
  assign tmp10409 = s8 ? tmp10410 : tmp10406;
  assign tmp10408 = s9 ? tmp10395 : tmp10409;
  assign tmp10407 = s10 ? tmp10322 : tmp10408;
  assign tmp10320 = s11 ? tmp10321 : tmp10407;
  assign tmp10182 = s12 ? tmp10183 : tmp10320;
  assign tmp10424 = ~(l4 ? 1 : 0);
  assign tmp10423 = l3 ? 1 : tmp10424;
  assign tmp10422 = ~(l2 ? 1 : tmp10423);
  assign tmp10421 = l1 ? tmp9172 : tmp10422;
  assign tmp10425 = s0 ? 1 : tmp10421;
  assign tmp10420 = s1 ? tmp10421 : tmp10425;
  assign tmp10427 = s1 ? tmp9657 : tmp10421;
  assign tmp10426 = s2 ? tmp10421 : tmp10427;
  assign tmp10419 = s3 ? tmp10420 : tmp10426;
  assign tmp10432 = l1 ? 1 : tmp10422;
  assign tmp10431 = s0 ? tmp10432 : 1;
  assign tmp10430 = s1 ? tmp10431 : tmp10421;
  assign tmp10434 = s0 ? tmp10421 : tmp9151;
  assign tmp10433 = s1 ? tmp10434 : 1;
  assign tmp10429 = s2 ? tmp10430 : tmp10433;
  assign tmp10436 = s1 ? 1 : tmp9254;
  assign tmp10438 = s0 ? tmp9610 : tmp10421;
  assign tmp10437 = s1 ? tmp10421 : tmp10438;
  assign tmp10435 = s2 ? tmp10436 : tmp10437;
  assign tmp10428 = s3 ? tmp10429 : tmp10435;
  assign tmp10418 = s4 ? tmp10419 : tmp10428;
  assign tmp10444 = s0 ? tmp10421 : 1;
  assign tmp10443 = s1 ? tmp10444 : 1;
  assign tmp10445 = s1 ? tmp10425 : tmp10421;
  assign tmp10442 = s2 ? tmp10443 : tmp10445;
  assign tmp10447 = s1 ? tmp10229 : tmp10421;
  assign tmp10446 = s2 ? tmp10421 : tmp10447;
  assign tmp10441 = s3 ? tmp10442 : tmp10446;
  assign tmp10452 = ~(l1 ? tmp9172 : tmp10422);
  assign tmp10451 = s0 ? 1 : tmp10452;
  assign tmp10450 = s1 ? tmp10451 : 0;
  assign tmp10453 = ~(s1 ? 1 : tmp10431);
  assign tmp10449 = s2 ? tmp10450 : tmp10453;
  assign tmp10454 = ~(s2 ? tmp10420 : 0);
  assign tmp10448 = ~(s3 ? tmp10449 : tmp10454);
  assign tmp10440 = s4 ? tmp10441 : tmp10448;
  assign tmp10459 = s0 ? tmp10421 : 0;
  assign tmp10458 = s1 ? tmp10459 : tmp9618;
  assign tmp10457 = s2 ? tmp10458 : tmp9475;
  assign tmp10463 = ~(l1 ? 1 : tmp10422);
  assign tmp10462 = s0 ? 1 : tmp10463;
  assign tmp10461 = ~(s1 ? 1 : tmp10462);
  assign tmp10460 = s2 ? tmp9476 : tmp10461;
  assign tmp10456 = s3 ? tmp10457 : tmp10460;
  assign tmp10467 = s0 ? tmp10432 : tmp9610;
  assign tmp10466 = s1 ? tmp10467 : tmp9610;
  assign tmp10468 = ~(s1 ? tmp10451 : 0);
  assign tmp10465 = s2 ? tmp10466 : tmp10468;
  assign tmp10471 = ~(s0 ? 1 : tmp10452);
  assign tmp10470 = s1 ? tmp9610 : tmp10471;
  assign tmp10474 = ~(l1 ? tmp9172 : 0);
  assign tmp10473 = s0 ? 1 : tmp10474;
  assign tmp10472 = ~(s1 ? tmp10462 : tmp10473);
  assign tmp10469 = s2 ? tmp10470 : tmp10472;
  assign tmp10464 = s3 ? tmp10465 : tmp10469;
  assign tmp10455 = s4 ? tmp10456 : tmp10464;
  assign tmp10439 = s5 ? tmp10440 : tmp10455;
  assign tmp10417 = s6 ? tmp10418 : tmp10439;
  assign tmp10478 = s2 ? tmp9816 : tmp10437;
  assign tmp10477 = s3 ? tmp10429 : tmp10478;
  assign tmp10476 = s4 ? tmp10419 : tmp10477;
  assign tmp10482 = s2 ? tmp10443 : tmp10421;
  assign tmp10481 = s3 ? tmp10482 : tmp10446;
  assign tmp10484 = s2 ? tmp10450 : tmp10463;
  assign tmp10485 = ~(s2 ? tmp10421 : 0);
  assign tmp10483 = ~(s3 ? tmp10484 : tmp10485);
  assign tmp10480 = s4 ? tmp10481 : tmp10483;
  assign tmp10489 = s1 ? tmp10459 : tmp9172;
  assign tmp10488 = s2 ? tmp10489 : 1;
  assign tmp10491 = s1 ? 1 : tmp10463;
  assign tmp10490 = ~(s2 ? 1 : tmp10491);
  assign tmp10487 = s3 ? tmp10488 : tmp10490;
  assign tmp10493 = s2 ? tmp9610 : tmp10421;
  assign tmp10495 = s1 ? tmp9610 : tmp10421;
  assign tmp10494 = s2 ? tmp10495 : tmp9610;
  assign tmp10492 = s3 ? tmp10493 : tmp10494;
  assign tmp10486 = s4 ? tmp10487 : tmp10492;
  assign tmp10479 = s5 ? tmp10480 : tmp10486;
  assign tmp10475 = s6 ? tmp10476 : tmp10479;
  assign tmp10416 = s7 ? tmp10417 : tmp10475;
  assign tmp10502 = ~(l3 ? 1 : tmp10424);
  assign tmp10501 = l1 ? tmp9172 : tmp10502;
  assign tmp10503 = s0 ? 1 : tmp10501;
  assign tmp10500 = s1 ? tmp10501 : tmp10503;
  assign tmp10505 = s1 ? tmp9662 : tmp10501;
  assign tmp10504 = s2 ? tmp10501 : tmp10505;
  assign tmp10499 = s3 ? tmp10500 : tmp10504;
  assign tmp10510 = l1 ? 1 : tmp10502;
  assign tmp10509 = s0 ? tmp10510 : 1;
  assign tmp10508 = s1 ? tmp10509 : tmp10501;
  assign tmp10512 = s0 ? tmp10501 : tmp9151;
  assign tmp10511 = s1 ? tmp10512 : 1;
  assign tmp10507 = s2 ? tmp10508 : tmp10511;
  assign tmp10515 = s0 ? tmp9172 : tmp10501;
  assign tmp10514 = s1 ? tmp10501 : tmp10515;
  assign tmp10513 = s2 ? tmp10436 : tmp10514;
  assign tmp10506 = s3 ? tmp10507 : tmp10513;
  assign tmp10498 = s4 ? tmp10499 : tmp10506;
  assign tmp10521 = s0 ? tmp10501 : 1;
  assign tmp10520 = s1 ? tmp10521 : 1;
  assign tmp10522 = s1 ? tmp10503 : tmp10521;
  assign tmp10519 = s2 ? tmp10520 : tmp10522;
  assign tmp10524 = s1 ? tmp9186 : tmp10501;
  assign tmp10523 = s2 ? tmp10503 : tmp10524;
  assign tmp10518 = s3 ? tmp10519 : tmp10523;
  assign tmp10529 = ~(l1 ? tmp9172 : tmp10502);
  assign tmp10528 = s0 ? 1 : tmp10529;
  assign tmp10527 = s1 ? tmp10528 : 0;
  assign tmp10530 = ~(s1 ? 1 : tmp10509);
  assign tmp10526 = s2 ? tmp10527 : tmp10530;
  assign tmp10532 = s1 ? tmp10501 : tmp10425;
  assign tmp10531 = ~(s2 ? tmp10532 : 0);
  assign tmp10525 = ~(s3 ? tmp10526 : tmp10531);
  assign tmp10517 = s4 ? tmp10518 : tmp10525;
  assign tmp10537 = s0 ? tmp10501 : 0;
  assign tmp10536 = s1 ? tmp10537 : tmp9839;
  assign tmp10535 = s2 ? tmp10536 : tmp9689;
  assign tmp10534 = s3 ? tmp10535 : tmp10460;
  assign tmp10540 = s1 ? tmp10467 : tmp9622;
  assign tmp10541 = ~(s1 ? tmp10528 : 0);
  assign tmp10539 = s2 ? tmp10540 : tmp10541;
  assign tmp10544 = s0 ? tmp9657 : tmp9610;
  assign tmp10543 = s1 ? tmp10544 : tmp10471;
  assign tmp10542 = s2 ? tmp10543 : tmp10472;
  assign tmp10538 = s3 ? tmp10539 : tmp10542;
  assign tmp10533 = s4 ? tmp10534 : tmp10538;
  assign tmp10516 = s5 ? tmp10517 : tmp10533;
  assign tmp10497 = s6 ? tmp10498 : tmp10516;
  assign tmp10548 = s2 ? tmp9816 : tmp10514;
  assign tmp10547 = s3 ? tmp10507 : tmp10548;
  assign tmp10546 = s4 ? tmp10499 : tmp10547;
  assign tmp10553 = s1 ? tmp10501 : tmp10521;
  assign tmp10552 = s2 ? tmp10520 : tmp10553;
  assign tmp10554 = s2 ? tmp10501 : tmp10524;
  assign tmp10551 = s3 ? tmp10552 : tmp10554;
  assign tmp10557 = ~(l1 ? 1 : tmp10502);
  assign tmp10556 = s2 ? tmp10527 : tmp10557;
  assign tmp10559 = s1 ? tmp10501 : tmp10421;
  assign tmp10558 = ~(s2 ? tmp10559 : 0);
  assign tmp10555 = ~(s3 ? tmp10556 : tmp10558);
  assign tmp10550 = s4 ? tmp10551 : tmp10555;
  assign tmp10563 = s1 ? tmp10537 : tmp9657;
  assign tmp10562 = s2 ? tmp10563 : 1;
  assign tmp10561 = s3 ? tmp10562 : tmp10490;
  assign tmp10566 = s1 ? tmp9610 : tmp9622;
  assign tmp10565 = s2 ? tmp10566 : tmp10501;
  assign tmp10564 = s3 ? tmp10565 : tmp10494;
  assign tmp10560 = s4 ? tmp10561 : tmp10564;
  assign tmp10549 = s5 ? tmp10550 : tmp10560;
  assign tmp10545 = s6 ? tmp10546 : tmp10549;
  assign tmp10496 = s7 ? tmp10497 : tmp10545;
  assign tmp10415 = s8 ? tmp10416 : tmp10496;
  assign tmp10573 = s0 ? 1 : tmp9610;
  assign tmp10572 = s1 ? tmp9610 : tmp10573;
  assign tmp10575 = s1 ? tmp9433 : tmp9610;
  assign tmp10574 = s2 ? tmp9610 : tmp10575;
  assign tmp10571 = s3 ? tmp10572 : tmp10574;
  assign tmp10578 = s1 ? tmp9159 : tmp9610;
  assign tmp10580 = s0 ? tmp9610 : tmp9151;
  assign tmp10579 = s1 ? tmp10580 : 1;
  assign tmp10577 = s2 ? tmp10578 : tmp10579;
  assign tmp10581 = s2 ? tmp10436 : tmp9610;
  assign tmp10576 = s3 ? tmp10577 : tmp10581;
  assign tmp10570 = s4 ? tmp10571 : tmp10576;
  assign tmp10586 = s1 ? tmp10573 : tmp9648;
  assign tmp10585 = s2 ? tmp9647 : tmp10586;
  assign tmp10588 = s1 ? tmp10229 : tmp9610;
  assign tmp10587 = s2 ? tmp10573 : tmp10588;
  assign tmp10584 = s3 ? tmp10585 : tmp10587;
  assign tmp10591 = s1 ? tmp10473 : 0;
  assign tmp10590 = s2 ? tmp10591 : tmp9258;
  assign tmp10594 = s0 ? tmp9151 : tmp9610;
  assign tmp10593 = s1 ? tmp9610 : tmp10594;
  assign tmp10592 = ~(s2 ? tmp10593 : 0);
  assign tmp10589 = ~(s3 ? tmp10590 : tmp10592);
  assign tmp10583 = s4 ? tmp10584 : tmp10589;
  assign tmp10598 = s1 ? tmp10229 : tmp9618;
  assign tmp10597 = s2 ? tmp10598 : tmp9172;
  assign tmp10596 = s3 ? tmp10597 : tmp9546;
  assign tmp10601 = ~(s1 ? tmp10473 : 0);
  assign tmp10600 = s2 ? tmp9610 : tmp10601;
  assign tmp10604 = ~(s0 ? 1 : tmp10474);
  assign tmp10603 = s1 ? tmp9610 : tmp10604;
  assign tmp10602 = s2 ? tmp10603 : tmp10604;
  assign tmp10599 = s3 ? tmp10600 : tmp10602;
  assign tmp10595 = s4 ? tmp10596 : tmp10599;
  assign tmp10582 = s5 ? tmp10583 : tmp10595;
  assign tmp10569 = s6 ? tmp10570 : tmp10582;
  assign tmp10608 = s2 ? tmp9816 : tmp9610;
  assign tmp10607 = s3 ? tmp10577 : tmp10608;
  assign tmp10606 = s4 ? tmp10571 : tmp10607;
  assign tmp10613 = s1 ? tmp9610 : tmp9648;
  assign tmp10612 = s2 ? tmp9647 : tmp10613;
  assign tmp10614 = s2 ? tmp9610 : tmp10588;
  assign tmp10611 = s3 ? tmp10612 : tmp10614;
  assign tmp10616 = s2 ? tmp10591 : tmp9257;
  assign tmp10617 = ~(s2 ? tmp9610 : 0);
  assign tmp10615 = ~(s3 ? tmp10616 : tmp10617);
  assign tmp10610 = s4 ? tmp10611 : tmp10615;
  assign tmp10621 = s1 ? tmp10229 : tmp9172;
  assign tmp10620 = s2 ? tmp10621 : 1;
  assign tmp10619 = s3 ? tmp10620 : tmp9565;
  assign tmp10618 = s4 ? tmp10619 : tmp9610;
  assign tmp10609 = s5 ? tmp10610 : tmp10618;
  assign tmp10605 = s6 ? tmp10606 : tmp10609;
  assign tmp10568 = s7 ? tmp10569 : tmp10605;
  assign tmp10567 = s8 ? tmp10496 : tmp10568;
  assign tmp10414 = s9 ? tmp10415 : tmp10567;
  assign tmp10629 = s1 ? tmp9662 : tmp10421;
  assign tmp10628 = s2 ? tmp10421 : tmp10629;
  assign tmp10627 = s3 ? tmp10420 : tmp10628;
  assign tmp10634 = ~(l2 ? tmp10423 : 1);
  assign tmp10633 = s0 ? tmp10421 : tmp10634;
  assign tmp10632 = s1 ? tmp10633 : 1;
  assign tmp10631 = s2 ? tmp10430 : tmp10632;
  assign tmp10630 = s3 ? tmp10631 : tmp10435;
  assign tmp10626 = s4 ? tmp10627 : tmp10630;
  assign tmp10639 = s1 ? tmp10425 : tmp10444;
  assign tmp10638 = s2 ? tmp10443 : tmp10639;
  assign tmp10640 = s2 ? tmp10425 : tmp10447;
  assign tmp10637 = s3 ? tmp10638 : tmp10640;
  assign tmp10644 = s0 ? tmp9151 : tmp10421;
  assign tmp10643 = s1 ? tmp10421 : tmp10644;
  assign tmp10642 = ~(s2 ? tmp10643 : 0);
  assign tmp10641 = ~(s3 ? tmp10449 : tmp10642);
  assign tmp10636 = s4 ? tmp10637 : tmp10641;
  assign tmp10635 = s5 ? tmp10636 : tmp10455;
  assign tmp10625 = s6 ? tmp10626 : tmp10635;
  assign tmp10647 = s3 ? tmp10631 : tmp10478;
  assign tmp10646 = s4 ? tmp10627 : tmp10647;
  assign tmp10652 = s1 ? tmp10421 : tmp10444;
  assign tmp10651 = s2 ? tmp10443 : tmp10652;
  assign tmp10650 = s3 ? tmp10651 : tmp10446;
  assign tmp10649 = s4 ? tmp10650 : tmp10483;
  assign tmp10648 = s5 ? tmp10649 : tmp10486;
  assign tmp10645 = s6 ? tmp10646 : tmp10648;
  assign tmp10624 = s7 ? tmp10625 : tmp10645;
  assign tmp10623 = s8 ? tmp10624 : tmp10625;
  assign tmp10658 = s3 ? tmp10493 : tmp10495;
  assign tmp10657 = s4 ? tmp10487 : tmp10658;
  assign tmp10656 = s5 ? tmp10480 : tmp10657;
  assign tmp10655 = s6 ? tmp10476 : tmp10656;
  assign tmp10654 = s7 ? tmp10655 : tmp10605;
  assign tmp10663 = s3 ? tmp10565 : tmp10495;
  assign tmp10662 = s4 ? tmp10561 : tmp10663;
  assign tmp10661 = s5 ? tmp10550 : tmp10662;
  assign tmp10660 = s6 ? tmp10546 : tmp10661;
  assign tmp10665 = s5 ? tmp10649 : tmp10657;
  assign tmp10664 = s6 ? tmp10646 : tmp10665;
  assign tmp10659 = s7 ? tmp10660 : tmp10664;
  assign tmp10653 = s8 ? tmp10654 : tmp10659;
  assign tmp10622 = s9 ? tmp10623 : tmp10653;
  assign tmp10413 = s10 ? tmp10414 : tmp10622;
  assign tmp10669 = s7 ? tmp10475 : tmp10605;
  assign tmp10670 = s7 ? tmp10545 : tmp10645;
  assign tmp10668 = s8 ? tmp10669 : tmp10670;
  assign tmp10667 = s9 ? tmp10623 : tmp10668;
  assign tmp10666 = s10 ? tmp10414 : tmp10667;
  assign tmp10412 = ~(s11 ? tmp10413 : tmp10666);
  assign tmp10411 = ~(s12 ? 1 : tmp10412);
  assign tmp10181 = s13 ? tmp10182 : tmp10411;
  assign tmp9898 = ~(s14 ? tmp9899 : tmp10181);
  assign tmp9136 = s15 ? tmp9137 : tmp9898;
  assign tmp10683 = s2 ? tmp9181 : tmp9187;
  assign tmp10682 = s3 ? tmp10683 : 0;
  assign tmp10681 = ~(s4 ? tmp10682 : tmp9209);
  assign tmp10680 = s5 ? tmp9166 : tmp10681;
  assign tmp10679 = s6 ? tmp9145 : tmp10680;
  assign tmp10687 = s3 ? tmp9181 : 0;
  assign tmp10686 = ~(s4 ? tmp10687 : tmp9209);
  assign tmp10685 = s5 ? tmp9198 : tmp10686;
  assign tmp10684 = s6 ? tmp9193 : tmp10685;
  assign tmp10678 = s7 ? tmp10679 : tmp10684;
  assign tmp10695 = s0 ? tmp9148 : 0;
  assign tmp10694 = s1 ? tmp9150 : tmp10695;
  assign tmp10693 = s2 ? tmp9169 : tmp10694;
  assign tmp10698 = s0 ? 1 : tmp9320;
  assign tmp10697 = s1 ? tmp10698 : tmp9174;
  assign tmp10696 = ~(s2 ? tmp10697 : tmp9175);
  assign tmp10692 = s3 ? tmp10693 : tmp10696;
  assign tmp10691 = s4 ? tmp10692 : tmp9226;
  assign tmp10690 = s5 ? tmp10691 : tmp10681;
  assign tmp10689 = s6 ? tmp9213 : tmp10690;
  assign tmp10704 = s1 ? tmp9148 : tmp10695;
  assign tmp10703 = s2 ? tmp9153 : tmp10704;
  assign tmp10702 = s3 ? tmp10703 : tmp9236;
  assign tmp10708 = ~(s0 ? tmp9148 : tmp9659);
  assign tmp10707 = ~(s1 ? tmp9657 : tmp10708);
  assign tmp10706 = s2 ? tmp9178 : tmp10707;
  assign tmp10705 = s3 ? tmp10706 : tmp9227;
  assign tmp10701 = s4 ? tmp10702 : tmp10705;
  assign tmp10700 = s5 ? tmp10701 : tmp10686;
  assign tmp10699 = s6 ? tmp9229 : tmp10700;
  assign tmp10688 = s7 ? tmp10689 : tmp10699;
  assign tmp10677 = s8 ? tmp10678 : tmp10688;
  assign tmp10714 = s2 ? tmp9657 : tmp9695;
  assign tmp10716 = s1 ? tmp9657 : tmp9186;
  assign tmp10715 = s2 ? tmp10716 : tmp10354;
  assign tmp10713 = s3 ? tmp10714 : tmp10715;
  assign tmp10712 = s4 ? tmp9657 : tmp10713;
  assign tmp10721 = s1 ? tmp9666 : tmp9658;
  assign tmp10722 = ~(s1 ? tmp10342 : tmp9659);
  assign tmp10720 = s2 ? tmp10721 : tmp10722;
  assign tmp10724 = s1 ? tmp9657 : tmp9256;
  assign tmp10726 = ~(s0 ? tmp9657 : tmp9172);
  assign tmp10725 = ~(s1 ? 1 : tmp10726);
  assign tmp10723 = s2 ? tmp10724 : tmp10725;
  assign tmp10719 = s3 ? tmp10720 : tmp10723;
  assign tmp10729 = s1 ? tmp9841 : tmp10726;
  assign tmp10730 = ~(s1 ? tmp9695 : tmp9657);
  assign tmp10728 = s2 ? tmp10729 : tmp10730;
  assign tmp10731 = s2 ? tmp9930 : 1;
  assign tmp10727 = ~(s3 ? tmp10728 : tmp10731);
  assign tmp10718 = s4 ? tmp10719 : tmp10727;
  assign tmp10734 = s2 ? tmp9161 : tmp9268;
  assign tmp10733 = s3 ? tmp10734 : 1;
  assign tmp10732 = ~(s4 ? tmp10733 : tmp9283);
  assign tmp10717 = s5 ? tmp10718 : tmp10732;
  assign tmp10711 = s6 ? tmp10712 : tmp10717;
  assign tmp10739 = s1 ? tmp9695 : tmp9657;
  assign tmp10738 = s2 ? tmp9657 : tmp10739;
  assign tmp10740 = s2 ? tmp9921 : tmp10354;
  assign tmp10737 = s3 ? tmp10738 : tmp10740;
  assign tmp10736 = s4 ? tmp9657 : tmp10737;
  assign tmp10744 = s2 ? tmp9665 : tmp9657;
  assign tmp10746 = s1 ? tmp9657 : tmp9257;
  assign tmp10745 = s2 ? tmp10746 : tmp10725;
  assign tmp10743 = s3 ? tmp10744 : tmp10745;
  assign tmp10748 = s2 ? tmp10729 : tmp9659;
  assign tmp10750 = s1 ? tmp9224 : 1;
  assign tmp10749 = s2 ? tmp10750 : 1;
  assign tmp10747 = ~(s3 ? tmp10748 : tmp10749);
  assign tmp10742 = s4 ? tmp10743 : tmp10747;
  assign tmp10752 = s3 ? tmp9161 : 1;
  assign tmp10751 = ~(s4 ? tmp10752 : tmp9283);
  assign tmp10741 = s5 ? tmp10742 : tmp10751;
  assign tmp10735 = s6 ? tmp10736 : tmp10741;
  assign tmp10710 = ~(s7 ? tmp10711 : tmp10735);
  assign tmp10709 = s8 ? tmp10688 : tmp10710;
  assign tmp10676 = s9 ? tmp10677 : tmp10709;
  assign tmp10760 = s1 ? tmp9691 : tmp9172;
  assign tmp10759 = s2 ? tmp9172 : tmp10760;
  assign tmp10758 = s3 ? tmp10255 : tmp10759;
  assign tmp10762 = s2 ? tmp10760 : tmp10255;
  assign tmp10763 = s2 ? tmp10716 : tmp9806;
  assign tmp10761 = s3 ? tmp10762 : tmp10763;
  assign tmp10757 = s4 ? tmp10758 : tmp10761;
  assign tmp10768 = s1 ? tmp9599 : tmp9454;
  assign tmp10769 = ~(s1 ? tmp9224 : tmp9171);
  assign tmp10767 = s2 ? tmp10768 : tmp10769;
  assign tmp10772 = ~(s0 ? tmp9172 : tmp9610);
  assign tmp10771 = ~(s1 ? 1 : tmp10772);
  assign tmp10770 = s2 ? tmp9174 : tmp10771;
  assign tmp10766 = s3 ? tmp10767 : tmp10770;
  assign tmp10775 = s1 ? tmp9188 : tmp10726;
  assign tmp10776 = ~(s1 ? tmp9695 : tmp9691);
  assign tmp10774 = s2 ? tmp10775 : tmp10776;
  assign tmp10778 = s1 ? tmp9609 : tmp9186;
  assign tmp10777 = ~(s2 ? tmp10778 : 0);
  assign tmp10773 = ~(s3 ? tmp10774 : tmp10777);
  assign tmp10765 = s4 ? tmp10766 : tmp10773;
  assign tmp10779 = s4 ? tmp10682 : tmp9209;
  assign tmp10764 = s5 ? tmp10765 : tmp10779;
  assign tmp10756 = s6 ? tmp10757 : tmp10764;
  assign tmp10783 = s2 ? tmp10760 : tmp10388;
  assign tmp10784 = s2 ? tmp9921 : tmp9806;
  assign tmp10782 = s3 ? tmp10783 : tmp10784;
  assign tmp10781 = s4 ? tmp10758 : tmp10782;
  assign tmp10788 = s2 ? tmp9598 : tmp9636;
  assign tmp10789 = s2 ? tmp9172 : tmp10771;
  assign tmp10787 = s3 ? tmp10788 : tmp10789;
  assign tmp10792 = ~(s1 ? tmp9657 : tmp9691);
  assign tmp10791 = s2 ? tmp10775 : tmp10792;
  assign tmp10794 = s1 ? tmp9609 : 0;
  assign tmp10793 = ~(s2 ? tmp10794 : 0);
  assign tmp10790 = ~(s3 ? tmp10791 : tmp10793);
  assign tmp10786 = s4 ? tmp10787 : tmp10790;
  assign tmp10795 = s4 ? tmp10687 : tmp9209;
  assign tmp10785 = s5 ? tmp10786 : tmp10795;
  assign tmp10780 = s6 ? tmp10781 : tmp10785;
  assign tmp10755 = s7 ? tmp10756 : tmp10780;
  assign tmp10754 = s8 ? tmp10755 : tmp10756;
  assign tmp10799 = s5 ? tmp9296 : tmp10686;
  assign tmp10798 = s6 ? tmp9193 : tmp10799;
  assign tmp10800 = ~(s6 ? tmp10736 : tmp10741);
  assign tmp10797 = s7 ? tmp10798 : tmp10800;
  assign tmp10807 = ~(s1 ? tmp9657 : tmp9320);
  assign tmp10806 = s2 ? tmp9178 : tmp10807;
  assign tmp10805 = s3 ? tmp10806 : tmp9227;
  assign tmp10804 = s4 ? tmp10702 : tmp10805;
  assign tmp10803 = s5 ? tmp10804 : tmp10686;
  assign tmp10802 = s6 ? tmp9229 : tmp10803;
  assign tmp10813 = ~(s1 ? tmp9657 : tmp9172);
  assign tmp10812 = s2 ? tmp10775 : tmp10813;
  assign tmp10811 = ~(s3 ? tmp10812 : tmp10793);
  assign tmp10810 = s4 ? tmp10787 : tmp10811;
  assign tmp10809 = s5 ? tmp10810 : tmp10795;
  assign tmp10808 = ~(s6 ? tmp10781 : tmp10809);
  assign tmp10801 = s7 ? tmp10802 : tmp10808;
  assign tmp10796 = ~(s8 ? tmp10797 : tmp10801);
  assign tmp10753 = ~(s9 ? tmp10754 : tmp10796);
  assign tmp10675 = s10 ? tmp10676 : tmp10753;
  assign tmp10817 = s7 ? tmp10684 : tmp10800;
  assign tmp10819 = ~(s6 ? tmp10781 : tmp10785);
  assign tmp10818 = s7 ? tmp10699 : tmp10819;
  assign tmp10816 = ~(s8 ? tmp10817 : tmp10818);
  assign tmp10815 = ~(s9 ? tmp10754 : tmp10816);
  assign tmp10814 = s10 ? tmp10676 : tmp10815;
  assign tmp10674 = s11 ? tmp10675 : tmp10814;
  assign tmp10830 = s1 ? 1 : tmp9350;
  assign tmp10829 = s2 ? tmp9796 : tmp10830;
  assign tmp10828 = s3 ? 1 : tmp10829;
  assign tmp10827 = s4 ? 1 : tmp10828;
  assign tmp10835 = ~(s1 ? 1 : tmp9350);
  assign tmp10834 = s2 ? tmp9796 : tmp10835;
  assign tmp10833 = s3 ? 1 : tmp10834;
  assign tmp10838 = ~(s1 ? tmp9317 : 1);
  assign tmp10837 = s2 ? tmp9349 : tmp10838;
  assign tmp10836 = ~(s3 ? tmp10837 : 1);
  assign tmp10832 = s4 ? tmp10833 : tmp10836;
  assign tmp10831 = s5 ? tmp10832 : 0;
  assign tmp10826 = s6 ? tmp10827 : tmp10831;
  assign tmp10843 = s2 ? tmp9816 : tmp10835;
  assign tmp10842 = s3 ? 1 : tmp10843;
  assign tmp10845 = s2 ? tmp9349 : 0;
  assign tmp10844 = ~(s3 ? tmp10845 : 1);
  assign tmp10841 = s4 ? tmp10842 : tmp10844;
  assign tmp10840 = s5 ? tmp10841 : 0;
  assign tmp10839 = s6 ? tmp10827 : tmp10840;
  assign tmp10825 = s7 ? tmp10826 : tmp10839;
  assign tmp10852 = ~(s1 ? 1 : 0);
  assign tmp10851 = s2 ? tmp9796 : tmp10852;
  assign tmp10850 = s3 ? 1 : tmp10851;
  assign tmp10854 = s2 ? tmp9476 : 0;
  assign tmp10853 = ~(s3 ? tmp10854 : 1);
  assign tmp10849 = s4 ? tmp10850 : tmp10853;
  assign tmp10848 = s5 ? tmp10849 : 0;
  assign tmp10847 = s6 ? tmp10827 : tmp10848;
  assign tmp10859 = s1 ? 1 : tmp10473;
  assign tmp10858 = s2 ? 1 : tmp10859;
  assign tmp10862 = ~(s0 ? tmp9610 : 1);
  assign tmp10861 = s1 ? 1 : tmp10862;
  assign tmp10860 = s2 ? tmp10861 : tmp10830;
  assign tmp10857 = s3 ? tmp10858 : tmp10860;
  assign tmp10856 = s4 ? 1 : tmp10857;
  assign tmp10866 = s2 ? tmp9816 : tmp10852;
  assign tmp10865 = s3 ? 1 : tmp10866;
  assign tmp10864 = s4 ? tmp10865 : tmp10853;
  assign tmp10863 = s5 ? tmp10864 : 0;
  assign tmp10855 = s6 ? tmp10856 : tmp10863;
  assign tmp10846 = s7 ? tmp10847 : tmp10855;
  assign tmp10824 = s8 ? tmp10825 : tmp10846;
  assign tmp10872 = s2 ? tmp10613 : tmp10572;
  assign tmp10871 = s3 ? tmp9610 : tmp10872;
  assign tmp10870 = s4 ? tmp9610 : tmp10871;
  assign tmp10877 = s1 ? tmp10229 : tmp10604;
  assign tmp10878 = ~(s1 ? tmp9188 : tmp9257);
  assign tmp10876 = s2 ? tmp10877 : tmp10878;
  assign tmp10880 = s1 ? tmp9151 : tmp9159;
  assign tmp10879 = s2 ? tmp10880 : tmp9425;
  assign tmp10875 = s3 ? tmp10876 : tmp10879;
  assign tmp10882 = s2 ? tmp9811 : tmp9172;
  assign tmp10881 = s3 ? tmp10882 : 1;
  assign tmp10874 = s4 ? tmp10875 : tmp10881;
  assign tmp10873 = s5 ? tmp10874 : 1;
  assign tmp10869 = s6 ? tmp10870 : tmp10873;
  assign tmp10888 = s1 ? tmp9172 : tmp9151;
  assign tmp10887 = s2 ? tmp10588 : tmp10888;
  assign tmp10889 = s2 ? tmp9161 : tmp9425;
  assign tmp10886 = s3 ? tmp10887 : tmp10889;
  assign tmp10885 = s4 ? tmp10886 : tmp10881;
  assign tmp10884 = s5 ? tmp10885 : 1;
  assign tmp10883 = s6 ? tmp10870 : tmp10884;
  assign tmp10868 = ~(s7 ? tmp10869 : tmp10883);
  assign tmp10867 = s8 ? tmp10846 : tmp10868;
  assign tmp10823 = s9 ? tmp10824 : tmp10867;
  assign tmp10892 = s7 ? tmp10869 : tmp10883;
  assign tmp10891 = s8 ? tmp10892 : tmp10869;
  assign tmp10898 = s2 ? tmp9816 : tmp10830;
  assign tmp10897 = s3 ? 1 : tmp10898;
  assign tmp10896 = s4 ? 1 : tmp10897;
  assign tmp10895 = s6 ? tmp10896 : tmp10840;
  assign tmp10903 = s1 ? tmp9610 : 1;
  assign tmp10902 = s2 ? tmp10903 : tmp10572;
  assign tmp10901 = s3 ? tmp9610 : tmp10902;
  assign tmp10900 = s4 ? tmp9610 : tmp10901;
  assign tmp10899 = ~(s6 ? tmp10900 : tmp10884);
  assign tmp10894 = s7 ? tmp10895 : tmp10899;
  assign tmp10907 = s3 ? tmp10858 : tmp10898;
  assign tmp10906 = s4 ? 1 : tmp10907;
  assign tmp10905 = s6 ? tmp10906 : tmp10863;
  assign tmp10904 = s7 ? tmp10905 : tmp10899;
  assign tmp10893 = ~(s8 ? tmp10894 : tmp10904);
  assign tmp10890 = ~(s9 ? tmp10891 : tmp10893);
  assign tmp10822 = s10 ? tmp10823 : tmp10890;
  assign tmp10912 = ~(s6 ? tmp10870 : tmp10884);
  assign tmp10911 = s7 ? tmp10839 : tmp10912;
  assign tmp10913 = s7 ? tmp10855 : tmp10912;
  assign tmp10910 = ~(s8 ? tmp10911 : tmp10913);
  assign tmp10909 = ~(s9 ? tmp10891 : tmp10910);
  assign tmp10908 = s10 ? tmp10823 : tmp10909;
  assign tmp10821 = s11 ? tmp10822 : tmp10908;
  assign tmp10820 = s12 ? tmp9306 : tmp10821;
  assign tmp10673 = s13 ? tmp10674 : tmp10820;
  assign tmp10924 = s2 ? tmp9969 : tmp9971;
  assign tmp10926 = s1 ? tmp9969 : tmp9159;
  assign tmp10927 = s1 ? tmp9969 : tmp9984;
  assign tmp10925 = s2 ? tmp10926 : tmp10927;
  assign tmp10923 = s3 ? tmp10924 : tmp10925;
  assign tmp10922 = s4 ? tmp9969 : tmp10923;
  assign tmp10933 = s0 ? tmp9969 : tmp9172;
  assign tmp10934 = s0 ? tmp9172 : tmp9969;
  assign tmp10932 = s1 ? tmp10933 : tmp10934;
  assign tmp10935 = s1 ? tmp9433 : tmp9969;
  assign tmp10931 = s2 ? tmp10932 : tmp10935;
  assign tmp10938 = s0 ? tmp9969 : 1;
  assign tmp10937 = s1 ? tmp9969 : tmp10938;
  assign tmp10936 = s2 ? tmp10937 : 1;
  assign tmp10930 = s3 ? tmp10931 : tmp10936;
  assign tmp10929 = s4 ? tmp10930 : 1;
  assign tmp10928 = s5 ? tmp10929 : 1;
  assign tmp10921 = s6 ? tmp10922 : tmp10928;
  assign tmp10943 = s1 ? tmp9971 : 1;
  assign tmp10942 = s2 ? tmp9969 : tmp10943;
  assign tmp10945 = s1 ? tmp9969 : 1;
  assign tmp10944 = s2 ? tmp10945 : tmp10927;
  assign tmp10941 = s3 ? tmp10942 : tmp10944;
  assign tmp10940 = s4 ? tmp9969 : tmp10941;
  assign tmp10950 = s1 ? tmp10933 : tmp9969;
  assign tmp10951 = s1 ? 1 : tmp9969;
  assign tmp10949 = s2 ? tmp10950 : tmp10951;
  assign tmp10948 = s3 ? tmp10949 : tmp10936;
  assign tmp10947 = s4 ? tmp10948 : 1;
  assign tmp10946 = s5 ? tmp10947 : 1;
  assign tmp10939 = s6 ? tmp10940 : tmp10946;
  assign tmp10920 = s7 ? tmp10921 : tmp10939;
  assign tmp10919 = s8 ? tmp9405 : tmp10920;
  assign tmp10918 = s9 ? tmp10919 : tmp10920;
  assign tmp10953 = s8 ? tmp10920 : tmp10921;
  assign tmp10960 = s2 ? tmp10945 : 1;
  assign tmp10959 = s3 ? tmp10949 : tmp10960;
  assign tmp10958 = s4 ? tmp10959 : 1;
  assign tmp10957 = s5 ? tmp10958 : 1;
  assign tmp10956 = s6 ? tmp10940 : tmp10957;
  assign tmp10955 = s7 ? tmp9438 : tmp10956;
  assign tmp10954 = s8 ? tmp10955 : tmp10956;
  assign tmp10952 = s9 ? tmp10953 : tmp10954;
  assign tmp10917 = s10 ? tmp10918 : tmp10952;
  assign tmp10964 = s7 ? tmp9417 : tmp10939;
  assign tmp10963 = s8 ? tmp10964 : tmp10939;
  assign tmp10962 = s9 ? tmp10953 : tmp10963;
  assign tmp10961 = s10 ? tmp10918 : tmp10962;
  assign tmp10916 = s11 ? tmp10917 : tmp10961;
  assign tmp10973 = s2 ? tmp9456 : tmp9600;
  assign tmp10972 = s3 ? tmp10973 : tmp9490;
  assign tmp10971 = s4 ? tmp9595 : tmp10972;
  assign tmp10978 = s1 ? tmp9433 : tmp9317;
  assign tmp10977 = s2 ? tmp10978 : tmp9606;
  assign tmp10979 = s2 ? tmp9174 : tmp9425;
  assign tmp10976 = s3 ? tmp10977 : tmp10979;
  assign tmp10975 = s4 ? tmp10976 : tmp9466;
  assign tmp10974 = s5 ? tmp10975 : tmp9472;
  assign tmp10970 = s6 ? tmp10971 : tmp10974;
  assign tmp10983 = s2 ? tmp9456 : tmp9631;
  assign tmp10982 = s3 ? tmp10983 : tmp9490;
  assign tmp10981 = s4 ? tmp9595 : tmp10982;
  assign tmp10988 = s1 ? tmp9433 : 0;
  assign tmp10987 = s2 ? tmp10988 : tmp9636;
  assign tmp10986 = s3 ? tmp10987 : tmp9424;
  assign tmp10985 = s4 ? tmp10986 : tmp9496;
  assign tmp10984 = s5 ? tmp10985 : tmp9499;
  assign tmp10980 = s6 ? tmp10981 : tmp10984;
  assign tmp10969 = s7 ? tmp10970 : tmp10980;
  assign tmp10992 = s3 ? tmp10255 : tmp9431;
  assign tmp10995 = s1 ? tmp9433 : tmp9662;
  assign tmp10994 = s2 ? tmp9172 : tmp10995;
  assign tmp10997 = s1 ? tmp9657 : 1;
  assign tmp10996 = s2 ? tmp10997 : tmp9412;
  assign tmp10993 = s3 ? tmp10994 : tmp10996;
  assign tmp10991 = s4 ? tmp10992 : tmp10993;
  assign tmp11000 = s3 ? tmp9604 : tmp10979;
  assign tmp11002 = s2 ? tmp10351 : tmp9710;
  assign tmp11003 = s2 ? tmp10255 : 1;
  assign tmp11001 = s3 ? tmp11002 : tmp11003;
  assign tmp10999 = s4 ? tmp11000 : tmp11001;
  assign tmp11006 = s2 ? tmp9475 : tmp9811;
  assign tmp11005 = s3 ? tmp11006 : tmp9477;
  assign tmp11007 = s3 ? tmp11006 : tmp9482;
  assign tmp11004 = s4 ? tmp11005 : tmp11007;
  assign tmp10998 = s5 ? tmp10999 : tmp11004;
  assign tmp10990 = s6 ? tmp10991 : tmp10998;
  assign tmp11012 = s1 ? tmp9433 : tmp9657;
  assign tmp11011 = s2 ? tmp9172 : tmp11012;
  assign tmp11010 = s3 ? tmp11011 : tmp10996;
  assign tmp11009 = s4 ? tmp10992 : tmp11010;
  assign tmp11015 = s3 ? tmp9635 : tmp9424;
  assign tmp11014 = s4 ? tmp11015 : tmp11001;
  assign tmp11018 = s2 ? tmp9475 : tmp9181;
  assign tmp11017 = s3 ? tmp11018 : tmp9502;
  assign tmp11016 = s4 ? tmp11017 : tmp9503;
  assign tmp11013 = s5 ? tmp11014 : tmp11016;
  assign tmp11008 = s6 ? tmp11009 : tmp11013;
  assign tmp10989 = s7 ? tmp10990 : tmp11008;
  assign tmp10968 = s8 ? tmp10969 : tmp10989;
  assign tmp11024 = s2 ? tmp9657 : tmp9662;
  assign tmp11025 = s2 ? tmp10997 : tmp10328;
  assign tmp11023 = s3 ? tmp11024 : tmp11025;
  assign tmp11022 = s4 ? tmp9657 : tmp11023;
  assign tmp11029 = s2 ? tmp9675 : tmp10330;
  assign tmp11030 = s2 ? tmp10724 : tmp9678;
  assign tmp11028 = s3 ? tmp11029 : tmp11030;
  assign tmp11032 = s2 ? tmp10330 : tmp9657;
  assign tmp11034 = s1 ? tmp10342 : tmp9683;
  assign tmp11033 = ~(s2 ? tmp11034 : 0);
  assign tmp11031 = s3 ? tmp11032 : tmp11033;
  assign tmp11027 = s4 ? tmp11028 : tmp11031;
  assign tmp11038 = ~(s1 ? tmp9256 : tmp9257);
  assign tmp11037 = s2 ? tmp9544 : tmp11038;
  assign tmp11036 = s3 ? tmp11037 : tmp9546;
  assign tmp11039 = s3 ? tmp11037 : tmp9551;
  assign tmp11035 = ~(s4 ? tmp11036 : tmp11039);
  assign tmp11026 = s5 ? tmp11027 : tmp11035;
  assign tmp11021 = s6 ? tmp11022 : tmp11026;
  assign tmp11042 = s3 ? tmp9660 : tmp11025;
  assign tmp11041 = s4 ? tmp9657 : tmp11042;
  assign tmp11046 = s2 ? tmp9661 : tmp9657;
  assign tmp11047 = s2 ? tmp10746 : tmp9678;
  assign tmp11045 = s3 ? tmp11046 : tmp11047;
  assign tmp11044 = s4 ? tmp11045 : tmp11031;
  assign tmp11050 = s2 ? tmp9544 : tmp9161;
  assign tmp11049 = s3 ? tmp11050 : tmp9565;
  assign tmp11048 = ~(s4 ? tmp11049 : tmp9567);
  assign tmp11043 = s5 ? tmp11044 : tmp11048;
  assign tmp11040 = s6 ? tmp11041 : tmp11043;
  assign tmp11020 = s7 ? tmp11021 : tmp11040;
  assign tmp11019 = s8 ? tmp10989 : tmp11020;
  assign tmp10967 = s9 ? tmp10968 : tmp11019;
  assign tmp11052 = s8 ? tmp10989 : tmp10990;
  assign tmp11057 = s4 ? tmp10986 : tmp9580;
  assign tmp11056 = s5 ? tmp11057 : tmp9499;
  assign tmp11055 = s6 ? tmp10981 : tmp11056;
  assign tmp11063 = s1 ? tmp10342 : tmp9151;
  assign tmp11062 = ~(s2 ? tmp11063 : 0);
  assign tmp11061 = s3 ? tmp11032 : tmp11062;
  assign tmp11060 = s4 ? tmp11045 : tmp11061;
  assign tmp11059 = s5 ? tmp11060 : tmp11048;
  assign tmp11058 = s6 ? tmp11041 : tmp11059;
  assign tmp11054 = s7 ? tmp11055 : tmp11058;
  assign tmp11067 = s3 ? tmp11002 : tmp9416;
  assign tmp11066 = s4 ? tmp11015 : tmp11067;
  assign tmp11065 = s5 ? tmp11066 : tmp11016;
  assign tmp11064 = s6 ? tmp11009 : tmp11065;
  assign tmp11053 = s8 ? tmp11054 : tmp11064;
  assign tmp11051 = s9 ? tmp11052 : tmp11053;
  assign tmp10966 = s10 ? tmp10967 : tmp11051;
  assign tmp11071 = s7 ? tmp10980 : tmp11040;
  assign tmp11070 = s8 ? tmp11071 : tmp11008;
  assign tmp11069 = s9 ? tmp11052 : tmp11070;
  assign tmp11068 = s10 ? tmp10967 : tmp11069;
  assign tmp10965 = s11 ? tmp10966 : tmp11068;
  assign tmp10915 = s12 ? tmp10916 : tmp10965;
  assign tmp11082 = s1 ? tmp9657 : tmp9618;
  assign tmp11081 = s2 ? tmp11082 : 1;
  assign tmp11080 = s3 ? tmp9680 : tmp11081;
  assign tmp11079 = s4 ? tmp9673 : tmp11080;
  assign tmp11085 = s2 ? tmp9689 : tmp10330;
  assign tmp11084 = s3 ? tmp11085 : tmp9623;
  assign tmp11087 = s2 ? tmp9172 : tmp10330;
  assign tmp11086 = s3 ? tmp11087 : tmp9482;
  assign tmp11083 = s4 ? tmp11084 : tmp11086;
  assign tmp11078 = s5 ? tmp11079 : tmp11083;
  assign tmp11077 = s6 ? tmp9654 : tmp11078;
  assign tmp11091 = s3 ? tmp9713 : tmp9502;
  assign tmp11090 = s4 ? tmp11091 : tmp9770;
  assign tmp11089 = s5 ? tmp9702 : tmp11090;
  assign tmp11088 = s6 ? tmp9697 : tmp11089;
  assign tmp11076 = s7 ? tmp11077 : tmp11088;
  assign tmp11097 = s2 ? tmp9383 : tmp10330;
  assign tmp11096 = s3 ? tmp11097 : tmp9482;
  assign tmp11095 = s4 ? tmp11084 : tmp11096;
  assign tmp11094 = s5 ? tmp9672 : tmp11095;
  assign tmp11093 = s6 ? tmp9654 : tmp11094;
  assign tmp11092 = s7 ? tmp11093 : tmp11088;
  assign tmp11075 = s8 ? tmp11076 : tmp11092;
  assign tmp11102 = s3 ? tmp9664 : tmp9858;
  assign tmp11101 = s4 ? tmp9655 : tmp11102;
  assign tmp11106 = s2 ? tmp9689 : tmp9657;
  assign tmp11105 = s3 ? tmp11106 : tmp9623;
  assign tmp11104 = s4 ? tmp11105 : tmp11096;
  assign tmp11103 = s5 ? tmp9672 : tmp11104;
  assign tmp11100 = s6 ? tmp11101 : tmp11103;
  assign tmp11109 = s3 ? tmp9699 : tmp9858;
  assign tmp11108 = s4 ? tmp9655 : tmp11109;
  assign tmp11112 = s3 ? tmp11106 : tmp9747;
  assign tmp11111 = s4 ? tmp11112 : tmp9770;
  assign tmp11110 = s5 ? tmp9702 : tmp11111;
  assign tmp11107 = s6 ? tmp11108 : tmp11110;
  assign tmp11099 = s7 ? tmp11100 : tmp11107;
  assign tmp11098 = s8 ? tmp11092 : tmp11099;
  assign tmp11074 = s9 ? tmp11075 : tmp11098;
  assign tmp11114 = s8 ? tmp11092 : tmp11093;
  assign tmp11116 = s7 ? tmp11088 : tmp11107;
  assign tmp11115 = s8 ? tmp11116 : tmp11088;
  assign tmp11113 = s9 ? tmp11114 : tmp11115;
  assign tmp11073 = s10 ? tmp11074 : tmp11113;
  assign tmp11125 = s3 ? tmp9757 : tmp9502;
  assign tmp11124 = s4 ? tmp11125 : tmp9766;
  assign tmp11123 = ~(s5 ? tmp9818 : tmp11124);
  assign tmp11122 = s6 ? tmp9813 : tmp11123;
  assign tmp11121 = s7 ? tmp9789 : tmp11122;
  assign tmp11128 = s5 ? tmp9860 : tmp11090;
  assign tmp11127 = s6 ? tmp9854 : tmp11128;
  assign tmp11126 = ~(s7 ? tmp9826 : tmp11127);
  assign tmp11120 = s8 ? tmp11121 : tmp11126;
  assign tmp11130 = s7 ? tmp9826 : tmp11127;
  assign tmp11129 = ~(s8 ? tmp11130 : tmp9867);
  assign tmp11119 = s9 ? tmp11120 : tmp11129;
  assign tmp11135 = ~(s5 ? tmp9875 : tmp11124);
  assign tmp11134 = s6 ? tmp9813 : tmp11135;
  assign tmp11133 = s7 ? tmp9868 : tmp11134;
  assign tmp11132 = s8 ? tmp11133 : tmp9868;
  assign tmp11140 = s4 ? tmp9879 : tmp9766;
  assign tmp11139 = ~(s5 ? tmp9875 : tmp11140);
  assign tmp11138 = s6 ? tmp9813 : tmp11139;
  assign tmp11137 = s7 ? tmp11122 : tmp11138;
  assign tmp11142 = ~(s6 ? tmp9813 : tmp11135);
  assign tmp11141 = ~(s7 ? tmp11127 : tmp11142);
  assign tmp11136 = s8 ? tmp11137 : tmp11141;
  assign tmp11131 = s9 ? tmp11132 : tmp11136;
  assign tmp11118 = s10 ? tmp11119 : tmp11131;
  assign tmp11146 = s7 ? tmp11122 : tmp9873;
  assign tmp11145 = s8 ? tmp11146 : tmp11141;
  assign tmp11144 = s9 ? tmp11132 : tmp11145;
  assign tmp11143 = s10 ? tmp11119 : tmp11144;
  assign tmp11117 = ~(s11 ? tmp11118 : tmp11143);
  assign tmp11072 = s12 ? tmp11073 : tmp11117;
  assign tmp10914 = ~(s13 ? tmp10915 : tmp11072);
  assign tmp10672 = s14 ? tmp10673 : tmp10914;
  assign tmp11160 = ~(s1 ? tmp9188 : tmp9615);
  assign tmp11159 = s2 ? tmp9801 : tmp11160;
  assign tmp11161 = ~(s2 ? tmp9224 : tmp10200);
  assign tmp11158 = s3 ? tmp11159 : tmp11161;
  assign tmp11157 = s4 ? tmp11158 : tmp10201;
  assign tmp11156 = s5 ? tmp11157 : tmp10206;
  assign tmp11155 = s6 ? tmp10277 : tmp11156;
  assign tmp11166 = s2 ? tmp9456 : tmp10057;
  assign tmp11165 = s3 ? tmp11166 : tmp9455;
  assign tmp11164 = s4 ? tmp11165 : tmp10223;
  assign tmp11168 = s3 ? tmp10075 : tmp10082;
  assign tmp11169 = s3 ? tmp10233 : tmp10077;
  assign tmp11167 = s4 ? tmp11168 : tmp11169;
  assign tmp11163 = s5 ? tmp11164 : tmp11167;
  assign tmp11162 = s6 ? tmp10282 : tmp11163;
  assign tmp11154 = s7 ? tmp11155 : tmp11162;
  assign tmp11174 = s2 ? tmp9744 : tmp10239;
  assign tmp11173 = s3 ? tmp9453 : tmp11174;
  assign tmp11172 = s4 ? tmp11173 : tmp10193;
  assign tmp11171 = s6 ? tmp11172 : tmp10240;
  assign tmp11176 = s4 ? tmp11173 : tmp10258;
  assign tmp11179 = s3 ? tmp10270 : tmp10082;
  assign tmp11181 = s2 ? tmp10009 : tmp9172;
  assign tmp11180 = s3 ? tmp11181 : tmp10077;
  assign tmp11178 = s4 ? tmp11179 : tmp11180;
  assign tmp11177 = s5 ? tmp10261 : tmp11178;
  assign tmp11175 = s6 ? tmp11176 : tmp11177;
  assign tmp11170 = s7 ? tmp11171 : tmp11175;
  assign tmp11153 = s8 ? tmp11154 : tmp11170;
  assign tmp11188 = s2 ? tmp9801 : tmp10245;
  assign tmp11189 = s2 ? tmp9174 : tmp9456;
  assign tmp11187 = s3 ? tmp11188 : tmp11189;
  assign tmp11186 = s4 ? tmp11187 : tmp10201;
  assign tmp11185 = s5 ? tmp11186 : tmp10206;
  assign tmp11184 = s6 ? tmp10277 : tmp11185;
  assign tmp11194 = s2 ? tmp9456 : tmp9636;
  assign tmp11193 = s3 ? tmp11194 : tmp9455;
  assign tmp11192 = s4 ? tmp11193 : tmp10266;
  assign tmp11191 = s5 ? tmp11192 : tmp10286;
  assign tmp11190 = s6 ? tmp10282 : tmp11191;
  assign tmp11183 = s7 ? tmp11184 : tmp11190;
  assign tmp11182 = s8 ? tmp11170 : tmp11183;
  assign tmp11152 = s9 ? tmp11153 : tmp11182;
  assign tmp11199 = s5 ? tmp11192 : tmp11167;
  assign tmp11198 = s6 ? tmp10282 : tmp11199;
  assign tmp11197 = s7 ? tmp11184 : tmp11198;
  assign tmp11196 = s8 ? tmp11197 : tmp11184;
  assign tmp11204 = s4 ? tmp11165 : tmp10301;
  assign tmp11203 = s5 ? tmp11204 : tmp11167;
  assign tmp11202 = s6 ? tmp10282 : tmp11203;
  assign tmp11206 = s5 ? tmp11192 : tmp10306;
  assign tmp11205 = s6 ? tmp10282 : tmp11206;
  assign tmp11201 = s7 ? tmp11202 : tmp11205;
  assign tmp11207 = s7 ? tmp11175 : tmp11198;
  assign tmp11200 = s8 ? tmp11201 : tmp11207;
  assign tmp11195 = s9 ? tmp11196 : tmp11200;
  assign tmp11151 = s10 ? tmp11152 : tmp11195;
  assign tmp11211 = s7 ? tmp11162 : tmp11190;
  assign tmp11210 = s8 ? tmp11211 : tmp11207;
  assign tmp11209 = s9 ? tmp11196 : tmp11210;
  assign tmp11208 = s10 ? tmp11152 : tmp11209;
  assign tmp11150 = s11 ? tmp11151 : tmp11208;
  assign tmp11219 = s3 ? tmp10328 : tmp9660;
  assign tmp11218 = s4 ? tmp11219 : tmp10331;
  assign tmp11223 = s2 ? tmp9838 : tmp9657;
  assign tmp11222 = s3 ? tmp11223 : tmp10347;
  assign tmp11221 = s4 ? tmp11222 : tmp10349;
  assign tmp11220 = s5 ? tmp10335 : tmp11221;
  assign tmp11217 = s6 ? tmp11218 : tmp11220;
  assign tmp11225 = s4 ? tmp11219 : tmp10358;
  assign tmp11229 = s2 ? tmp9830 : tmp10997;
  assign tmp11228 = s3 ? tmp11229 : tmp10371;
  assign tmp11227 = s4 ? tmp11228 : tmp9657;
  assign tmp11226 = s5 ? tmp10361 : tmp11227;
  assign tmp11224 = s6 ? tmp11225 : tmp11226;
  assign tmp11216 = s7 ? tmp11217 : tmp11224;
  assign tmp11215 = s8 ? tmp10324 : tmp11216;
  assign tmp11214 = s9 ? tmp10324 : tmp11215;
  assign tmp11233 = s6 ? tmp11218 : tmp10334;
  assign tmp11234 = s6 ? tmp11225 : tmp10360;
  assign tmp11232 = s7 ? tmp11233 : tmp11234;
  assign tmp11231 = s8 ? tmp11232 : tmp11233;
  assign tmp11236 = s7 ? tmp10403 : tmp11224;
  assign tmp11237 = s6 ? tmp11225 : tmp10404;
  assign tmp11235 = s8 ? tmp11236 : tmp11237;
  assign tmp11230 = s9 ? tmp11231 : tmp11235;
  assign tmp11213 = s10 ? tmp11214 : tmp11230;
  assign tmp11241 = s7 ? tmp10356 : tmp11224;
  assign tmp11240 = s8 ? tmp11241 : tmp11234;
  assign tmp11239 = s9 ? tmp11231 : tmp11240;
  assign tmp11238 = s10 ? tmp11214 : tmp11239;
  assign tmp11212 = s11 ? tmp11213 : tmp11238;
  assign tmp11149 = s12 ? tmp11150 : tmp11212;
  assign tmp11148 = s13 ? tmp11149 : tmp10411;
  assign tmp11147 = ~(s14 ? tmp9899 : tmp11148);
  assign tmp10671 = s15 ? tmp10672 : tmp11147;
  assign tmp9135 = s16 ? tmp9136 : tmp10671;
  assign tmp11253 = s4 ? tmp10733 : tmp9283;
  assign tmp11252 = s5 ? tmp9250 : tmp11253;
  assign tmp11251 = s6 ? tmp9243 : tmp11252;
  assign tmp11256 = s4 ? tmp10752 : tmp9283;
  assign tmp11255 = s5 ? tmp9273 : tmp11256;
  assign tmp11254 = s6 ? tmp9243 : tmp11255;
  assign tmp11250 = s7 ? tmp11251 : tmp11254;
  assign tmp11249 = s8 ? tmp10688 : tmp11250;
  assign tmp11248 = s9 ? tmp10677 : tmp11249;
  assign tmp11261 = s5 ? tmp9290 : tmp10686;
  assign tmp11260 = s6 ? tmp9193 : tmp11261;
  assign tmp11259 = s7 ? tmp10679 : tmp11260;
  assign tmp11258 = s8 ? tmp11259 : tmp10679;
  assign tmp11263 = s7 ? tmp10798 : tmp11254;
  assign tmp11264 = s7 ? tmp10802 : tmp11260;
  assign tmp11262 = s8 ? tmp11263 : tmp11264;
  assign tmp11257 = s9 ? tmp11258 : tmp11262;
  assign tmp11247 = s10 ? tmp11248 : tmp11257;
  assign tmp11268 = s7 ? tmp10684 : tmp11254;
  assign tmp11269 = s7 ? tmp10699 : tmp11260;
  assign tmp11267 = s8 ? tmp11268 : tmp11269;
  assign tmp11266 = s9 ? tmp11258 : tmp11267;
  assign tmp11265 = s10 ? tmp11248 : tmp11266;
  assign tmp11246 = s11 ? tmp11247 : tmp11265;
  assign tmp11275 = s7 ? tmp10826 : tmp10895;
  assign tmp11274 = s8 ? tmp10846 : tmp11275;
  assign tmp11273 = s9 ? tmp10824 : tmp11274;
  assign tmp11277 = s8 ? tmp11275 : tmp10826;
  assign tmp11279 = s7 ? tmp10905 : tmp10895;
  assign tmp11278 = s8 ? tmp10895 : tmp11279;
  assign tmp11276 = s9 ? tmp11277 : tmp11278;
  assign tmp11272 = s10 ? tmp11273 : tmp11276;
  assign tmp11283 = s7 ? tmp10839 : tmp10895;
  assign tmp11284 = s7 ? tmp10855 : tmp10895;
  assign tmp11282 = s8 ? tmp11283 : tmp11284;
  assign tmp11281 = s9 ? tmp11277 : tmp11282;
  assign tmp11280 = s10 ? tmp11273 : tmp11281;
  assign tmp11271 = s11 ? tmp11272 : tmp11280;
  assign tmp11270 = s12 ? tmp9306 : tmp11271;
  assign tmp11245 = s13 ? tmp11246 : tmp11270;
  assign tmp11290 = s8 ? tmp10920 : tmp9426;
  assign tmp11289 = s9 ? tmp10919 : tmp11290;
  assign tmp11293 = s7 ? tmp10956 : tmp9417;
  assign tmp11292 = s8 ? tmp9437 : tmp11293;
  assign tmp11291 = s9 ? tmp9435 : tmp11292;
  assign tmp11288 = s10 ? tmp11289 : tmp11291;
  assign tmp11297 = s7 ? tmp10939 : tmp9417;
  assign tmp11296 = s8 ? tmp9417 : tmp11297;
  assign tmp11295 = s9 ? tmp9435 : tmp11296;
  assign tmp11294 = s10 ? tmp11289 : tmp11295;
  assign tmp11287 = s11 ? tmp11288 : tmp11294;
  assign tmp11307 = s1 ? tmp9254 : tmp9151;
  assign tmp11306 = s2 ? tmp9151 : tmp11307;
  assign tmp11305 = s3 ? tmp9151 : tmp11306;
  assign tmp11309 = s2 ? tmp9151 : tmp9254;
  assign tmp11308 = s3 ? tmp11309 : tmp9557;
  assign tmp11304 = s4 ? tmp11305 : tmp11308;
  assign tmp11314 = s1 ? tmp9254 : tmp9350;
  assign tmp11315 = ~(s1 ? tmp9256 : tmp9326);
  assign tmp11313 = s2 ? tmp11314 : tmp11315;
  assign tmp11316 = ~(s2 ? tmp9256 : tmp9566);
  assign tmp11312 = s3 ? tmp11313 : tmp11316;
  assign tmp11311 = s4 ? tmp11312 : tmp9537;
  assign tmp11310 = s5 ? tmp11311 : tmp9541;
  assign tmp11303 = s6 ? tmp11304 : tmp11310;
  assign tmp11319 = s3 ? tmp11306 : tmp9557;
  assign tmp11318 = s4 ? tmp11305 : tmp11319;
  assign tmp11324 = s1 ? tmp9254 : 1;
  assign tmp11323 = s2 ? tmp11324 : tmp9253;
  assign tmp11322 = s3 ? tmp11323 : tmp9535;
  assign tmp11321 = s4 ? tmp11322 : tmp9537;
  assign tmp11320 = s5 ? tmp11321 : tmp9562;
  assign tmp11317 = s6 ? tmp11318 : tmp11320;
  assign tmp11302 = ~(s7 ? tmp11303 : tmp11317);
  assign tmp11301 = s8 ? tmp10989 : tmp11302;
  assign tmp11300 = s9 ? tmp10968 : tmp11301;
  assign tmp11330 = s4 ? tmp10986 : tmp9520;
  assign tmp11329 = s5 ? tmp11330 : tmp9499;
  assign tmp11328 = s6 ? tmp10981 : tmp11329;
  assign tmp11327 = s7 ? tmp10970 : tmp11328;
  assign tmp11326 = s8 ? tmp11327 : tmp10970;
  assign tmp11333 = ~(s6 ? tmp11318 : tmp11320);
  assign tmp11332 = s7 ? tmp11055 : tmp11333;
  assign tmp11334 = s7 ? tmp11064 : tmp11328;
  assign tmp11331 = s8 ? tmp11332 : tmp11334;
  assign tmp11325 = s9 ? tmp11326 : tmp11331;
  assign tmp11299 = s10 ? tmp11300 : tmp11325;
  assign tmp11338 = s7 ? tmp10980 : tmp11333;
  assign tmp11339 = s7 ? tmp11008 : tmp11328;
  assign tmp11337 = s8 ? tmp11338 : tmp11339;
  assign tmp11336 = s9 ? tmp11326 : tmp11337;
  assign tmp11335 = s10 ? tmp11300 : tmp11336;
  assign tmp11298 = s11 ? tmp11299 : tmp11335;
  assign tmp11286 = s12 ? tmp11287 : tmp11298;
  assign tmp11351 = s1 ? tmp10212 : tmp9343;
  assign tmp11350 = s2 ? tmp11351 : tmp9614;
  assign tmp11349 = s3 ? tmp11350 : tmp9616;
  assign tmp11348 = s4 ? tmp9603 : tmp11349;
  assign tmp11347 = s5 ? tmp11348 : tmp9619;
  assign tmp11346 = s6 ? tmp9594 : tmp11347;
  assign tmp11356 = s2 ? tmp11351 : tmp9172;
  assign tmp11355 = s3 ? tmp11356 : tmp9640;
  assign tmp11354 = s4 ? tmp9634 : tmp11355;
  assign tmp11353 = s5 ? tmp11354 : tmp9642;
  assign tmp11352 = s6 ? tmp9628 : tmp11353;
  assign tmp11345 = s7 ? tmp11346 : tmp11352;
  assign tmp11363 = s1 ? tmp10212 : tmp9257;
  assign tmp11364 = ~(s1 ? tmp9151 : tmp9615);
  assign tmp11362 = s2 ? tmp11363 : tmp11364;
  assign tmp11361 = s3 ? tmp11362 : tmp9471;
  assign tmp11360 = s4 ? tmp11000 : tmp11361;
  assign tmp11368 = s1 ? tmp9174 : tmp9622;
  assign tmp11367 = s2 ? tmp9475 : tmp11368;
  assign tmp11366 = s3 ? tmp11367 : tmp9623;
  assign tmp11370 = s2 ? tmp9383 : tmp9626;
  assign tmp11369 = s3 ? tmp11370 : tmp9482;
  assign tmp11365 = s4 ? tmp11366 : tmp11369;
  assign tmp11359 = s5 ? tmp11360 : tmp11365;
  assign tmp11358 = s6 ? tmp9594 : tmp11359;
  assign tmp11375 = s2 ? tmp11363 : tmp9172;
  assign tmp11374 = s3 ? tmp11375 : tmp9416;
  assign tmp11373 = s4 ? tmp11015 : tmp11374;
  assign tmp11372 = s5 ? tmp11373 : tmp9642;
  assign tmp11371 = s6 ? tmp9628 : tmp11372;
  assign tmp11357 = s7 ? tmp11358 : tmp11371;
  assign tmp11344 = s8 ? tmp11345 : tmp11357;
  assign tmp11384 = s0 ? tmp9151 : tmp9657;
  assign tmp11383 = s1 ? tmp11384 : tmp9343;
  assign tmp11382 = s2 ? tmp11383 : tmp9728;
  assign tmp11381 = s3 ? tmp11382 : tmp9729;
  assign tmp11380 = s4 ? tmp9722 : tmp11381;
  assign tmp11379 = s5 ? tmp11380 : tmp9731;
  assign tmp11378 = s6 ? tmp9654 : tmp11379;
  assign tmp11389 = s2 ? tmp11383 : tmp9657;
  assign tmp11388 = s3 ? tmp11389 : tmp9743;
  assign tmp11387 = s4 ? tmp9739 : tmp11388;
  assign tmp11386 = s5 ? tmp11387 : tmp9745;
  assign tmp11385 = s6 ? tmp9697 : tmp11386;
  assign tmp11377 = s7 ? tmp11378 : tmp11385;
  assign tmp11376 = s8 ? tmp11357 : tmp11377;
  assign tmp11343 = s9 ? tmp11344 : tmp11376;
  assign tmp11394 = s5 ? tmp11354 : tmp9755;
  assign tmp11393 = s6 ? tmp9628 : tmp11394;
  assign tmp11392 = s7 ? tmp11346 : tmp11393;
  assign tmp11391 = s8 ? tmp11392 : tmp11346;
  assign tmp11398 = s5 ? tmp11354 : tmp9765;
  assign tmp11397 = s6 ? tmp9628 : tmp11398;
  assign tmp11400 = s5 ? tmp11387 : tmp9769;
  assign tmp11399 = s6 ? tmp9697 : tmp11400;
  assign tmp11396 = s7 ? tmp11397 : tmp11399;
  assign tmp11403 = s5 ? tmp11373 : tmp9765;
  assign tmp11402 = s6 ? tmp9628 : tmp11403;
  assign tmp11405 = s5 ? tmp11354 : tmp9778;
  assign tmp11404 = s6 ? tmp9628 : tmp11405;
  assign tmp11401 = s7 ? tmp11402 : tmp11404;
  assign tmp11395 = s8 ? tmp11396 : tmp11401;
  assign tmp11390 = s9 ? tmp11391 : tmp11395;
  assign tmp11342 = s10 ? tmp11343 : tmp11390;
  assign tmp11409 = s7 ? tmp11352 : tmp11385;
  assign tmp11410 = s7 ? tmp11371 : tmp11393;
  assign tmp11408 = s8 ? tmp11409 : tmp11410;
  assign tmp11407 = s9 ? tmp11391 : tmp11408;
  assign tmp11406 = s10 ? tmp11343 : tmp11407;
  assign tmp11341 = s11 ? tmp11342 : tmp11406;
  assign tmp11340 = s12 ? tmp11341 : tmp9784;
  assign tmp11285 = ~(s13 ? tmp11286 : tmp11340);
  assign tmp11244 = s14 ? tmp11245 : tmp11285;
  assign tmp11417 = s8 ? tmp10324 : tmp10390;
  assign tmp11416 = s9 ? tmp10324 : tmp11417;
  assign tmp11420 = s7 ? tmp10403 : tmp10397;
  assign tmp11419 = s8 ? tmp10402 : tmp11420;
  assign tmp11418 = s9 ? tmp10395 : tmp11419;
  assign tmp11415 = s10 ? tmp11416 : tmp11418;
  assign tmp11424 = s7 ? tmp10356 : tmp10397;
  assign tmp11423 = s8 ? tmp10410 : tmp11424;
  assign tmp11422 = s9 ? tmp10395 : tmp11423;
  assign tmp11421 = s10 ? tmp11416 : tmp11422;
  assign tmp11414 = s11 ? tmp11415 : tmp11421;
  assign tmp11413 = s12 ? tmp10183 : tmp11414;
  assign tmp11412 = s13 ? tmp11413 : tmp10411;
  assign tmp11411 = ~(s14 ? tmp9899 : tmp11412);
  assign tmp11243 = s15 ? tmp11244 : tmp11411;
  assign tmp11439 = s1 ? tmp11384 : tmp9257;
  assign tmp11438 = s2 ? tmp11439 : tmp9682;
  assign tmp11437 = s3 ? tmp11438 : tmp9684;
  assign tmp11436 = s4 ? tmp9673 : tmp11437;
  assign tmp11435 = s5 ? tmp11436 : tmp9686;
  assign tmp11434 = s6 ? tmp9654 : tmp11435;
  assign tmp11444 = s2 ? tmp11439 : tmp9657;
  assign tmp11443 = s3 ? tmp11444 : tmp9709;
  assign tmp11442 = s4 ? tmp9703 : tmp11443;
  assign tmp11446 = s3 ? tmp9851 : tmp9747;
  assign tmp11449 = s1 ? tmp9657 : tmp9695;
  assign tmp11448 = s2 ? 1 : tmp11449;
  assign tmp11447 = s3 ? tmp11448 : tmp9172;
  assign tmp11445 = s4 ? tmp11446 : tmp11447;
  assign tmp11441 = s5 ? tmp11442 : tmp11445;
  assign tmp11440 = s6 ? tmp9697 : tmp11441;
  assign tmp11433 = s7 ? tmp11434 : tmp11440;
  assign tmp11432 = s8 ? tmp11357 : tmp11433;
  assign tmp11431 = s9 ? tmp11344 : tmp11432;
  assign tmp11451 = s8 ? tmp11357 : tmp11358;
  assign tmp11456 = s4 ? tmp11446 : tmp9770;
  assign tmp11455 = s5 ? tmp11442 : tmp11456;
  assign tmp11454 = s6 ? tmp9697 : tmp11455;
  assign tmp11453 = s7 ? tmp11397 : tmp11454;
  assign tmp11452 = s8 ? tmp11453 : tmp11402;
  assign tmp11450 = s9 ? tmp11451 : tmp11452;
  assign tmp11430 = s10 ? tmp11431 : tmp11450;
  assign tmp11460 = s7 ? tmp11352 : tmp11440;
  assign tmp11459 = s8 ? tmp11460 : tmp11371;
  assign tmp11458 = s9 ? tmp11451 : tmp11459;
  assign tmp11457 = s10 ? tmp11431 : tmp11458;
  assign tmp11429 = s11 ? tmp11430 : tmp11457;
  assign tmp11428 = s12 ? tmp11429 : tmp9784;
  assign tmp11427 = ~(s13 ? tmp10915 : tmp11428);
  assign tmp11426 = s14 ? tmp10673 : tmp11427;
  assign tmp11463 = s12 ? tmp10183 : tmp11212;
  assign tmp11462 = s13 ? tmp11463 : tmp10411;
  assign tmp11461 = ~(s14 ? tmp9899 : tmp11462);
  assign tmp11425 = s15 ? tmp11426 : tmp11461;
  assign tmp11242 = s16 ? tmp11243 : tmp11425;
  assign tmp9134 = ~(s17 ? tmp9135 : tmp11242);
  assign l2__1 = tmp9134;

  assign tmp11479 = l3 ? 1 : 0;
  assign tmp11480 = l2 ? 1 : 0;
  assign tmp11478 = l1 ? tmp11479 : tmp11480;
  assign tmp11482 = l1 ? tmp11479 : 1;
  assign tmp11481 = s0 ? tmp11482 : tmp11478;
  assign tmp11477 = s1 ? tmp11478 : tmp11481;
  assign tmp11485 = s0 ? tmp11478 : 1;
  assign tmp11484 = s1 ? tmp11485 : tmp11478;
  assign tmp11483 = s2 ? tmp11478 : tmp11484;
  assign tmp11476 = s3 ? tmp11477 : tmp11483;
  assign tmp11489 = s0 ? tmp11478 : tmp11482;
  assign tmp11488 = s1 ? tmp11489 : tmp11478;
  assign tmp11491 = s0 ? tmp11482 : 1;
  assign tmp11490 = s1 ? tmp11485 : tmp11491;
  assign tmp11487 = s2 ? tmp11488 : tmp11490;
  assign tmp11494 = s0 ? 1 : 0;
  assign tmp11493 = s1 ? tmp11482 : tmp11494;
  assign tmp11496 = s0 ? tmp11478 : tmp11480;
  assign tmp11498 = ~(l1 ? tmp11479 : tmp11480);
  assign tmp11497 = ~(s0 ? 1 : tmp11498);
  assign tmp11495 = s1 ? tmp11496 : tmp11497;
  assign tmp11492 = s2 ? tmp11493 : tmp11495;
  assign tmp11486 = s3 ? tmp11487 : tmp11492;
  assign tmp11475 = s4 ? tmp11476 : tmp11486;
  assign tmp11504 = s0 ? 1 : tmp11478;
  assign tmp11503 = s1 ? tmp11485 : tmp11504;
  assign tmp11506 = s0 ? tmp11480 : 1;
  assign tmp11505 = s1 ? tmp11504 : tmp11506;
  assign tmp11502 = s2 ? tmp11503 : tmp11505;
  assign tmp11508 = s0 ? 1 : tmp11480;
  assign tmp11510 = ~(s0 ? tmp11478 : 0);
  assign tmp11509 = ~(s1 ? 1 : tmp11510);
  assign tmp11507 = s2 ? tmp11508 : tmp11509;
  assign tmp11501 = s3 ? tmp11502 : tmp11507;
  assign tmp11514 = s0 ? 1 : tmp11498;
  assign tmp11515 = ~(s0 ? tmp11482 : 0);
  assign tmp11513 = s1 ? tmp11514 : tmp11515;
  assign tmp11517 = s0 ? tmp11482 : 0;
  assign tmp11516 = ~(s1 ? tmp11517 : tmp11489);
  assign tmp11512 = s2 ? tmp11513 : tmp11516;
  assign tmp11519 = s1 ? tmp11480 : 0;
  assign tmp11518 = ~(s2 ? tmp11519 : 0);
  assign tmp11511 = ~(s3 ? tmp11512 : tmp11518);
  assign tmp11500 = s4 ? tmp11501 : tmp11511;
  assign tmp11524 = s0 ? tmp11480 : 0;
  assign tmp11523 = s1 ? tmp11524 : 0;
  assign tmp11527 = ~(l2 ? 1 : 0);
  assign tmp11526 = s0 ? 1 : tmp11527;
  assign tmp11525 = ~(s1 ? tmp11526 : tmp11527);
  assign tmp11522 = s2 ? tmp11523 : tmp11525;
  assign tmp11521 = s3 ? tmp11522 : 0;
  assign tmp11530 = s1 ? tmp11526 : tmp11527;
  assign tmp11529 = s2 ? 1 : tmp11530;
  assign tmp11528 = ~(s3 ? tmp11529 : 1);
  assign tmp11520 = s4 ? tmp11521 : tmp11528;
  assign tmp11499 = s5 ? tmp11500 : tmp11520;
  assign tmp11474 = s6 ? tmp11475 : tmp11499;
  assign tmp11535 = s1 ? tmp11485 : tmp11482;
  assign tmp11534 = s2 ? tmp11488 : tmp11535;
  assign tmp11537 = s1 ? tmp11482 : 0;
  assign tmp11536 = s2 ? tmp11537 : tmp11495;
  assign tmp11533 = s3 ? tmp11534 : tmp11536;
  assign tmp11532 = s4 ? tmp11476 : tmp11533;
  assign tmp11542 = s1 ? tmp11478 : tmp11506;
  assign tmp11541 = s2 ? tmp11484 : tmp11542;
  assign tmp11543 = s2 ? tmp11480 : tmp11509;
  assign tmp11540 = s3 ? tmp11541 : tmp11543;
  assign tmp11546 = ~(s1 ? tmp11482 : tmp11489);
  assign tmp11545 = s2 ? tmp11513 : tmp11546;
  assign tmp11544 = ~(s3 ? tmp11545 : tmp11518);
  assign tmp11539 = s4 ? tmp11540 : tmp11544;
  assign tmp11549 = s2 ? tmp11523 : tmp11519;
  assign tmp11548 = s3 ? tmp11549 : 0;
  assign tmp11551 = s2 ? 1 : tmp11527;
  assign tmp11550 = ~(s3 ? tmp11551 : 1);
  assign tmp11547 = s4 ? tmp11548 : tmp11550;
  assign tmp11538 = s5 ? tmp11539 : tmp11547;
  assign tmp11531 = s6 ? tmp11532 : tmp11538;
  assign tmp11473 = s7 ? tmp11474 : tmp11531;
  assign tmp11558 = l2 ? 1 : tmp11479;
  assign tmp11557 = l1 ? tmp11558 : tmp11480;
  assign tmp11560 = l1 ? tmp11558 : 1;
  assign tmp11559 = s0 ? tmp11560 : tmp11557;
  assign tmp11556 = s1 ? tmp11557 : tmp11559;
  assign tmp11563 = s0 ? tmp11557 : 1;
  assign tmp11562 = s1 ? tmp11563 : tmp11557;
  assign tmp11561 = s2 ? tmp11557 : tmp11562;
  assign tmp11555 = s3 ? tmp11556 : tmp11561;
  assign tmp11567 = s0 ? tmp11557 : tmp11560;
  assign tmp11566 = s1 ? tmp11567 : tmp11557;
  assign tmp11569 = s0 ? tmp11560 : 1;
  assign tmp11568 = s1 ? tmp11563 : tmp11569;
  assign tmp11565 = s2 ? tmp11566 : tmp11568;
  assign tmp11571 = s1 ? tmp11560 : tmp11494;
  assign tmp11573 = s0 ? tmp11557 : tmp11480;
  assign tmp11575 = ~(l1 ? tmp11558 : tmp11480);
  assign tmp11574 = ~(s0 ? 1 : tmp11575);
  assign tmp11572 = s1 ? tmp11573 : tmp11574;
  assign tmp11570 = s2 ? tmp11571 : tmp11572;
  assign tmp11564 = s3 ? tmp11565 : tmp11570;
  assign tmp11554 = s4 ? tmp11555 : tmp11564;
  assign tmp11581 = s0 ? 1 : tmp11557;
  assign tmp11580 = s1 ? tmp11563 : tmp11581;
  assign tmp11582 = s1 ? tmp11581 : tmp11506;
  assign tmp11579 = s2 ? tmp11580 : tmp11582;
  assign tmp11586 = l1 ? tmp11480 : 0;
  assign tmp11585 = ~(s0 ? tmp11557 : tmp11586);
  assign tmp11584 = ~(s1 ? 1 : tmp11585);
  assign tmp11583 = s2 ? tmp11508 : tmp11584;
  assign tmp11578 = s3 ? tmp11579 : tmp11583;
  assign tmp11590 = s0 ? 1 : tmp11575;
  assign tmp11591 = ~(s0 ? tmp11560 : tmp11480);
  assign tmp11589 = s1 ? tmp11590 : tmp11591;
  assign tmp11593 = s0 ? tmp11560 : tmp11480;
  assign tmp11592 = ~(s1 ? tmp11593 : tmp11567);
  assign tmp11588 = s2 ? tmp11589 : tmp11592;
  assign tmp11596 = s0 ? tmp11480 : tmp11586;
  assign tmp11595 = s1 ? tmp11596 : tmp11524;
  assign tmp11594 = ~(s2 ? tmp11595 : 0);
  assign tmp11587 = ~(s3 ? tmp11588 : tmp11594);
  assign tmp11577 = s4 ? tmp11578 : tmp11587;
  assign tmp11576 = s5 ? tmp11577 : tmp11520;
  assign tmp11553 = s6 ? tmp11554 : tmp11576;
  assign tmp11601 = s1 ? tmp11563 : tmp11560;
  assign tmp11600 = s2 ? tmp11566 : tmp11601;
  assign tmp11603 = s1 ? tmp11560 : 0;
  assign tmp11602 = s2 ? tmp11603 : tmp11572;
  assign tmp11599 = s3 ? tmp11600 : tmp11602;
  assign tmp11598 = s4 ? tmp11555 : tmp11599;
  assign tmp11608 = s1 ? tmp11557 : tmp11506;
  assign tmp11607 = s2 ? tmp11562 : tmp11608;
  assign tmp11609 = s2 ? tmp11480 : tmp11584;
  assign tmp11606 = s3 ? tmp11607 : tmp11609;
  assign tmp11611 = s2 ? tmp11589 : tmp11575;
  assign tmp11613 = s1 ? tmp11596 : 0;
  assign tmp11612 = ~(s2 ? tmp11613 : 0);
  assign tmp11610 = ~(s3 ? tmp11611 : tmp11612);
  assign tmp11605 = s4 ? tmp11606 : tmp11610;
  assign tmp11604 = s5 ? tmp11605 : tmp11547;
  assign tmp11597 = s6 ? tmp11598 : tmp11604;
  assign tmp11552 = s7 ? tmp11553 : tmp11597;
  assign tmp11472 = s8 ? tmp11473 : tmp11552;
  assign tmp11619 = s2 ? tmp11482 : tmp11491;
  assign tmp11623 = ~(l1 ? 1 : 0);
  assign tmp11622 = s0 ? tmp11482 : tmp11623;
  assign tmp11625 = ~(l1 ? tmp11479 : 1);
  assign tmp11624 = ~(s0 ? 1 : tmp11625);
  assign tmp11621 = s1 ? tmp11622 : tmp11624;
  assign tmp11620 = s2 ? tmp11493 : tmp11621;
  assign tmp11618 = s3 ? tmp11619 : tmp11620;
  assign tmp11617 = s4 ? tmp11482 : tmp11618;
  assign tmp11632 = l1 ? 1 : 0;
  assign tmp11631 = ~(s0 ? tmp11632 : 0);
  assign tmp11630 = s1 ? tmp11482 : tmp11631;
  assign tmp11629 = s2 ? tmp11482 : tmp11630;
  assign tmp11634 = s0 ? 1 : tmp11623;
  assign tmp11635 = ~(s1 ? 1 : tmp11515);
  assign tmp11633 = s2 ? tmp11634 : tmp11635;
  assign tmp11628 = s3 ? tmp11629 : tmp11633;
  assign tmp11639 = s0 ? 1 : tmp11625;
  assign tmp11638 = s1 ? tmp11639 : tmp11515;
  assign tmp11640 = ~(s1 ? tmp11517 : tmp11482);
  assign tmp11637 = s2 ? tmp11638 : tmp11640;
  assign tmp11641 = s2 ? tmp11632 : 1;
  assign tmp11636 = ~(s3 ? tmp11637 : tmp11641);
  assign tmp11627 = s4 ? tmp11628 : tmp11636;
  assign tmp11646 = s0 ? tmp11632 : 1;
  assign tmp11645 = s1 ? tmp11646 : 1;
  assign tmp11648 = s0 ? 1 : tmp11632;
  assign tmp11647 = s1 ? tmp11648 : tmp11632;
  assign tmp11644 = s2 ? tmp11645 : tmp11647;
  assign tmp11643 = s3 ? tmp11644 : 1;
  assign tmp11650 = s2 ? 1 : tmp11647;
  assign tmp11649 = s3 ? tmp11650 : 1;
  assign tmp11642 = ~(s4 ? tmp11643 : tmp11649);
  assign tmp11626 = s5 ? tmp11627 : tmp11642;
  assign tmp11616 = s6 ? tmp11617 : tmp11626;
  assign tmp11655 = s1 ? tmp11491 : tmp11482;
  assign tmp11654 = s2 ? tmp11482 : tmp11655;
  assign tmp11656 = s2 ? tmp11537 : tmp11621;
  assign tmp11653 = s3 ? tmp11654 : tmp11656;
  assign tmp11652 = s4 ? tmp11482 : tmp11653;
  assign tmp11661 = s1 ? 1 : tmp11515;
  assign tmp11660 = ~(s2 ? tmp11632 : tmp11661);
  assign tmp11659 = s3 ? tmp11629 : tmp11660;
  assign tmp11663 = s2 ? tmp11638 : tmp11625;
  assign tmp11665 = s1 ? tmp11632 : 1;
  assign tmp11664 = s2 ? tmp11665 : 1;
  assign tmp11662 = ~(s3 ? tmp11663 : tmp11664);
  assign tmp11658 = s4 ? tmp11659 : tmp11662;
  assign tmp11668 = s2 ? tmp11645 : tmp11665;
  assign tmp11667 = s3 ? tmp11668 : 1;
  assign tmp11670 = s2 ? 1 : tmp11632;
  assign tmp11669 = s3 ? tmp11670 : 1;
  assign tmp11666 = ~(s4 ? tmp11667 : tmp11669);
  assign tmp11657 = s5 ? tmp11658 : tmp11666;
  assign tmp11651 = s6 ? tmp11652 : tmp11657;
  assign tmp11615 = s7 ? tmp11616 : tmp11651;
  assign tmp11614 = s8 ? tmp11552 : tmp11615;
  assign tmp11471 = s9 ? tmp11472 : tmp11614;
  assign tmp11678 = s2 ? tmp11513 : tmp11498;
  assign tmp11677 = ~(s3 ? tmp11678 : tmp11518);
  assign tmp11676 = s4 ? tmp11540 : tmp11677;
  assign tmp11675 = s5 ? tmp11676 : tmp11547;
  assign tmp11674 = s6 ? tmp11532 : tmp11675;
  assign tmp11673 = s7 ? tmp11474 : tmp11674;
  assign tmp11672 = s8 ? tmp11673 : tmp11474;
  assign tmp11686 = ~(s1 ? tmp11482 : tmp11478);
  assign tmp11685 = s2 ? tmp11513 : tmp11686;
  assign tmp11684 = ~(s3 ? tmp11685 : tmp11518);
  assign tmp11683 = s4 ? tmp11540 : tmp11684;
  assign tmp11682 = s5 ? tmp11683 : tmp11547;
  assign tmp11681 = s6 ? tmp11532 : tmp11682;
  assign tmp11680 = s7 ? tmp11681 : tmp11651;
  assign tmp11687 = s7 ? tmp11597 : tmp11674;
  assign tmp11679 = s8 ? tmp11680 : tmp11687;
  assign tmp11671 = s9 ? tmp11672 : tmp11679;
  assign tmp11470 = s10 ? tmp11471 : tmp11671;
  assign tmp11691 = s7 ? tmp11531 : tmp11651;
  assign tmp11690 = s8 ? tmp11691 : tmp11687;
  assign tmp11689 = s9 ? tmp11672 : tmp11690;
  assign tmp11688 = s10 ? tmp11471 : tmp11689;
  assign tmp11469 = s11 ? tmp11470 : tmp11688;
  assign tmp11468 = s13 ? tmp11469 : 1;
  assign tmp11693 = s12 ? 1 : 0;
  assign tmp11704 = l1 ? 1 : tmp11527;
  assign tmp11705 = s0 ? tmp11632 : tmp11704;
  assign tmp11703 = s1 ? tmp11704 : tmp11705;
  assign tmp11708 = s0 ? tmp11704 : 0;
  assign tmp11707 = s1 ? tmp11708 : tmp11704;
  assign tmp11706 = s2 ? tmp11704 : tmp11707;
  assign tmp11702 = s3 ? tmp11703 : tmp11706;
  assign tmp11712 = s0 ? tmp11704 : tmp11632;
  assign tmp11711 = s1 ? tmp11712 : tmp11704;
  assign tmp11714 = s0 ? tmp11632 : 0;
  assign tmp11713 = s1 ? tmp11708 : tmp11714;
  assign tmp11710 = s2 ? tmp11711 : tmp11713;
  assign tmp11717 = ~(s0 ? 1 : 0);
  assign tmp11716 = s1 ? tmp11632 : tmp11717;
  assign tmp11719 = s0 ? 1 : tmp11704;
  assign tmp11718 = s1 ? tmp11704 : tmp11719;
  assign tmp11715 = s2 ? tmp11716 : tmp11718;
  assign tmp11709 = s3 ? tmp11710 : tmp11715;
  assign tmp11701 = s4 ? tmp11702 : tmp11709;
  assign tmp11726 = ~(l1 ? 1 : tmp11527);
  assign tmp11725 = ~(s0 ? 1 : tmp11726);
  assign tmp11724 = s1 ? tmp11708 : tmp11725;
  assign tmp11728 = s0 ? 1 : tmp11726;
  assign tmp11729 = ~(s0 ? tmp11704 : 0);
  assign tmp11727 = ~(s1 ? tmp11728 : tmp11729);
  assign tmp11723 = s2 ? tmp11724 : tmp11727;
  assign tmp11732 = s0 ? tmp11704 : 1;
  assign tmp11731 = ~(s1 ? 1 : tmp11732);
  assign tmp11730 = ~(s2 ? tmp11728 : tmp11731);
  assign tmp11722 = s3 ? tmp11723 : tmp11730;
  assign tmp11735 = s1 ? tmp11719 : tmp11646;
  assign tmp11736 = s1 ? tmp11646 : tmp11712;
  assign tmp11734 = s2 ? tmp11735 : tmp11736;
  assign tmp11738 = s1 ? tmp11732 : 1;
  assign tmp11737 = s2 ? tmp11738 : 1;
  assign tmp11733 = s3 ? tmp11734 : tmp11737;
  assign tmp11721 = s4 ? tmp11722 : tmp11733;
  assign tmp11741 = s2 ? tmp11738 : tmp11719;
  assign tmp11740 = s3 ? tmp11741 : 1;
  assign tmp11744 = s1 ? tmp11719 : tmp11732;
  assign tmp11743 = s2 ? 1 : tmp11744;
  assign tmp11742 = s3 ? tmp11743 : 1;
  assign tmp11739 = s4 ? tmp11740 : tmp11742;
  assign tmp11720 = s5 ? tmp11721 : tmp11739;
  assign tmp11700 = s6 ? tmp11701 : tmp11720;
  assign tmp11749 = s1 ? tmp11708 : tmp11632;
  assign tmp11748 = s2 ? tmp11711 : tmp11749;
  assign tmp11750 = s2 ? tmp11665 : tmp11718;
  assign tmp11747 = s3 ? tmp11748 : tmp11750;
  assign tmp11746 = s4 ? tmp11702 : tmp11747;
  assign tmp11755 = s1 ? tmp11704 : tmp11708;
  assign tmp11754 = s2 ? tmp11707 : tmp11755;
  assign tmp11757 = s1 ? 1 : tmp11732;
  assign tmp11756 = s2 ? tmp11704 : tmp11757;
  assign tmp11753 = s3 ? tmp11754 : tmp11756;
  assign tmp11759 = s2 ? tmp11735 : tmp11704;
  assign tmp11758 = s3 ? tmp11759 : tmp11737;
  assign tmp11752 = s4 ? tmp11753 : tmp11758;
  assign tmp11763 = s1 ? tmp11704 : tmp11732;
  assign tmp11762 = s2 ? 1 : tmp11763;
  assign tmp11761 = s3 ? tmp11762 : 1;
  assign tmp11760 = s4 ? tmp11740 : tmp11761;
  assign tmp11751 = s5 ? tmp11752 : tmp11760;
  assign tmp11745 = s6 ? tmp11746 : tmp11751;
  assign tmp11699 = s7 ? tmp11700 : tmp11745;
  assign tmp11769 = ~(l3 ? 1 : 0);
  assign tmp11768 = l1 ? 1 : tmp11769;
  assign tmp11772 = s0 ? tmp11768 : tmp11769;
  assign tmp11771 = s1 ? tmp11772 : tmp11768;
  assign tmp11770 = s2 ? tmp11768 : tmp11771;
  assign tmp11767 = s3 ? tmp11768 : tmp11770;
  assign tmp11776 = s0 ? tmp11768 : tmp11632;
  assign tmp11775 = s1 ? tmp11776 : tmp11768;
  assign tmp11777 = s0 ? tmp11768 : 0;
  assign tmp11774 = s2 ? tmp11775 : tmp11777;
  assign tmp11779 = s1 ? tmp11768 : tmp11717;
  assign tmp11781 = s0 ? 1 : tmp11768;
  assign tmp11780 = s1 ? tmp11768 : tmp11781;
  assign tmp11778 = s2 ? tmp11779 : tmp11780;
  assign tmp11773 = s3 ? tmp11774 : tmp11778;
  assign tmp11766 = s4 ? tmp11767 : tmp11773;
  assign tmp11788 = ~(l1 ? 1 : tmp11769);
  assign tmp11787 = ~(s0 ? 1 : tmp11788);
  assign tmp11786 = s1 ? tmp11777 : tmp11787;
  assign tmp11790 = s0 ? 1 : tmp11788;
  assign tmp11791 = ~(s0 ? tmp11768 : tmp11769);
  assign tmp11789 = ~(s1 ? tmp11790 : tmp11791);
  assign tmp11785 = s2 ? tmp11786 : tmp11789;
  assign tmp11793 = s0 ? tmp11479 : tmp11788;
  assign tmp11794 = ~(s1 ? 1 : tmp11768);
  assign tmp11792 = ~(s2 ? tmp11793 : tmp11794);
  assign tmp11784 = s3 ? tmp11785 : tmp11792;
  assign tmp11797 = s1 ? tmp11781 : tmp11646;
  assign tmp11798 = s1 ? tmp11646 : tmp11776;
  assign tmp11796 = s2 ? tmp11797 : tmp11798;
  assign tmp11800 = s1 ? tmp11768 : 1;
  assign tmp11799 = s2 ? tmp11800 : 1;
  assign tmp11795 = s3 ? tmp11796 : tmp11799;
  assign tmp11783 = s4 ? tmp11784 : tmp11795;
  assign tmp11805 = s0 ? tmp11768 : 1;
  assign tmp11804 = s1 ? tmp11805 : 1;
  assign tmp11803 = s2 ? tmp11804 : tmp11781;
  assign tmp11802 = s3 ? tmp11803 : 1;
  assign tmp11808 = s1 ? tmp11781 : tmp11805;
  assign tmp11807 = s2 ? 1 : tmp11808;
  assign tmp11806 = s3 ? tmp11807 : 1;
  assign tmp11801 = s4 ? tmp11802 : tmp11806;
  assign tmp11782 = s5 ? tmp11783 : tmp11801;
  assign tmp11765 = s6 ? tmp11766 : tmp11782;
  assign tmp11813 = s1 ? tmp11777 : tmp11768;
  assign tmp11812 = s2 ? tmp11775 : tmp11813;
  assign tmp11814 = s2 ? tmp11800 : tmp11780;
  assign tmp11811 = s3 ? tmp11812 : tmp11814;
  assign tmp11810 = s4 ? tmp11767 : tmp11811;
  assign tmp11819 = s1 ? tmp11768 : tmp11772;
  assign tmp11818 = s2 ? tmp11813 : tmp11819;
  assign tmp11821 = s1 ? 1 : tmp11768;
  assign tmp11820 = s2 ? tmp11768 : tmp11821;
  assign tmp11817 = s3 ? tmp11818 : tmp11820;
  assign tmp11823 = s2 ? tmp11797 : tmp11768;
  assign tmp11822 = s3 ? tmp11823 : tmp11799;
  assign tmp11816 = s4 ? tmp11817 : tmp11822;
  assign tmp11826 = s2 ? tmp11804 : tmp11800;
  assign tmp11825 = s3 ? tmp11826 : 1;
  assign tmp11828 = s2 ? 1 : tmp11800;
  assign tmp11827 = s3 ? tmp11828 : 1;
  assign tmp11824 = s4 ? tmp11825 : tmp11827;
  assign tmp11815 = s5 ? tmp11816 : tmp11824;
  assign tmp11809 = s6 ? tmp11810 : tmp11815;
  assign tmp11764 = s7 ? tmp11765 : tmp11809;
  assign tmp11698 = s8 ? tmp11699 : tmp11764;
  assign tmp11835 = s1 ? tmp11714 : tmp11632;
  assign tmp11834 = s2 ? tmp11632 : tmp11835;
  assign tmp11833 = s3 ? tmp11632 : tmp11834;
  assign tmp11837 = s2 ? tmp11632 : tmp11714;
  assign tmp11839 = s1 ? tmp11632 : tmp11648;
  assign tmp11838 = s2 ? tmp11716 : tmp11839;
  assign tmp11836 = s3 ? tmp11837 : tmp11838;
  assign tmp11832 = s4 ? tmp11833 : tmp11836;
  assign tmp11845 = ~(s0 ? 1 : tmp11623);
  assign tmp11844 = s1 ? tmp11714 : tmp11845;
  assign tmp11846 = ~(s1 ? tmp11634 : tmp11631);
  assign tmp11843 = s2 ? tmp11844 : tmp11846;
  assign tmp11848 = ~(s1 ? 1 : tmp11705);
  assign tmp11847 = ~(s2 ? tmp11634 : tmp11848);
  assign tmp11842 = s3 ? tmp11843 : tmp11847;
  assign tmp11851 = s1 ? tmp11648 : tmp11646;
  assign tmp11852 = s1 ? tmp11646 : tmp11632;
  assign tmp11850 = s2 ? tmp11851 : tmp11852;
  assign tmp11854 = s1 ? tmp11705 : 1;
  assign tmp11853 = s2 ? tmp11854 : 1;
  assign tmp11849 = s3 ? tmp11850 : tmp11853;
  assign tmp11841 = s4 ? tmp11842 : tmp11849;
  assign tmp11858 = s1 ? tmp11648 : tmp11712;
  assign tmp11857 = s2 ? tmp11645 : tmp11858;
  assign tmp11856 = s3 ? tmp11857 : 1;
  assign tmp11861 = s1 ? tmp11648 : tmp11705;
  assign tmp11860 = s2 ? 1 : tmp11861;
  assign tmp11859 = s3 ? tmp11860 : 1;
  assign tmp11855 = s4 ? tmp11856 : tmp11859;
  assign tmp11840 = s5 ? tmp11841 : tmp11855;
  assign tmp11831 = s6 ? tmp11832 : tmp11840;
  assign tmp11865 = s2 ? tmp11665 : tmp11839;
  assign tmp11864 = s3 ? tmp11834 : tmp11865;
  assign tmp11863 = s4 ? tmp11833 : tmp11864;
  assign tmp11870 = s1 ? tmp11632 : tmp11714;
  assign tmp11869 = s2 ? tmp11835 : tmp11870;
  assign tmp11872 = s1 ? 1 : tmp11705;
  assign tmp11871 = s2 ? tmp11632 : tmp11872;
  assign tmp11868 = s3 ? tmp11869 : tmp11871;
  assign tmp11874 = s2 ? tmp11851 : tmp11632;
  assign tmp11873 = s3 ? tmp11874 : tmp11853;
  assign tmp11867 = s4 ? tmp11868 : tmp11873;
  assign tmp11878 = s1 ? tmp11632 : tmp11704;
  assign tmp11877 = s2 ? 1 : tmp11878;
  assign tmp11876 = s3 ? tmp11877 : 1;
  assign tmp11875 = s4 ? tmp11667 : tmp11876;
  assign tmp11866 = s5 ? tmp11867 : tmp11875;
  assign tmp11862 = s6 ? tmp11863 : tmp11866;
  assign tmp11830 = s7 ? tmp11831 : tmp11862;
  assign tmp11829 = s8 ? tmp11764 : tmp11830;
  assign tmp11697 = s9 ? tmp11698 : tmp11829;
  assign tmp11887 = s1 ? tmp11704 : 1;
  assign tmp11886 = s2 ? tmp11738 : tmp11887;
  assign tmp11885 = s3 ? tmp11886 : 1;
  assign tmp11889 = s2 ? 1 : tmp11887;
  assign tmp11888 = s3 ? tmp11889 : 1;
  assign tmp11884 = s4 ? tmp11885 : tmp11888;
  assign tmp11883 = s5 ? tmp11752 : tmp11884;
  assign tmp11882 = s6 ? tmp11746 : tmp11883;
  assign tmp11881 = s7 ? tmp11700 : tmp11882;
  assign tmp11880 = s8 ? tmp11881 : tmp11700;
  assign tmp11896 = s2 ? 1 : tmp11704;
  assign tmp11895 = s3 ? tmp11896 : 1;
  assign tmp11894 = s4 ? tmp11740 : tmp11895;
  assign tmp11893 = s5 ? tmp11752 : tmp11894;
  assign tmp11892 = s6 ? tmp11746 : tmp11893;
  assign tmp11899 = s4 ? tmp11667 : tmp11669;
  assign tmp11898 = s5 ? tmp11867 : tmp11899;
  assign tmp11897 = s6 ? tmp11863 : tmp11898;
  assign tmp11891 = s7 ? tmp11892 : tmp11897;
  assign tmp11905 = s2 ? 1 : tmp11768;
  assign tmp11904 = s3 ? tmp11905 : 1;
  assign tmp11903 = s4 ? tmp11825 : tmp11904;
  assign tmp11902 = s5 ? tmp11816 : tmp11903;
  assign tmp11901 = s6 ? tmp11810 : tmp11902;
  assign tmp11908 = s4 ? tmp11885 : tmp11895;
  assign tmp11907 = s5 ? tmp11752 : tmp11908;
  assign tmp11906 = s6 ? tmp11746 : tmp11907;
  assign tmp11900 = s7 ? tmp11901 : tmp11906;
  assign tmp11890 = s8 ? tmp11891 : tmp11900;
  assign tmp11879 = s9 ? tmp11880 : tmp11890;
  assign tmp11696 = s10 ? tmp11697 : tmp11879;
  assign tmp11912 = s7 ? tmp11745 : tmp11862;
  assign tmp11913 = s7 ? tmp11809 : tmp11882;
  assign tmp11911 = s8 ? tmp11912 : tmp11913;
  assign tmp11910 = s9 ? tmp11880 : tmp11911;
  assign tmp11909 = s10 ? tmp11697 : tmp11910;
  assign tmp11695 = s11 ? tmp11696 : tmp11909;
  assign tmp11694 = ~(s12 ? tmp11695 : 1);
  assign tmp11692 = s13 ? tmp11693 : tmp11694;
  assign tmp11467 = s14 ? tmp11468 : tmp11692;
  assign tmp11924 = ~(l2 ? 1 : tmp11769);
  assign tmp11923 = l1 ? 1 : tmp11924;
  assign tmp11922 = s1 ? tmp11923 : tmp11845;
  assign tmp11928 = ~(l1 ? 1 : tmp11924);
  assign tmp11927 = s0 ? 1 : tmp11928;
  assign tmp11929 = ~(s0 ? tmp11632 : tmp11923);
  assign tmp11926 = s1 ? tmp11927 : tmp11929;
  assign tmp11930 = ~(s1 ? tmp11714 : tmp11923);
  assign tmp11925 = ~(s2 ? tmp11926 : tmp11930);
  assign tmp11921 = s3 ? tmp11922 : tmp11925;
  assign tmp11933 = s1 ? 1 : tmp11928;
  assign tmp11935 = s0 ? tmp11923 : 0;
  assign tmp11934 = ~(s1 ? tmp11935 : 0);
  assign tmp11932 = s2 ? tmp11933 : tmp11934;
  assign tmp11937 = s1 ? 1 : tmp11927;
  assign tmp11936 = s2 ? tmp11937 : tmp11928;
  assign tmp11931 = ~(s3 ? tmp11932 : tmp11936);
  assign tmp11920 = s4 ? tmp11921 : tmp11931;
  assign tmp11942 = s1 ? tmp11714 : 0;
  assign tmp11944 = ~(s0 ? tmp11923 : 0);
  assign tmp11943 = ~(s1 ? tmp11634 : tmp11944);
  assign tmp11941 = s2 ? tmp11942 : tmp11943;
  assign tmp11946 = s1 ? tmp11634 : tmp11927;
  assign tmp11945 = ~(s2 ? tmp11946 : tmp11928);
  assign tmp11940 = s3 ? tmp11941 : tmp11945;
  assign tmp11949 = s1 ? tmp11923 : 0;
  assign tmp11948 = s2 ? tmp11949 : 0;
  assign tmp11950 = ~(s2 ? tmp11927 : tmp11928);
  assign tmp11947 = s3 ? tmp11948 : tmp11950;
  assign tmp11939 = s4 ? tmp11940 : tmp11947;
  assign tmp11955 = s0 ? tmp11923 : tmp11632;
  assign tmp11954 = s1 ? tmp11955 : tmp11648;
  assign tmp11953 = s2 ? tmp11954 : tmp11942;
  assign tmp11958 = s0 ? 1 : tmp11769;
  assign tmp11959 = ~(s0 ? tmp11479 : 1);
  assign tmp11957 = s1 ? tmp11958 : tmp11959;
  assign tmp11960 = ~(s1 ? tmp11923 : tmp11935);
  assign tmp11956 = ~(s2 ? tmp11957 : tmp11960);
  assign tmp11952 = s3 ? tmp11953 : tmp11956;
  assign tmp11963 = s1 ? tmp11634 : tmp11929;
  assign tmp11964 = ~(s1 ? tmp11648 : 0);
  assign tmp11962 = s2 ? tmp11963 : tmp11964;
  assign tmp11968 = l1 ? 1 : tmp11479;
  assign tmp11967 = s0 ? tmp11632 : tmp11968;
  assign tmp11966 = s1 ? tmp11967 : tmp11923;
  assign tmp11970 = s0 ? tmp11479 : tmp11632;
  assign tmp11969 = s1 ? tmp11935 : tmp11970;
  assign tmp11965 = ~(s2 ? tmp11966 : tmp11969);
  assign tmp11961 = ~(s3 ? tmp11962 : tmp11965);
  assign tmp11951 = s4 ? tmp11952 : tmp11961;
  assign tmp11938 = s5 ? tmp11939 : tmp11951;
  assign tmp11919 = s6 ? tmp11920 : tmp11938;
  assign tmp11974 = s2 ? tmp11933 : tmp11928;
  assign tmp11973 = ~(s3 ? tmp11932 : tmp11974);
  assign tmp11972 = s4 ? tmp11921 : tmp11973;
  assign tmp11979 = s1 ? tmp11632 : tmp11935;
  assign tmp11978 = s2 ? tmp11942 : tmp11979;
  assign tmp11981 = s1 ? tmp11632 : tmp11923;
  assign tmp11980 = s2 ? tmp11981 : tmp11923;
  assign tmp11977 = s3 ? tmp11978 : tmp11980;
  assign tmp11976 = s4 ? tmp11977 : tmp11947;
  assign tmp11985 = s1 ? tmp11955 : tmp11632;
  assign tmp11984 = s2 ? tmp11985 : 0;
  assign tmp11987 = s1 ? tmp11479 : 1;
  assign tmp11988 = s1 ? tmp11923 : tmp11935;
  assign tmp11986 = s2 ? tmp11987 : tmp11988;
  assign tmp11983 = s3 ? tmp11984 : tmp11986;
  assign tmp11990 = s2 ? tmp11981 : tmp11632;
  assign tmp11989 = s3 ? tmp11990 : tmp11923;
  assign tmp11982 = s4 ? tmp11983 : tmp11989;
  assign tmp11975 = s5 ? tmp11976 : tmp11982;
  assign tmp11971 = s6 ? tmp11972 : tmp11975;
  assign tmp11918 = s7 ? tmp11919 : tmp11971;
  assign tmp11992 = s8 ? tmp11918 : tmp11919;
  assign tmp11991 = s9 ? tmp11992 : tmp11971;
  assign tmp11917 = s10 ? tmp11918 : tmp11991;
  assign tmp12001 = s0 ? 1 : tmp11479;
  assign tmp12000 = s1 ? 1 : tmp12001;
  assign tmp12003 = s0 ? 1 : tmp11482;
  assign tmp12004 = s1 ? 1 : tmp11482;
  assign tmp12002 = s2 ? tmp12003 : tmp12004;
  assign tmp11999 = s3 ? tmp12000 : tmp12002;
  assign tmp12006 = s2 ? tmp12004 : 1;
  assign tmp12007 = s2 ? tmp12004 : tmp11482;
  assign tmp12005 = s3 ? tmp12006 : tmp12007;
  assign tmp11998 = s4 ? tmp11999 : tmp12005;
  assign tmp12012 = s1 ? tmp11479 : tmp11491;
  assign tmp12011 = s2 ? tmp11987 : tmp12012;
  assign tmp12014 = s1 ? 1 : tmp12003;
  assign tmp12013 = s2 ? tmp12014 : tmp11482;
  assign tmp12010 = s3 ? tmp12011 : tmp12013;
  assign tmp12017 = s1 ? tmp11482 : 1;
  assign tmp12016 = s2 ? tmp12017 : 1;
  assign tmp12019 = s1 ? 1 : tmp11491;
  assign tmp12018 = s2 ? tmp12014 : tmp12019;
  assign tmp12015 = s3 ? tmp12016 : tmp12018;
  assign tmp12009 = s4 ? tmp12010 : tmp12015;
  assign tmp12022 = s2 ? tmp11482 : 1;
  assign tmp12025 = s0 ? tmp11632 : tmp11625;
  assign tmp12024 = s1 ? tmp11632 : tmp12025;
  assign tmp12026 = ~(s1 ? tmp11482 : 1);
  assign tmp12023 = ~(s2 ? tmp12024 : tmp12026);
  assign tmp12021 = s3 ? tmp12022 : tmp12023;
  assign tmp12029 = s1 ? tmp12001 : tmp11482;
  assign tmp12030 = s1 ? tmp12001 : 1;
  assign tmp12028 = s2 ? tmp12029 : tmp12030;
  assign tmp12032 = s1 ? tmp12003 : tmp11482;
  assign tmp12034 = ~(s0 ? tmp11632 : tmp11769);
  assign tmp12033 = s1 ? 1 : tmp12034;
  assign tmp12031 = s2 ? tmp12032 : tmp12033;
  assign tmp12027 = s3 ? tmp12028 : tmp12031;
  assign tmp12020 = s4 ? tmp12021 : tmp12027;
  assign tmp12008 = s5 ? tmp12009 : tmp12020;
  assign tmp11997 = s6 ? tmp11998 : tmp12008;
  assign tmp12038 = s3 ? tmp12011 : tmp12007;
  assign tmp12039 = s3 ? tmp12016 : tmp12004;
  assign tmp12037 = s4 ? tmp12038 : tmp12039;
  assign tmp12043 = s1 ? tmp11632 : tmp11625;
  assign tmp12042 = ~(s2 ? tmp12043 : tmp12026);
  assign tmp12041 = s3 ? tmp12016 : tmp12042;
  assign tmp12045 = s2 ? tmp11482 : tmp11479;
  assign tmp12044 = s3 ? tmp12045 : tmp11482;
  assign tmp12040 = s4 ? tmp12041 : tmp12044;
  assign tmp12036 = s5 ? tmp12037 : tmp12040;
  assign tmp12035 = s6 ? tmp11998 : tmp12036;
  assign tmp11996 = s7 ? tmp11997 : tmp12035;
  assign tmp12049 = s3 ? tmp12006 : tmp12013;
  assign tmp12048 = s4 ? tmp11999 : tmp12049;
  assign tmp12047 = s6 ? tmp12048 : tmp12008;
  assign tmp12046 = s7 ? tmp12047 : tmp12035;
  assign tmp11995 = s8 ? tmp11996 : tmp12046;
  assign tmp11994 = s9 ? tmp11995 : tmp12046;
  assign tmp12051 = s8 ? tmp12046 : tmp12047;
  assign tmp12050 = s9 ? tmp12051 : tmp12035;
  assign tmp11993 = s10 ? tmp11994 : tmp12050;
  assign tmp11916 = s12 ? tmp11917 : tmp11993;
  assign tmp11915 = s13 ? 1 : tmp11916;
  assign tmp12063 = l1 ? tmp11480 : 1;
  assign tmp12062 = s0 ? 1 : tmp12063;
  assign tmp12065 = s1 ? tmp12062 : tmp12063;
  assign tmp12067 = s0 ? tmp12063 : 1;
  assign tmp12066 = s1 ? tmp12067 : tmp12063;
  assign tmp12064 = s2 ? tmp12065 : tmp12066;
  assign tmp12061 = s3 ? tmp12062 : tmp12064;
  assign tmp12070 = s1 ? 1 : tmp12063;
  assign tmp12071 = s1 ? tmp12067 : 1;
  assign tmp12069 = s2 ? tmp12070 : tmp12071;
  assign tmp12073 = s1 ? 1 : tmp11634;
  assign tmp12072 = s2 ? tmp12073 : tmp12063;
  assign tmp12068 = s3 ? tmp12069 : tmp12072;
  assign tmp12060 = s4 ? tmp12061 : tmp12068;
  assign tmp12078 = s1 ? tmp12062 : tmp12067;
  assign tmp12077 = s2 ? tmp12071 : tmp12078;
  assign tmp12081 = s0 ? tmp12063 : 0;
  assign tmp12080 = s1 ? tmp12081 : tmp12063;
  assign tmp12079 = s2 ? tmp12062 : tmp12080;
  assign tmp12076 = s3 ? tmp12077 : tmp12079;
  assign tmp12086 = ~(l1 ? tmp11480 : 1);
  assign tmp12085 = s0 ? tmp11632 : tmp12086;
  assign tmp12084 = s1 ? tmp12085 : 0;
  assign tmp12083 = s2 ? tmp12084 : 0;
  assign tmp12088 = s1 ? tmp12063 : tmp12062;
  assign tmp12089 = ~(s1 ? 1 : tmp11646);
  assign tmp12087 = ~(s2 ? tmp12088 : tmp12089);
  assign tmp12082 = ~(s3 ? tmp12083 : tmp12087);
  assign tmp12075 = s4 ? tmp12076 : tmp12082;
  assign tmp12094 = ~(s0 ? 1 : tmp12086);
  assign tmp12093 = s1 ? tmp12081 : tmp12094;
  assign tmp12092 = s2 ? tmp12093 : tmp12071;
  assign tmp12096 = s1 ? tmp11494 : 0;
  assign tmp12097 = ~(s1 ? tmp11632 : tmp11714);
  assign tmp12095 = s2 ? tmp12096 : tmp12097;
  assign tmp12091 = s3 ? tmp12092 : tmp12095;
  assign tmp12100 = s1 ? tmp11508 : tmp12063;
  assign tmp12102 = s0 ? 1 : tmp12086;
  assign tmp12101 = ~(s1 ? tmp12102 : 0);
  assign tmp12099 = s2 ? tmp12100 : tmp12101;
  assign tmp12104 = s1 ? tmp12063 : tmp12094;
  assign tmp12105 = ~(s1 ? tmp11714 : tmp11526);
  assign tmp12103 = s2 ? tmp12104 : tmp12105;
  assign tmp12098 = s3 ? tmp12099 : tmp12103;
  assign tmp12090 = s4 ? tmp12091 : tmp12098;
  assign tmp12074 = s5 ? tmp12075 : tmp12090;
  assign tmp12059 = s6 ? tmp12060 : tmp12074;
  assign tmp12110 = s1 ? 1 : tmp11623;
  assign tmp12109 = s2 ? tmp12110 : tmp12063;
  assign tmp12108 = s3 ? tmp12069 : tmp12109;
  assign tmp12107 = s4 ? tmp12061 : tmp12108;
  assign tmp12115 = s1 ? tmp12063 : tmp12067;
  assign tmp12114 = s2 ? tmp12071 : tmp12115;
  assign tmp12116 = s2 ? tmp12063 : tmp12080;
  assign tmp12113 = s3 ? tmp12114 : tmp12116;
  assign tmp12119 = ~(s1 ? 1 : tmp11632);
  assign tmp12118 = ~(s2 ? tmp12063 : tmp12119);
  assign tmp12117 = ~(s3 ? tmp12083 : tmp12118);
  assign tmp12112 = s4 ? tmp12113 : tmp12117;
  assign tmp12122 = s2 ? tmp12080 : tmp12071;
  assign tmp12124 = s1 ? tmp11632 : 0;
  assign tmp12123 = ~(s2 ? 1 : tmp12124);
  assign tmp12121 = s3 ? tmp12122 : tmp12123;
  assign tmp12120 = s4 ? tmp12121 : tmp12063;
  assign tmp12111 = s5 ? tmp12112 : tmp12120;
  assign tmp12106 = s6 ? tmp12107 : tmp12111;
  assign tmp12058 = s7 ? tmp12059 : tmp12106;
  assign tmp12132 = s0 ? tmp11480 : tmp12063;
  assign tmp12131 = s1 ? tmp11508 : tmp12132;
  assign tmp12130 = s2 ? tmp12131 : tmp12101;
  assign tmp12135 = s0 ? tmp12063 : tmp11480;
  assign tmp12134 = s1 ? tmp12135 : tmp12094;
  assign tmp12133 = s2 ? tmp12134 : tmp12105;
  assign tmp12129 = s3 ? tmp12130 : tmp12133;
  assign tmp12128 = s4 ? tmp12091 : tmp12129;
  assign tmp12127 = s5 ? tmp12075 : tmp12128;
  assign tmp12126 = s6 ? tmp12060 : tmp12127;
  assign tmp12140 = s2 ? tmp12080 : 1;
  assign tmp12139 = s3 ? tmp12140 : tmp12123;
  assign tmp12143 = s1 ? tmp11480 : tmp12063;
  assign tmp12142 = s2 ? tmp12143 : tmp12063;
  assign tmp12141 = s3 ? tmp12142 : tmp12143;
  assign tmp12138 = s4 ? tmp12139 : tmp12141;
  assign tmp12137 = s5 ? tmp12112 : tmp12138;
  assign tmp12136 = s6 ? tmp12107 : tmp12137;
  assign tmp12125 = s7 ? tmp12126 : tmp12136;
  assign tmp12057 = s8 ? tmp12058 : tmp12125;
  assign tmp12148 = s4 ? tmp12139 : tmp12063;
  assign tmp12147 = s5 ? tmp12112 : tmp12148;
  assign tmp12146 = s6 ? tmp12107 : tmp12147;
  assign tmp12145 = s7 ? tmp12059 : tmp12146;
  assign tmp12144 = s8 ? tmp12125 : tmp12145;
  assign tmp12056 = s9 ? tmp12057 : tmp12144;
  assign tmp12155 = s3 ? tmp12063 : tmp12143;
  assign tmp12154 = s4 ? tmp12139 : tmp12155;
  assign tmp12153 = s5 ? tmp12112 : tmp12154;
  assign tmp12152 = s6 ? tmp12107 : tmp12153;
  assign tmp12151 = s7 ? tmp12059 : tmp12152;
  assign tmp12150 = s8 ? tmp12151 : tmp12059;
  assign tmp12160 = s4 ? tmp12121 : tmp12155;
  assign tmp12159 = s5 ? tmp12112 : tmp12160;
  assign tmp12158 = s6 ? tmp12107 : tmp12159;
  assign tmp12157 = s7 ? tmp12158 : tmp12146;
  assign tmp12161 = s7 ? tmp12136 : tmp12152;
  assign tmp12156 = s8 ? tmp12157 : tmp12161;
  assign tmp12149 = s9 ? tmp12150 : tmp12156;
  assign tmp12055 = s10 ? tmp12056 : tmp12149;
  assign tmp12165 = s7 ? tmp12106 : tmp12146;
  assign tmp12164 = s8 ? tmp12165 : tmp12161;
  assign tmp12163 = s9 ? tmp12150 : tmp12164;
  assign tmp12162 = s10 ? tmp12056 : tmp12163;
  assign tmp12054 = s11 ? tmp12055 : tmp12162;
  assign tmp12053 = s12 ? 1 : tmp12054;
  assign tmp12172 = s1 ? tmp11479 : 0;
  assign tmp12173 = ~(s2 ? tmp11781 : tmp11821);
  assign tmp12171 = s3 ? tmp12172 : tmp12173;
  assign tmp12177 = s0 ? tmp11479 : 0;
  assign tmp12176 = ~(s1 ? tmp12177 : 0);
  assign tmp12175 = s2 ? tmp11821 : tmp12176;
  assign tmp12179 = s1 ? 1 : tmp11781;
  assign tmp12178 = s2 ? tmp12179 : tmp11768;
  assign tmp12174 = ~(s3 ? tmp12175 : tmp12178);
  assign tmp12170 = s4 ? tmp12171 : tmp12174;
  assign tmp12184 = s1 ? 1 : tmp11805;
  assign tmp12183 = s2 ? 1 : tmp12184;
  assign tmp12182 = s3 ? tmp12183 : tmp12178;
  assign tmp12186 = s2 ? tmp11781 : tmp11768;
  assign tmp12185 = s3 ? tmp11799 : tmp12186;
  assign tmp12181 = s4 ? tmp12182 : tmp12185;
  assign tmp12190 = s1 ? tmp11777 : tmp11717;
  assign tmp12189 = s2 ? tmp12190 : 1;
  assign tmp12192 = s1 ? tmp11781 : tmp11768;
  assign tmp12194 = ~(s0 ? tmp11479 : 0);
  assign tmp12193 = s1 ? tmp11768 : tmp12194;
  assign tmp12191 = s2 ? tmp12192 : tmp12193;
  assign tmp12188 = s3 ? tmp12189 : tmp12191;
  assign tmp12197 = ~(s1 ? tmp11494 : 0);
  assign tmp12196 = s2 ? tmp12179 : tmp12197;
  assign tmp12198 = s2 ? tmp12192 : tmp11805;
  assign tmp12195 = s3 ? tmp12196 : tmp12198;
  assign tmp12187 = s4 ? tmp12188 : tmp12195;
  assign tmp12180 = ~(s5 ? tmp12181 : tmp12187);
  assign tmp12169 = s6 ? tmp12170 : tmp12180;
  assign tmp12202 = s2 ? tmp11821 : tmp11768;
  assign tmp12201 = ~(s3 ? tmp12175 : tmp12202);
  assign tmp12200 = s4 ? tmp12171 : tmp12201;
  assign tmp12205 = s3 ? tmp12183 : tmp12202;
  assign tmp12204 = s4 ? tmp12205 : tmp12185;
  assign tmp12209 = s1 ? tmp11777 : 1;
  assign tmp12208 = s2 ? tmp12209 : 1;
  assign tmp12211 = ~(s1 ? tmp11479 : 0);
  assign tmp12210 = s2 ? tmp11768 : tmp12211;
  assign tmp12207 = s3 ? tmp12208 : tmp12210;
  assign tmp12213 = s2 ? tmp11821 : 1;
  assign tmp12212 = s3 ? tmp12213 : tmp11768;
  assign tmp12206 = s4 ? tmp12207 : tmp12212;
  assign tmp12203 = ~(s5 ? tmp12204 : tmp12206);
  assign tmp12199 = s6 ? tmp12200 : tmp12203;
  assign tmp12168 = s7 ? tmp12169 : tmp12199;
  assign tmp12215 = s8 ? tmp12168 : tmp12169;
  assign tmp12214 = s9 ? tmp12215 : tmp12199;
  assign tmp12167 = s10 ? tmp12168 : tmp12214;
  assign tmp12225 = l2 ? 1 : tmp11769;
  assign tmp12224 = l1 ? tmp12225 : 1;
  assign tmp12223 = s0 ? 1 : tmp12224;
  assign tmp12227 = s1 ? tmp12223 : tmp12224;
  assign tmp12228 = s1 ? tmp12063 : tmp12224;
  assign tmp12226 = s2 ? tmp12227 : tmp12228;
  assign tmp12222 = s3 ? tmp12223 : tmp12226;
  assign tmp12231 = s1 ? 1 : tmp12224;
  assign tmp12230 = s2 ? tmp12231 : tmp12071;
  assign tmp12235 = ~(l1 ? tmp11479 : 0);
  assign tmp12234 = s0 ? 1 : tmp12235;
  assign tmp12233 = s1 ? 1 : tmp12234;
  assign tmp12232 = s2 ? tmp12233 : tmp12224;
  assign tmp12229 = s3 ? tmp12230 : tmp12232;
  assign tmp12221 = s4 ? tmp12222 : tmp12229;
  assign tmp12241 = s0 ? tmp12224 : 1;
  assign tmp12240 = s1 ? tmp12241 : 1;
  assign tmp12246 = ~(l4 ? 1 : 0);
  assign tmp12245 = ~(l2 ? 1 : tmp12246);
  assign tmp12244 = l1 ? tmp11480 : tmp12245;
  assign tmp12243 = s0 ? tmp12224 : tmp12244;
  assign tmp12242 = s1 ? tmp12223 : tmp12243;
  assign tmp12239 = s2 ? tmp12240 : tmp12242;
  assign tmp12248 = s0 ? tmp12244 : tmp12224;
  assign tmp12247 = s2 ? tmp12248 : tmp12224;
  assign tmp12238 = s3 ? tmp12239 : tmp12247;
  assign tmp12251 = s1 ? tmp12224 : 1;
  assign tmp12250 = s2 ? tmp12251 : 1;
  assign tmp12255 = l1 ? tmp11479 : 0;
  assign tmp12254 = s0 ? tmp12255 : 1;
  assign tmp12253 = ~(s1 ? 1 : tmp12254);
  assign tmp12252 = s2 ? tmp12223 : tmp12253;
  assign tmp12249 = s3 ? tmp12250 : tmp12252;
  assign tmp12237 = s4 ? tmp12238 : tmp12249;
  assign tmp12258 = s2 ? tmp12224 : tmp12071;
  assign tmp12260 = s1 ? 1 : tmp11958;
  assign tmp12261 = ~(s1 ? tmp12255 : tmp11714);
  assign tmp12259 = s2 ? tmp12260 : tmp12261;
  assign tmp12257 = s3 ? tmp12258 : tmp12259;
  assign tmp12263 = s2 ? tmp12227 : tmp12251;
  assign tmp12266 = ~(s0 ? 1 : tmp12224);
  assign tmp12265 = ~(s1 ? tmp11714 : tmp12266);
  assign tmp12264 = s2 ? tmp12224 : tmp12265;
  assign tmp12262 = s3 ? tmp12263 : tmp12264;
  assign tmp12256 = s4 ? tmp12257 : tmp12262;
  assign tmp12236 = s5 ? tmp12237 : tmp12256;
  assign tmp12220 = s6 ? tmp12221 : tmp12236;
  assign tmp12271 = s1 ? 1 : tmp12235;
  assign tmp12270 = s2 ? tmp12271 : tmp12224;
  assign tmp12269 = s3 ? tmp12230 : tmp12270;
  assign tmp12268 = s4 ? tmp12222 : tmp12269;
  assign tmp12276 = s1 ? tmp12224 : tmp12243;
  assign tmp12275 = s2 ? tmp12240 : tmp12276;
  assign tmp12274 = s3 ? tmp12275 : tmp12224;
  assign tmp12279 = ~(s1 ? 1 : tmp12255);
  assign tmp12278 = s2 ? tmp12223 : tmp12279;
  assign tmp12277 = s3 ? tmp12250 : tmp12278;
  assign tmp12273 = s4 ? tmp12274 : tmp12277;
  assign tmp12283 = s1 ? tmp12224 : tmp12063;
  assign tmp12282 = s2 ? tmp12283 : 1;
  assign tmp12285 = s1 ? 1 : tmp11769;
  assign tmp12286 = ~(s1 ? tmp11632 : 0);
  assign tmp12284 = s2 ? tmp12285 : tmp12286;
  assign tmp12281 = s3 ? tmp12282 : tmp12284;
  assign tmp12280 = s4 ? tmp12281 : tmp12224;
  assign tmp12272 = s5 ? tmp12273 : tmp12280;
  assign tmp12267 = s6 ? tmp12268 : tmp12272;
  assign tmp12219 = s7 ? tmp12220 : tmp12267;
  assign tmp12292 = s1 ? tmp12067 : tmp12224;
  assign tmp12291 = s2 ? tmp12227 : tmp12292;
  assign tmp12290 = s3 ? tmp12223 : tmp12291;
  assign tmp12299 = l3 ? 1 : tmp12246;
  assign tmp12298 = l2 ? tmp12299 : 1;
  assign tmp12297 = l1 ? 1 : tmp12298;
  assign tmp12296 = s0 ? tmp12063 : tmp12297;
  assign tmp12295 = s1 ? tmp12296 : 1;
  assign tmp12294 = s2 ? tmp12231 : tmp12295;
  assign tmp12293 = s3 ? tmp12294 : tmp12232;
  assign tmp12289 = s4 ? tmp12290 : tmp12293;
  assign tmp12304 = s1 ? tmp12223 : tmp12241;
  assign tmp12303 = s2 ? tmp12240 : tmp12304;
  assign tmp12305 = s2 ? tmp12223 : tmp12224;
  assign tmp12302 = s3 ? tmp12303 : tmp12305;
  assign tmp12301 = s4 ? tmp12302 : tmp12249;
  assign tmp12300 = s5 ? tmp12301 : tmp12256;
  assign tmp12288 = s6 ? tmp12289 : tmp12300;
  assign tmp12308 = s3 ? tmp12294 : tmp12270;
  assign tmp12307 = s4 ? tmp12290 : tmp12308;
  assign tmp12313 = s1 ? tmp12224 : tmp12241;
  assign tmp12312 = s2 ? tmp12240 : tmp12313;
  assign tmp12311 = s3 ? tmp12312 : tmp12224;
  assign tmp12310 = s4 ? tmp12311 : tmp12277;
  assign tmp12309 = s5 ? tmp12310 : tmp12280;
  assign tmp12306 = s6 ? tmp12307 : tmp12309;
  assign tmp12287 = s7 ? tmp12288 : tmp12306;
  assign tmp12218 = s8 ? tmp12219 : tmp12287;
  assign tmp12317 = s4 ? tmp12290 : tmp12229;
  assign tmp12316 = s6 ? tmp12317 : tmp12300;
  assign tmp12319 = s4 ? tmp12290 : tmp12269;
  assign tmp12318 = s6 ? tmp12319 : tmp12309;
  assign tmp12315 = s7 ? tmp12316 : tmp12318;
  assign tmp12314 = s8 ? tmp12287 : tmp12315;
  assign tmp12217 = s9 ? tmp12218 : tmp12314;
  assign tmp12330 = l1 ? 1 : tmp12246;
  assign tmp12329 = s0 ? tmp12330 : tmp12224;
  assign tmp12328 = s1 ? tmp12062 : tmp12329;
  assign tmp12327 = s2 ? tmp12328 : tmp12253;
  assign tmp12326 = s3 ? tmp12250 : tmp12327;
  assign tmp12325 = s4 ? tmp12302 : tmp12326;
  assign tmp12324 = s5 ? tmp12325 : tmp12256;
  assign tmp12323 = s6 ? tmp12317 : tmp12324;
  assign tmp12322 = s7 ? tmp12323 : tmp12318;
  assign tmp12321 = s8 ? tmp12322 : tmp12323;
  assign tmp12332 = s7 ? tmp12267 : tmp12318;
  assign tmp12333 = s7 ? tmp12306 : tmp12318;
  assign tmp12331 = s8 ? tmp12332 : tmp12333;
  assign tmp12320 = s9 ? tmp12321 : tmp12331;
  assign tmp12216 = ~(s10 ? tmp12217 : tmp12320);
  assign tmp12166 = ~(s12 ? tmp12167 : tmp12216);
  assign tmp12052 = ~(s13 ? tmp12053 : tmp12166);
  assign tmp11914 = s14 ? tmp11915 : tmp12052;
  assign tmp11466 = s15 ? tmp11467 : tmp11914;
  assign tmp12348 = s0 ? tmp11480 : tmp11623;
  assign tmp12347 = s1 ? tmp11581 : tmp12348;
  assign tmp12346 = s2 ? tmp11580 : tmp12347;
  assign tmp12350 = s0 ? tmp11632 : tmp11527;
  assign tmp12351 = s1 ? 1 : tmp11585;
  assign tmp12349 = ~(s2 ? tmp12350 : tmp12351);
  assign tmp12345 = s3 ? tmp12346 : tmp12349;
  assign tmp12344 = s4 ? tmp12345 : tmp11587;
  assign tmp12343 = s5 ? tmp12344 : tmp11520;
  assign tmp12342 = s6 ? tmp11554 : tmp12343;
  assign tmp12357 = s1 ? tmp11557 : tmp12348;
  assign tmp12356 = s2 ? tmp11562 : tmp12357;
  assign tmp12355 = s3 ? tmp12356 : tmp11609;
  assign tmp12361 = l1 ? tmp12225 : 0;
  assign tmp12363 = ~(l1 ? tmp12225 : 0);
  assign tmp12362 = ~(s0 ? tmp11557 : tmp12363);
  assign tmp12360 = s1 ? tmp12361 : tmp12362;
  assign tmp12359 = s2 ? tmp11589 : tmp12360;
  assign tmp12358 = ~(s3 ? tmp12359 : tmp11612);
  assign tmp12354 = s4 ? tmp12355 : tmp12358;
  assign tmp12353 = s5 ? tmp12354 : tmp11547;
  assign tmp12352 = s6 ? tmp11598 : tmp12353;
  assign tmp12341 = s7 ? tmp12342 : tmp12352;
  assign tmp12340 = s8 ? tmp11473 : tmp12341;
  assign tmp12370 = s0 ? tmp12361 : tmp12063;
  assign tmp12369 = s2 ? tmp12361 : tmp12370;
  assign tmp12372 = s1 ? tmp12361 : tmp12067;
  assign tmp12374 = s0 ? tmp12361 : tmp11632;
  assign tmp12375 = s0 ? 1 : tmp12361;
  assign tmp12373 = s1 ? tmp12374 : tmp12375;
  assign tmp12371 = s2 ? tmp12372 : tmp12373;
  assign tmp12368 = s3 ? tmp12369 : tmp12371;
  assign tmp12367 = s4 ? tmp12361 : tmp12368;
  assign tmp12380 = s1 ? tmp12361 : tmp11632;
  assign tmp12379 = s2 ? tmp12361 : tmp12380;
  assign tmp12383 = s0 ? tmp12361 : 1;
  assign tmp12382 = s1 ? 1 : tmp12383;
  assign tmp12381 = s2 ? tmp11632 : tmp12382;
  assign tmp12378 = s3 ? tmp12379 : tmp12381;
  assign tmp12386 = s1 ? tmp12375 : tmp12383;
  assign tmp12387 = s1 ? tmp12383 : tmp12361;
  assign tmp12385 = s2 ? tmp12386 : tmp12387;
  assign tmp12388 = s2 ? tmp11645 : 1;
  assign tmp12384 = s3 ? tmp12385 : tmp12388;
  assign tmp12377 = s4 ? tmp12378 : tmp12384;
  assign tmp12389 = s4 ? tmp11643 : tmp11649;
  assign tmp12376 = s5 ? tmp12377 : tmp12389;
  assign tmp12366 = s6 ? tmp12367 : tmp12376;
  assign tmp12394 = s1 ? tmp12370 : tmp12361;
  assign tmp12393 = s2 ? tmp12361 : tmp12394;
  assign tmp12396 = s1 ? tmp12361 : 1;
  assign tmp12395 = s2 ? tmp12396 : tmp12373;
  assign tmp12392 = s3 ? tmp12393 : tmp12395;
  assign tmp12391 = s4 ? tmp12361 : tmp12392;
  assign tmp12400 = s2 ? tmp12386 : tmp12361;
  assign tmp12399 = s3 ? tmp12400 : tmp12388;
  assign tmp12398 = s4 ? tmp12378 : tmp12399;
  assign tmp12397 = s5 ? tmp12398 : tmp11899;
  assign tmp12390 = s6 ? tmp12391 : tmp12397;
  assign tmp12365 = ~(s7 ? tmp12366 : tmp12390);
  assign tmp12364 = s8 ? tmp12341 : tmp12365;
  assign tmp12339 = s9 ? tmp12340 : tmp12364;
  assign tmp12408 = l1 ? tmp12225 : tmp11527;
  assign tmp12409 = s0 ? tmp12361 : tmp12408;
  assign tmp12407 = s1 ? tmp12408 : tmp12409;
  assign tmp12412 = s0 ? tmp12408 : tmp11586;
  assign tmp12411 = s1 ? tmp12412 : tmp12408;
  assign tmp12410 = s2 ? tmp12408 : tmp12411;
  assign tmp12406 = s3 ? tmp12407 : tmp12410;
  assign tmp12416 = s0 ? tmp12408 : tmp12361;
  assign tmp12415 = s1 ? tmp12416 : tmp12408;
  assign tmp12418 = s0 ? tmp12408 : tmp12063;
  assign tmp12417 = s1 ? tmp12418 : tmp12370;
  assign tmp12414 = s2 ? tmp12415 : tmp12417;
  assign tmp12421 = s0 ? tmp12408 : tmp11704;
  assign tmp12422 = s0 ? 1 : tmp12408;
  assign tmp12420 = s1 ? tmp12421 : tmp12422;
  assign tmp12419 = s2 ? tmp12372 : tmp12420;
  assign tmp12413 = s3 ? tmp12414 : tmp12419;
  assign tmp12405 = s4 ? tmp12406 : tmp12413;
  assign tmp12428 = s0 ? tmp12408 : 0;
  assign tmp12430 = ~(l1 ? tmp12225 : tmp11527);
  assign tmp12429 = ~(s0 ? 1 : tmp12430);
  assign tmp12427 = s1 ? tmp12428 : tmp12429;
  assign tmp12432 = s0 ? 1 : tmp12430;
  assign tmp12433 = ~(s0 ? tmp11704 : tmp11632);
  assign tmp12431 = ~(s1 ? tmp12432 : tmp12433);
  assign tmp12426 = s2 ? tmp12427 : tmp12431;
  assign tmp12435 = s1 ? tmp11705 : tmp12350;
  assign tmp12437 = s0 ? tmp12408 : 1;
  assign tmp12436 = s1 ? 1 : tmp12437;
  assign tmp12434 = s2 ? tmp12435 : tmp12436;
  assign tmp12425 = s3 ? tmp12426 : tmp12434;
  assign tmp12440 = s1 ? tmp12422 : tmp12383;
  assign tmp12441 = s1 ? tmp12383 : tmp12416;
  assign tmp12439 = s2 ? tmp12440 : tmp12441;
  assign tmp12442 = ~(s2 ? tmp11523 : 0);
  assign tmp12438 = s3 ? tmp12439 : tmp12442;
  assign tmp12424 = s4 ? tmp12425 : tmp12438;
  assign tmp12443 = ~(s4 ? tmp11521 : tmp11528);
  assign tmp12423 = s5 ? tmp12424 : tmp12443;
  assign tmp12404 = s6 ? tmp12405 : tmp12423;
  assign tmp12448 = s1 ? tmp12418 : tmp12361;
  assign tmp12447 = s2 ? tmp12415 : tmp12448;
  assign tmp12449 = s2 ? tmp12396 : tmp12420;
  assign tmp12446 = s3 ? tmp12447 : tmp12449;
  assign tmp12445 = s4 ? tmp12406 : tmp12446;
  assign tmp12454 = s1 ? tmp12428 : tmp12408;
  assign tmp12455 = s1 ? tmp12408 : tmp11712;
  assign tmp12453 = s2 ? tmp12454 : tmp12455;
  assign tmp12457 = s1 ? tmp11704 : tmp11527;
  assign tmp12456 = s2 ? tmp12457 : tmp12436;
  assign tmp12452 = s3 ? tmp12453 : tmp12456;
  assign tmp12460 = s1 ? tmp12361 : tmp12416;
  assign tmp12459 = s2 ? tmp12440 : tmp12460;
  assign tmp12458 = s3 ? tmp12459 : tmp12442;
  assign tmp12451 = s4 ? tmp12452 : tmp12458;
  assign tmp12461 = ~(s4 ? tmp11548 : tmp11550);
  assign tmp12450 = s5 ? tmp12451 : tmp12461;
  assign tmp12444 = s6 ? tmp12445 : tmp12450;
  assign tmp12403 = s7 ? tmp12404 : tmp12444;
  assign tmp12402 = s8 ? tmp12403 : tmp12404;
  assign tmp12464 = ~(s6 ? tmp12391 : tmp12397);
  assign tmp12463 = s7 ? tmp11681 : tmp12464;
  assign tmp12471 = s1 ? tmp12361 : tmp11575;
  assign tmp12470 = s2 ? tmp11589 : tmp12471;
  assign tmp12469 = ~(s3 ? tmp12470 : tmp11612);
  assign tmp12468 = s4 ? tmp12355 : tmp12469;
  assign tmp12467 = s5 ? tmp12468 : tmp11547;
  assign tmp12466 = s6 ? tmp11598 : tmp12467;
  assign tmp12477 = s1 ? tmp12361 : tmp12408;
  assign tmp12476 = s2 ? tmp12440 : tmp12477;
  assign tmp12475 = s3 ? tmp12476 : tmp12442;
  assign tmp12474 = s4 ? tmp12452 : tmp12475;
  assign tmp12473 = s5 ? tmp12474 : tmp12461;
  assign tmp12472 = ~(s6 ? tmp12445 : tmp12473);
  assign tmp12465 = s7 ? tmp12466 : tmp12472;
  assign tmp12462 = ~(s8 ? tmp12463 : tmp12465);
  assign tmp12401 = ~(s9 ? tmp12402 : tmp12462);
  assign tmp12338 = s10 ? tmp12339 : tmp12401;
  assign tmp12481 = s7 ? tmp11531 : tmp12464;
  assign tmp12483 = ~(s6 ? tmp12445 : tmp12450);
  assign tmp12482 = s7 ? tmp12352 : tmp12483;
  assign tmp12480 = ~(s8 ? tmp12481 : tmp12482);
  assign tmp12479 = ~(s9 ? tmp12402 : tmp12480);
  assign tmp12478 = s10 ? tmp12339 : tmp12479;
  assign tmp12337 = s11 ? tmp12338 : tmp12478;
  assign tmp12494 = s1 ? 1 : tmp11494;
  assign tmp12495 = s1 ? 1 : tmp11717;
  assign tmp12493 = s2 ? tmp12494 : tmp12495;
  assign tmp12492 = s3 ? 1 : tmp12493;
  assign tmp12491 = s4 ? 1 : tmp12492;
  assign tmp12500 = ~(s1 ? 1 : tmp11717);
  assign tmp12499 = s2 ? tmp12494 : tmp12500;
  assign tmp12498 = s3 ? 1 : tmp12499;
  assign tmp12503 = s1 ? tmp11494 : tmp11717;
  assign tmp12504 = ~(s1 ? tmp11494 : 1);
  assign tmp12502 = s2 ? tmp12503 : tmp12504;
  assign tmp12501 = ~(s3 ? tmp12502 : 1);
  assign tmp12497 = s4 ? tmp12498 : tmp12501;
  assign tmp12496 = s5 ? tmp12497 : 0;
  assign tmp12490 = s6 ? tmp12491 : tmp12496;
  assign tmp12510 = s1 ? 1 : 0;
  assign tmp12509 = s2 ? tmp12510 : tmp12500;
  assign tmp12508 = s3 ? 1 : tmp12509;
  assign tmp12512 = s2 ? tmp12503 : 0;
  assign tmp12511 = ~(s3 ? tmp12512 : 1);
  assign tmp12507 = s4 ? tmp12508 : tmp12511;
  assign tmp12506 = s5 ? tmp12507 : 0;
  assign tmp12505 = s6 ? tmp12491 : tmp12506;
  assign tmp12489 = s7 ? tmp12490 : tmp12505;
  assign tmp12519 = ~(s1 ? 1 : 0);
  assign tmp12518 = s2 ? tmp12494 : tmp12519;
  assign tmp12517 = s3 ? 1 : tmp12518;
  assign tmp12521 = s2 ? tmp12096 : 0;
  assign tmp12520 = ~(s3 ? tmp12521 : 1);
  assign tmp12516 = s4 ? tmp12517 : tmp12520;
  assign tmp12515 = s5 ? tmp12516 : 0;
  assign tmp12514 = s6 ? tmp12491 : tmp12515;
  assign tmp12528 = ~(l1 ? tmp11480 : 0);
  assign tmp12527 = s0 ? 1 : tmp12528;
  assign tmp12526 = s1 ? 1 : tmp12527;
  assign tmp12525 = s2 ? 1 : tmp12526;
  assign tmp12531 = ~(s0 ? tmp11586 : 1);
  assign tmp12530 = s1 ? 1 : tmp12531;
  assign tmp12529 = s2 ? tmp12530 : tmp12495;
  assign tmp12524 = s3 ? tmp12525 : tmp12529;
  assign tmp12523 = s4 ? 1 : tmp12524;
  assign tmp12535 = s2 ? tmp12510 : tmp12519;
  assign tmp12534 = s3 ? 1 : tmp12535;
  assign tmp12533 = s4 ? tmp12534 : tmp12520;
  assign tmp12532 = s5 ? tmp12533 : 0;
  assign tmp12522 = s6 ? tmp12523 : tmp12532;
  assign tmp12513 = s7 ? tmp12514 : tmp12522;
  assign tmp12488 = s8 ? tmp12489 : tmp12513;
  assign tmp12543 = s0 ? tmp11586 : 1;
  assign tmp12542 = s1 ? tmp11586 : tmp12543;
  assign tmp12545 = s0 ? 1 : tmp11586;
  assign tmp12544 = s1 ? tmp11586 : tmp12545;
  assign tmp12541 = s2 ? tmp12542 : tmp12544;
  assign tmp12540 = s3 ? tmp11586 : tmp12541;
  assign tmp12539 = s4 ? tmp11586 : tmp12540;
  assign tmp12551 = s0 ? tmp11586 : 0;
  assign tmp12552 = ~(s0 ? 1 : tmp12528);
  assign tmp12550 = s1 ? tmp12551 : tmp12552;
  assign tmp12553 = ~(s1 ? tmp11526 : tmp11623);
  assign tmp12549 = s2 ? tmp12550 : tmp12553;
  assign tmp12555 = s1 ? tmp11632 : tmp11646;
  assign tmp12556 = s1 ? 1 : tmp11480;
  assign tmp12554 = s2 ? tmp12555 : tmp12556;
  assign tmp12548 = s3 ? tmp12549 : tmp12554;
  assign tmp12559 = s1 ? tmp11508 : tmp11480;
  assign tmp12558 = s2 ? tmp12559 : tmp11480;
  assign tmp12557 = s3 ? tmp12558 : 1;
  assign tmp12547 = s4 ? tmp12548 : tmp12557;
  assign tmp12546 = s5 ? tmp12547 : 1;
  assign tmp12538 = s6 ? tmp12539 : tmp12546;
  assign tmp12565 = s1 ? tmp12551 : tmp11586;
  assign tmp12566 = s1 ? tmp11480 : tmp11632;
  assign tmp12564 = s2 ? tmp12565 : tmp12566;
  assign tmp12567 = s2 ? tmp11665 : tmp12556;
  assign tmp12563 = s3 ? tmp12564 : tmp12567;
  assign tmp12562 = s4 ? tmp12563 : tmp12557;
  assign tmp12561 = s5 ? tmp12562 : 1;
  assign tmp12560 = s6 ? tmp12539 : tmp12561;
  assign tmp12537 = ~(s7 ? tmp12538 : tmp12560);
  assign tmp12536 = s8 ? tmp12513 : tmp12537;
  assign tmp12487 = s9 ? tmp12488 : tmp12536;
  assign tmp12570 = s7 ? tmp12538 : tmp12560;
  assign tmp12569 = s8 ? tmp12570 : tmp12538;
  assign tmp12576 = s2 ? tmp12510 : tmp12495;
  assign tmp12575 = s3 ? 1 : tmp12576;
  assign tmp12574 = s4 ? 1 : tmp12575;
  assign tmp12573 = s6 ? tmp12574 : tmp12506;
  assign tmp12581 = s1 ? tmp11586 : 1;
  assign tmp12580 = s2 ? tmp12581 : tmp12544;
  assign tmp12579 = s3 ? tmp11586 : tmp12580;
  assign tmp12578 = s4 ? tmp11586 : tmp12579;
  assign tmp12577 = ~(s6 ? tmp12578 : tmp12561);
  assign tmp12572 = s7 ? tmp12573 : tmp12577;
  assign tmp12585 = s3 ? tmp12525 : tmp12576;
  assign tmp12584 = s4 ? 1 : tmp12585;
  assign tmp12583 = s6 ? tmp12584 : tmp12532;
  assign tmp12582 = s7 ? tmp12583 : tmp12577;
  assign tmp12571 = ~(s8 ? tmp12572 : tmp12582);
  assign tmp12568 = ~(s9 ? tmp12569 : tmp12571);
  assign tmp12486 = s10 ? tmp12487 : tmp12568;
  assign tmp12590 = ~(s6 ? tmp12539 : tmp12561);
  assign tmp12589 = s7 ? tmp12505 : tmp12590;
  assign tmp12591 = s7 ? tmp12522 : tmp12590;
  assign tmp12588 = ~(s8 ? tmp12589 : tmp12591);
  assign tmp12587 = ~(s9 ? tmp12569 : tmp12588);
  assign tmp12586 = s10 ? tmp12487 : tmp12587;
  assign tmp12485 = s11 ? tmp12486 : tmp12586;
  assign tmp12484 = s12 ? 1 : tmp12485;
  assign tmp12336 = s13 ? tmp12337 : tmp12484;
  assign tmp12604 = ~(s1 ? tmp11634 : tmp11623);
  assign tmp12603 = s2 ? tmp11844 : tmp12604;
  assign tmp12605 = s2 ? tmp11870 : tmp11646;
  assign tmp12602 = s3 ? tmp12603 : tmp12605;
  assign tmp12607 = s2 ? tmp12555 : tmp11852;
  assign tmp12606 = s3 ? tmp12607 : tmp12197;
  assign tmp12601 = s4 ? tmp12602 : tmp12606;
  assign tmp12600 = s5 ? tmp12601 : 0;
  assign tmp12599 = s6 ? tmp11632 : tmp12600;
  assign tmp12612 = s2 ? tmp11835 : tmp11632;
  assign tmp12616 = ~(l2 ? tmp11479 : 1);
  assign tmp12615 = l1 ? 1 : tmp12616;
  assign tmp12617 = s0 ? tmp12615 : 0;
  assign tmp12614 = s1 ? tmp12615 : tmp12617;
  assign tmp12613 = s2 ? tmp12614 : tmp11646;
  assign tmp12611 = s3 ? tmp12612 : tmp12613;
  assign tmp12619 = s2 ? tmp12555 : tmp11632;
  assign tmp12618 = s3 ? tmp12619 : tmp11717;
  assign tmp12610 = s4 ? tmp12611 : tmp12618;
  assign tmp12609 = s5 ? tmp12610 : 0;
  assign tmp12608 = s6 ? tmp11632 : tmp12609;
  assign tmp12598 = ~(s7 ? tmp12599 : tmp12608);
  assign tmp12597 = s8 ? 1 : tmp12598;
  assign tmp12596 = s9 ? tmp12597 : tmp12598;
  assign tmp12622 = s7 ? tmp12599 : tmp12608;
  assign tmp12621 = s8 ? tmp12622 : tmp12599;
  assign tmp12630 = s1 ? tmp12615 : 0;
  assign tmp12629 = s2 ? tmp12630 : tmp11646;
  assign tmp12628 = s3 ? tmp12612 : tmp12629;
  assign tmp12627 = s4 ? tmp12628 : tmp12618;
  assign tmp12626 = s5 ? tmp12627 : 0;
  assign tmp12625 = ~(s6 ? tmp11632 : tmp12626);
  assign tmp12624 = s7 ? 1 : tmp12625;
  assign tmp12623 = ~(s8 ? tmp12624 : tmp12625);
  assign tmp12620 = ~(s9 ? tmp12621 : tmp12623);
  assign tmp12595 = s10 ? tmp12596 : tmp12620;
  assign tmp12635 = ~(s6 ? tmp11632 : tmp12609);
  assign tmp12634 = s7 ? 1 : tmp12635;
  assign tmp12633 = ~(s8 ? tmp12634 : tmp12635);
  assign tmp12632 = ~(s9 ? tmp12621 : tmp12633);
  assign tmp12631 = s10 ? tmp12596 : tmp12632;
  assign tmp12594 = s11 ? tmp12595 : tmp12631;
  assign tmp12593 = s12 ? tmp12594 : 0;
  assign tmp12644 = ~(l2 ? tmp11479 : 0);
  assign tmp12643 = l1 ? 1 : tmp12644;
  assign tmp12647 = s0 ? tmp12643 : 0;
  assign tmp12646 = s2 ? tmp12643 : tmp12647;
  assign tmp12650 = s0 ? 1 : tmp12643;
  assign tmp12649 = s1 ? tmp12643 : tmp12650;
  assign tmp12648 = s2 ? tmp11779 : tmp12649;
  assign tmp12645 = s3 ? tmp12646 : tmp12648;
  assign tmp12642 = s4 ? tmp12643 : tmp12645;
  assign tmp12656 = s0 ? tmp12643 : 1;
  assign tmp12655 = s1 ? 1 : tmp12656;
  assign tmp12654 = s2 ? tmp12643 : tmp12655;
  assign tmp12653 = s3 ? tmp12643 : tmp12654;
  assign tmp12659 = s1 ? tmp12650 : tmp11646;
  assign tmp12660 = s1 ? tmp11646 : tmp12643;
  assign tmp12658 = s2 ? tmp12659 : tmp12660;
  assign tmp12662 = s1 ? tmp12656 : 1;
  assign tmp12661 = s2 ? tmp12662 : 1;
  assign tmp12657 = s3 ? tmp12658 : tmp12661;
  assign tmp12652 = s4 ? tmp12653 : tmp12657;
  assign tmp12665 = s2 ? tmp12662 : tmp12650;
  assign tmp12664 = s3 ? tmp12665 : 1;
  assign tmp12668 = s1 ? tmp12650 : tmp12656;
  assign tmp12667 = s2 ? 1 : tmp12668;
  assign tmp12666 = s3 ? tmp12667 : 1;
  assign tmp12663 = s4 ? tmp12664 : tmp12666;
  assign tmp12651 = s5 ? tmp12652 : tmp12663;
  assign tmp12641 = s6 ? tmp12642 : tmp12651;
  assign tmp12673 = s1 ? tmp12647 : tmp11768;
  assign tmp12672 = s2 ? tmp12643 : tmp12673;
  assign tmp12674 = s2 ? tmp11800 : tmp12649;
  assign tmp12671 = s3 ? tmp12672 : tmp12674;
  assign tmp12670 = s4 ? tmp12643 : tmp12671;
  assign tmp12678 = s2 ? tmp12659 : tmp12643;
  assign tmp12677 = s3 ? tmp12678 : tmp12661;
  assign tmp12676 = s4 ? tmp12653 : tmp12677;
  assign tmp12682 = s1 ? tmp12643 : 1;
  assign tmp12681 = s2 ? tmp12662 : tmp12682;
  assign tmp12680 = s3 ? tmp12681 : 1;
  assign tmp12684 = s2 ? 1 : tmp12643;
  assign tmp12683 = s3 ? tmp12684 : 1;
  assign tmp12679 = s4 ? tmp12680 : tmp12683;
  assign tmp12675 = s5 ? tmp12676 : tmp12679;
  assign tmp12669 = s6 ? tmp12670 : tmp12675;
  assign tmp12640 = s7 ? tmp12641 : tmp12669;
  assign tmp12690 = s2 ? tmp11768 : tmp11777;
  assign tmp12689 = s3 ? tmp12690 : tmp11778;
  assign tmp12688 = s4 ? tmp11768 : tmp12689;
  assign tmp12694 = s2 ? tmp11768 : tmp12184;
  assign tmp12693 = s3 ? tmp11768 : tmp12694;
  assign tmp12697 = s1 ? tmp11646 : tmp11768;
  assign tmp12696 = s2 ? tmp11797 : tmp12697;
  assign tmp12698 = s2 ? tmp11804 : 1;
  assign tmp12695 = s3 ? tmp12696 : tmp12698;
  assign tmp12692 = s4 ? tmp12693 : tmp12695;
  assign tmp12691 = s5 ? tmp12692 : tmp11801;
  assign tmp12687 = s6 ? tmp12688 : tmp12691;
  assign tmp12702 = s2 ? tmp11768 : tmp11813;
  assign tmp12701 = s3 ? tmp12702 : tmp11814;
  assign tmp12700 = s4 ? tmp11768 : tmp12701;
  assign tmp12705 = s3 ? tmp11823 : tmp12698;
  assign tmp12704 = s4 ? tmp12693 : tmp12705;
  assign tmp12709 = s1 ? tmp11768 : tmp11805;
  assign tmp12708 = s2 ? 1 : tmp12709;
  assign tmp12707 = s3 ? tmp12708 : 1;
  assign tmp12706 = s4 ? tmp11802 : tmp12707;
  assign tmp12703 = s5 ? tmp12704 : tmp12706;
  assign tmp12699 = s6 ? tmp12700 : tmp12703;
  assign tmp12686 = s7 ? tmp12687 : tmp12699;
  assign tmp12685 = s8 ? tmp12640 : tmp12686;
  assign tmp12639 = s9 ? tmp12640 : tmp12685;
  assign tmp12711 = s8 ? tmp12640 : tmp12641;
  assign tmp12717 = s2 ? tmp11704 : tmp11749;
  assign tmp12716 = s3 ? tmp12717 : tmp11750;
  assign tmp12715 = s4 ? tmp11704 : tmp12716;
  assign tmp12720 = s3 ? tmp11704 : tmp11756;
  assign tmp12719 = s4 ? tmp12720 : tmp11758;
  assign tmp12718 = s5 ? tmp12719 : tmp11908;
  assign tmp12714 = s6 ? tmp12715 : tmp12718;
  assign tmp12723 = s4 ? tmp11802 : tmp11904;
  assign tmp12722 = s5 ? tmp12704 : tmp12723;
  assign tmp12721 = s6 ? tmp12700 : tmp12722;
  assign tmp12713 = s7 ? tmp12714 : tmp12721;
  assign tmp12712 = s8 ? tmp12713 : tmp12669;
  assign tmp12710 = s9 ? tmp12711 : tmp12712;
  assign tmp12638 = s10 ? tmp12639 : tmp12710;
  assign tmp12727 = s7 ? tmp12714 : tmp12699;
  assign tmp12726 = s8 ? tmp12727 : tmp12669;
  assign tmp12725 = s9 ? tmp12711 : tmp12726;
  assign tmp12724 = s10 ? tmp12639 : tmp12725;
  assign tmp12637 = s11 ? tmp12638 : tmp12724;
  assign tmp12636 = ~(s12 ? tmp12637 : 1);
  assign tmp12592 = s13 ? tmp12593 : tmp12636;
  assign tmp12335 = s14 ? tmp12336 : tmp12592;
  assign tmp12739 = s2 ? tmp12063 : tmp12066;
  assign tmp12738 = s3 ? tmp12062 : tmp12739;
  assign tmp12737 = s4 ? tmp12738 : tmp12068;
  assign tmp12743 = s2 ? tmp12093 : tmp12063;
  assign tmp12742 = s3 ? tmp12743 : tmp12095;
  assign tmp12741 = s4 ? tmp12742 : tmp12098;
  assign tmp12740 = s5 ? tmp12075 : tmp12741;
  assign tmp12736 = s6 ? tmp12737 : tmp12740;
  assign tmp12745 = s4 ? tmp12738 : tmp12108;
  assign tmp12750 = s1 ? tmp12063 : 1;
  assign tmp12749 = s2 ? tmp12080 : tmp12750;
  assign tmp12748 = s3 ? tmp12749 : tmp12123;
  assign tmp12747 = s4 ? tmp12748 : tmp12063;
  assign tmp12746 = s5 ? tmp12112 : tmp12747;
  assign tmp12744 = s6 ? tmp12745 : tmp12746;
  assign tmp12735 = s7 ? tmp12736 : tmp12744;
  assign tmp12734 = s8 ? tmp12058 : tmp12735;
  assign tmp12733 = s9 ? tmp12058 : tmp12734;
  assign tmp12754 = s6 ? tmp12737 : tmp12074;
  assign tmp12755 = s6 ? tmp12745 : tmp12111;
  assign tmp12753 = s7 ? tmp12754 : tmp12755;
  assign tmp12752 = s8 ? tmp12753 : tmp12754;
  assign tmp12757 = s7 ? tmp12158 : tmp12744;
  assign tmp12758 = s6 ? tmp12745 : tmp12159;
  assign tmp12756 = s8 ? tmp12757 : tmp12758;
  assign tmp12751 = s9 ? tmp12752 : tmp12756;
  assign tmp12732 = s10 ? tmp12733 : tmp12751;
  assign tmp12762 = s7 ? tmp12106 : tmp12744;
  assign tmp12761 = s8 ? tmp12762 : tmp12755;
  assign tmp12760 = s9 ? tmp12752 : tmp12761;
  assign tmp12759 = s10 ? tmp12733 : tmp12760;
  assign tmp12731 = s11 ? tmp12732 : tmp12759;
  assign tmp12730 = s12 ? 1 : tmp12731;
  assign tmp12729 = ~(s13 ? tmp12730 : tmp12166);
  assign tmp12728 = s14 ? tmp11915 : tmp12729;
  assign tmp12334 = s15 ? tmp12335 : tmp12728;
  assign tmp11465 = s16 ? tmp11466 : tmp12334;
  assign tmp12770 = s8 ? tmp12341 : tmp11615;
  assign tmp12769 = s9 ? tmp12340 : tmp12770;
  assign tmp12773 = s7 ? tmp12466 : tmp11674;
  assign tmp12772 = s8 ? tmp11680 : tmp12773;
  assign tmp12771 = s9 ? tmp11672 : tmp12772;
  assign tmp12768 = s10 ? tmp12769 : tmp12771;
  assign tmp12777 = s7 ? tmp12352 : tmp11674;
  assign tmp12776 = s8 ? tmp11691 : tmp12777;
  assign tmp12775 = s9 ? tmp11672 : tmp12776;
  assign tmp12774 = s10 ? tmp12769 : tmp12775;
  assign tmp12767 = s11 ? tmp12768 : tmp12774;
  assign tmp12783 = s7 ? tmp12490 : tmp12573;
  assign tmp12782 = s8 ? tmp12513 : tmp12783;
  assign tmp12781 = s9 ? tmp12488 : tmp12782;
  assign tmp12785 = s8 ? tmp12783 : tmp12490;
  assign tmp12787 = s7 ? tmp12583 : tmp12573;
  assign tmp12786 = s8 ? tmp12573 : tmp12787;
  assign tmp12784 = s9 ? tmp12785 : tmp12786;
  assign tmp12780 = s10 ? tmp12781 : tmp12784;
  assign tmp12791 = s7 ? tmp12505 : tmp12573;
  assign tmp12792 = s7 ? tmp12522 : tmp12573;
  assign tmp12790 = s8 ? tmp12791 : tmp12792;
  assign tmp12789 = s9 ? tmp12785 : tmp12790;
  assign tmp12788 = s10 ? tmp12781 : tmp12789;
  assign tmp12779 = s11 ? tmp12780 : tmp12788;
  assign tmp12778 = s12 ? 1 : tmp12779;
  assign tmp12766 = s13 ? tmp12767 : tmp12778;
  assign tmp12798 = ~(s8 ? tmp12622 : 0);
  assign tmp12797 = s9 ? tmp12597 : tmp12798;
  assign tmp12802 = s6 ? tmp11632 : tmp12626;
  assign tmp12801 = ~(s7 ? tmp12802 : 0);
  assign tmp12800 = s8 ? 1 : tmp12801;
  assign tmp12799 = s9 ? 1 : tmp12800;
  assign tmp12796 = s10 ? tmp12797 : tmp12799;
  assign tmp12806 = ~(s7 ? tmp12608 : 0);
  assign tmp12805 = s8 ? 1 : tmp12806;
  assign tmp12804 = s9 ? 1 : tmp12805;
  assign tmp12803 = s10 ? tmp12797 : tmp12804;
  assign tmp12795 = s11 ? tmp12796 : tmp12803;
  assign tmp12794 = s12 ? tmp12795 : 0;
  assign tmp12817 = s1 ? tmp12643 : tmp12656;
  assign tmp12816 = s2 ? 1 : tmp12817;
  assign tmp12815 = s3 ? tmp12816 : 1;
  assign tmp12814 = s4 ? tmp12664 : tmp12815;
  assign tmp12813 = s5 ? tmp12676 : tmp12814;
  assign tmp12812 = s6 ? tmp12670 : tmp12813;
  assign tmp12811 = s7 ? tmp12641 : tmp12812;
  assign tmp12821 = s4 ? tmp11632 : tmp11836;
  assign tmp12826 = s1 ? 1 : tmp11646;
  assign tmp12825 = s2 ? tmp11632 : tmp12826;
  assign tmp12824 = s3 ? tmp11632 : tmp12825;
  assign tmp12827 = s3 ? tmp11850 : tmp12388;
  assign tmp12823 = s4 ? tmp12824 : tmp12827;
  assign tmp12830 = s2 ? tmp11645 : tmp11648;
  assign tmp12829 = s3 ? tmp12830 : 1;
  assign tmp12832 = s2 ? 1 : tmp11851;
  assign tmp12831 = s3 ? tmp12832 : 1;
  assign tmp12828 = s4 ? tmp12829 : tmp12831;
  assign tmp12822 = s5 ? tmp12823 : tmp12828;
  assign tmp12820 = s6 ? tmp12821 : tmp12822;
  assign tmp12834 = s4 ? tmp11632 : tmp11864;
  assign tmp12837 = s3 ? tmp11874 : tmp12388;
  assign tmp12836 = s4 ? tmp12824 : tmp12837;
  assign tmp12840 = s2 ? 1 : tmp11665;
  assign tmp12839 = s3 ? tmp12840 : 1;
  assign tmp12838 = s4 ? tmp11667 : tmp12839;
  assign tmp12835 = s5 ? tmp12836 : tmp12838;
  assign tmp12833 = s6 ? tmp12834 : tmp12835;
  assign tmp12819 = s7 ? tmp12820 : tmp12833;
  assign tmp12818 = s8 ? tmp12811 : tmp12819;
  assign tmp12810 = s9 ? tmp12811 : tmp12818;
  assign tmp12847 = s2 ? tmp11704 : tmp11708;
  assign tmp12846 = s3 ? tmp12847 : tmp11715;
  assign tmp12845 = s4 ? tmp11704 : tmp12846;
  assign tmp12852 = s1 ? tmp11646 : tmp11704;
  assign tmp12851 = s2 ? tmp11735 : tmp12852;
  assign tmp12850 = s3 ? tmp12851 : tmp11737;
  assign tmp12849 = s4 ? tmp12720 : tmp12850;
  assign tmp12848 = s5 ? tmp12849 : tmp11739;
  assign tmp12844 = s6 ? tmp12845 : tmp12848;
  assign tmp12854 = s5 ? tmp12719 : tmp11884;
  assign tmp12853 = s6 ? tmp12715 : tmp12854;
  assign tmp12843 = s7 ? tmp12844 : tmp12853;
  assign tmp12842 = s8 ? tmp12843 : tmp12844;
  assign tmp12858 = s4 ? tmp12664 : tmp12683;
  assign tmp12857 = s5 ? tmp12676 : tmp12858;
  assign tmp12856 = s6 ? tmp12670 : tmp12857;
  assign tmp12855 = s7 ? tmp12856 : tmp12714;
  assign tmp12841 = s9 ? tmp12842 : tmp12855;
  assign tmp12809 = s10 ? tmp12810 : tmp12841;
  assign tmp12861 = s7 ? tmp12812 : tmp12853;
  assign tmp12860 = s9 ? tmp12842 : tmp12861;
  assign tmp12859 = s10 ? tmp12810 : tmp12860;
  assign tmp12808 = s11 ? tmp12809 : tmp12859;
  assign tmp12807 = ~(s12 ? tmp12808 : 1);
  assign tmp12793 = s13 ? tmp12794 : tmp12807;
  assign tmp12765 = s14 ? tmp12766 : tmp12793;
  assign tmp12868 = s8 ? tmp12058 : tmp12145;
  assign tmp12867 = s9 ? tmp12058 : tmp12868;
  assign tmp12871 = s7 ? tmp12158 : tmp12152;
  assign tmp12870 = s8 ? tmp12157 : tmp12871;
  assign tmp12869 = s9 ? tmp12150 : tmp12870;
  assign tmp12866 = s10 ? tmp12867 : tmp12869;
  assign tmp12875 = s7 ? tmp12106 : tmp12152;
  assign tmp12874 = s8 ? tmp12165 : tmp12875;
  assign tmp12873 = s9 ? tmp12150 : tmp12874;
  assign tmp12872 = s10 ? tmp12867 : tmp12873;
  assign tmp12865 = s11 ? tmp12866 : tmp12872;
  assign tmp12864 = s12 ? 1 : tmp12865;
  assign tmp12863 = ~(s13 ? tmp12864 : tmp12166);
  assign tmp12862 = s14 ? tmp11915 : tmp12863;
  assign tmp12764 = s15 ? tmp12765 : tmp12862;
  assign tmp12883 = s8 ? tmp12811 : tmp12686;
  assign tmp12882 = s9 ? tmp12811 : tmp12883;
  assign tmp12885 = s8 ? tmp12811 : tmp12641;
  assign tmp12884 = s9 ? tmp12885 : tmp12856;
  assign tmp12881 = s10 ? tmp12882 : tmp12884;
  assign tmp12887 = s9 ? tmp12885 : tmp12812;
  assign tmp12886 = s10 ? tmp12882 : tmp12887;
  assign tmp12880 = s11 ? tmp12881 : tmp12886;
  assign tmp12879 = ~(s12 ? tmp12880 : 1);
  assign tmp12878 = s13 ? tmp12593 : tmp12879;
  assign tmp12877 = s14 ? tmp12336 : tmp12878;
  assign tmp12876 = s15 ? tmp12877 : tmp12728;
  assign tmp12763 = s16 ? tmp12764 : tmp12876;
  assign tmp11464 = s17 ? tmp11465 : tmp12763;
  assign l3__1 = tmp11464;

  assign tmp12903 = l2 ? 1 : 0;
  assign tmp12905 = l1 ? 1 : 0;
  assign tmp12906 = ~(l2 ? 1 : 0);
  assign tmp12904 = ~(s0 ? tmp12905 : tmp12906);
  assign tmp12902 = s1 ? tmp12903 : tmp12904;
  assign tmp12909 = s0 ? tmp12903 : 0;
  assign tmp12908 = s1 ? tmp12909 : tmp12903;
  assign tmp12907 = s2 ? tmp12903 : tmp12908;
  assign tmp12901 = s3 ? tmp12902 : tmp12907;
  assign tmp12913 = ~(s0 ? tmp12905 : 1);
  assign tmp12912 = s1 ? tmp12909 : tmp12913;
  assign tmp12911 = s2 ? tmp12908 : tmp12912;
  assign tmp12916 = s0 ? 1 : 0;
  assign tmp12915 = s1 ? tmp12905 : tmp12916;
  assign tmp12918 = s0 ? 1 : tmp12903;
  assign tmp12917 = ~(s1 ? tmp12903 : tmp12918);
  assign tmp12914 = ~(s2 ? tmp12915 : tmp12917);
  assign tmp12910 = s3 ? tmp12911 : tmp12914;
  assign tmp12900 = s4 ? tmp12901 : tmp12910;
  assign tmp12923 = s1 ? tmp12909 : 0;
  assign tmp12925 = s0 ? 1 : tmp12906;
  assign tmp12924 = ~(s1 ? tmp12925 : tmp12906);
  assign tmp12922 = s2 ? tmp12923 : tmp12924;
  assign tmp12927 = s1 ? 1 : tmp12903;
  assign tmp12926 = s2 ? tmp12903 : tmp12927;
  assign tmp12921 = s3 ? tmp12922 : tmp12926;
  assign tmp12931 = ~(l1 ? 1 : 0);
  assign tmp12930 = s1 ? tmp12918 : tmp12931;
  assign tmp12933 = ~(s0 ? tmp12903 : 0);
  assign tmp12932 = ~(s1 ? tmp12905 : tmp12933);
  assign tmp12929 = s2 ? tmp12930 : tmp12932;
  assign tmp12934 = s2 ? tmp12902 : 1;
  assign tmp12928 = s3 ? tmp12929 : tmp12934;
  assign tmp12920 = s4 ? tmp12921 : tmp12928;
  assign tmp12939 = s0 ? tmp12903 : 1;
  assign tmp12938 = s1 ? tmp12939 : 1;
  assign tmp12940 = s1 ? tmp12916 : 0;
  assign tmp12937 = s2 ? tmp12938 : tmp12940;
  assign tmp12942 = ~(s1 ? 1 : tmp12918);
  assign tmp12941 = ~(s2 ? tmp12940 : tmp12942);
  assign tmp12936 = s3 ? tmp12937 : tmp12941;
  assign tmp12945 = s1 ? tmp12918 : 0;
  assign tmp12944 = s2 ? tmp12938 : tmp12945;
  assign tmp12947 = s1 ? 1 : tmp12918;
  assign tmp12948 = s1 ? tmp12918 : 1;
  assign tmp12946 = s2 ? tmp12947 : tmp12948;
  assign tmp12943 = s3 ? tmp12944 : tmp12946;
  assign tmp12935 = s4 ? tmp12936 : tmp12943;
  assign tmp12919 = s5 ? tmp12920 : tmp12935;
  assign tmp12899 = s6 ? tmp12900 : tmp12919;
  assign tmp12953 = s1 ? tmp12909 : tmp12931;
  assign tmp12952 = s2 ? tmp12908 : tmp12953;
  assign tmp12955 = s1 ? tmp12905 : 0;
  assign tmp12954 = ~(s2 ? tmp12955 : tmp12917);
  assign tmp12951 = s3 ? tmp12952 : tmp12954;
  assign tmp12950 = s4 ? tmp12901 : tmp12951;
  assign tmp12959 = s2 ? tmp12923 : tmp12903;
  assign tmp12958 = s3 ? tmp12959 : tmp12926;
  assign tmp12962 = ~(s1 ? tmp12905 : tmp12906);
  assign tmp12961 = s2 ? tmp12930 : tmp12962;
  assign tmp12960 = s3 ? tmp12961 : tmp12934;
  assign tmp12957 = s4 ? tmp12958 : tmp12960;
  assign tmp12965 = s2 ? tmp12938 : 0;
  assign tmp12966 = s2 ? 1 : tmp12927;
  assign tmp12964 = s3 ? tmp12965 : tmp12966;
  assign tmp12968 = s2 ? 1 : tmp12903;
  assign tmp12967 = s3 ? tmp12968 : tmp12927;
  assign tmp12963 = s4 ? tmp12964 : tmp12967;
  assign tmp12956 = s5 ? tmp12957 : tmp12963;
  assign tmp12949 = s6 ? tmp12950 : tmp12956;
  assign tmp12898 = s7 ? tmp12899 : tmp12949;
  assign tmp12975 = ~(s1 ? tmp12925 : tmp12933);
  assign tmp12974 = s2 ? tmp12923 : tmp12975;
  assign tmp12977 = ~(s1 ? 1 : tmp12903);
  assign tmp12976 = ~(s2 ? tmp12925 : tmp12977);
  assign tmp12973 = s3 ? tmp12974 : tmp12976;
  assign tmp12972 = s4 ? tmp12973 : tmp12928;
  assign tmp12971 = s5 ? tmp12972 : tmp12935;
  assign tmp12970 = s6 ? tmp12900 : tmp12971;
  assign tmp12983 = s1 ? tmp12903 : tmp12909;
  assign tmp12982 = s2 ? tmp12923 : tmp12983;
  assign tmp12981 = s3 ? tmp12982 : tmp12926;
  assign tmp12985 = s2 ? tmp12930 : tmp12903;
  assign tmp12986 = s2 ? tmp12903 : 1;
  assign tmp12984 = s3 ? tmp12985 : tmp12986;
  assign tmp12980 = s4 ? tmp12981 : tmp12984;
  assign tmp12979 = s5 ? tmp12980 : tmp12963;
  assign tmp12978 = s6 ? tmp12950 : tmp12979;
  assign tmp12969 = s7 ? tmp12970 : tmp12978;
  assign tmp12897 = s8 ? tmp12898 : tmp12969;
  assign tmp12994 = s0 ? tmp12905 : 1;
  assign tmp12993 = s1 ? tmp12994 : tmp12905;
  assign tmp12992 = s2 ? tmp12905 : tmp12993;
  assign tmp12991 = s3 ? tmp12905 : tmp12992;
  assign tmp12996 = s2 ? tmp12905 : tmp12994;
  assign tmp12999 = ~(s0 ? 1 : tmp12931);
  assign tmp12998 = s1 ? tmp12905 : tmp12999;
  assign tmp12997 = s2 ? tmp12915 : tmp12998;
  assign tmp12995 = s3 ? tmp12996 : tmp12997;
  assign tmp12990 = s4 ? tmp12991 : tmp12995;
  assign tmp13004 = s1 ? tmp12994 : 1;
  assign tmp13006 = s0 ? 1 : tmp12905;
  assign tmp13005 = s1 ? tmp13006 : tmp12905;
  assign tmp13003 = s2 ? tmp13004 : tmp13005;
  assign tmp13008 = ~(s1 ? 1 : tmp12931);
  assign tmp13007 = s2 ? tmp12905 : tmp13008;
  assign tmp13002 = s3 ? tmp13003 : tmp13007;
  assign tmp13012 = s0 ? 1 : tmp12931;
  assign tmp13011 = s1 ? tmp13012 : tmp12931;
  assign tmp13010 = s2 ? tmp13011 : tmp12931;
  assign tmp13013 = ~(s2 ? tmp12905 : 0);
  assign tmp13009 = ~(s3 ? tmp13010 : tmp13013);
  assign tmp13001 = s4 ? tmp13002 : tmp13009;
  assign tmp13018 = s0 ? tmp12905 : 0;
  assign tmp13017 = s1 ? tmp13018 : 0;
  assign tmp13019 = ~(s1 ? tmp12916 : 0);
  assign tmp13016 = s2 ? tmp13017 : tmp13019;
  assign tmp13021 = ~(s1 ? 1 : tmp13012);
  assign tmp13020 = s2 ? tmp12940 : tmp13021;
  assign tmp13015 = s3 ? tmp13016 : tmp13020;
  assign tmp13024 = ~(s1 ? tmp13012 : 0);
  assign tmp13023 = s2 ? tmp13017 : tmp13024;
  assign tmp13026 = s1 ? 1 : tmp13012;
  assign tmp13027 = s1 ? tmp13012 : 1;
  assign tmp13025 = ~(s2 ? tmp13026 : tmp13027);
  assign tmp13022 = s3 ? tmp13023 : tmp13025;
  assign tmp13014 = s4 ? tmp13015 : tmp13022;
  assign tmp13000 = s5 ? tmp13001 : tmp13014;
  assign tmp12989 = s6 ? tmp12990 : tmp13000;
  assign tmp13031 = s2 ? tmp12955 : tmp12998;
  assign tmp13030 = s3 ? tmp12992 : tmp13031;
  assign tmp13029 = s4 ? tmp12991 : tmp13030;
  assign tmp13035 = s2 ? tmp13004 : tmp12905;
  assign tmp13034 = s3 ? tmp13035 : tmp13007;
  assign tmp13033 = s4 ? tmp13034 : tmp13009;
  assign tmp13038 = s2 ? tmp13017 : 1;
  assign tmp13040 = s1 ? 1 : tmp12931;
  assign tmp13039 = ~(s2 ? 1 : tmp13040);
  assign tmp13037 = s3 ? tmp13038 : tmp13039;
  assign tmp13042 = s2 ? 1 : tmp12931;
  assign tmp13041 = ~(s3 ? tmp13042 : tmp13040);
  assign tmp13036 = s4 ? tmp13037 : tmp13041;
  assign tmp13032 = s5 ? tmp13033 : tmp13036;
  assign tmp13028 = s6 ? tmp13029 : tmp13032;
  assign tmp12988 = ~(s7 ? tmp12989 : tmp13028);
  assign tmp12987 = s8 ? tmp12969 : tmp12988;
  assign tmp12896 = s9 ? tmp12897 : tmp12987;
  assign tmp13048 = s4 ? tmp12958 : tmp12984;
  assign tmp13047 = s5 ? tmp13048 : tmp12963;
  assign tmp13046 = s6 ? tmp12950 : tmp13047;
  assign tmp13045 = s7 ? tmp12899 : tmp13046;
  assign tmp13044 = s8 ? tmp13045 : tmp12899;
  assign tmp13054 = s3 ? tmp12961 : tmp12986;
  assign tmp13053 = s4 ? tmp12958 : tmp13054;
  assign tmp13052 = s5 ? tmp13053 : tmp12963;
  assign tmp13051 = s6 ? tmp12950 : tmp13052;
  assign tmp13055 = ~(s6 ? tmp13029 : tmp13032);
  assign tmp13050 = s7 ? tmp13051 : tmp13055;
  assign tmp13056 = s7 ? tmp12978 : tmp13046;
  assign tmp13049 = s8 ? tmp13050 : tmp13056;
  assign tmp13043 = s9 ? tmp13044 : tmp13049;
  assign tmp12895 = s10 ? tmp12896 : tmp13043;
  assign tmp13060 = s7 ? tmp12949 : tmp13055;
  assign tmp13059 = s8 ? tmp13060 : tmp13056;
  assign tmp13058 = s9 ? tmp13044 : tmp13059;
  assign tmp13057 = s10 ? tmp12896 : tmp13058;
  assign tmp12894 = ~(s11 ? tmp12895 : tmp13057);
  assign tmp12893 = s12 ? 1 : tmp12894;
  assign tmp13071 = l1 ? tmp12903 : 0;
  assign tmp13073 = ~(l1 ? tmp12903 : 0);
  assign tmp13072 = ~(s0 ? 1 : tmp13073);
  assign tmp13070 = s1 ? tmp13071 : tmp13072;
  assign tmp13076 = s0 ? tmp13071 : 0;
  assign tmp13075 = s1 ? tmp13076 : tmp13071;
  assign tmp13074 = s2 ? tmp13071 : tmp13075;
  assign tmp13069 = s3 ? tmp13070 : tmp13074;
  assign tmp13079 = s1 ? tmp13076 : 0;
  assign tmp13078 = s2 ? tmp13075 : tmp13079;
  assign tmp13081 = s1 ? 1 : tmp12916;
  assign tmp13083 = s0 ? 1 : tmp13071;
  assign tmp13082 = ~(s1 ? tmp13071 : tmp13083);
  assign tmp13080 = ~(s2 ? tmp13081 : tmp13082);
  assign tmp13077 = s3 ? tmp13078 : tmp13080;
  assign tmp13068 = s4 ? tmp13069 : tmp13077;
  assign tmp13088 = s1 ? tmp13076 : tmp13072;
  assign tmp13090 = s0 ? 1 : tmp13073;
  assign tmp13091 = ~(s0 ? tmp13071 : 0);
  assign tmp13089 = ~(s1 ? tmp13090 : tmp13091);
  assign tmp13087 = s2 ? tmp13088 : tmp13089;
  assign tmp13093 = ~(s1 ? 1 : tmp13071);
  assign tmp13092 = ~(s2 ? tmp13090 : tmp13093);
  assign tmp13086 = s3 ? tmp13087 : tmp13092;
  assign tmp13096 = s1 ? tmp13083 : 0;
  assign tmp13097 = ~(s1 ? 1 : tmp13091);
  assign tmp13095 = s2 ? tmp13096 : tmp13097;
  assign tmp13100 = ~(s0 ? 1 : tmp12906);
  assign tmp13099 = s1 ? tmp13071 : tmp13100;
  assign tmp13098 = s2 ? tmp13099 : 1;
  assign tmp13094 = s3 ? tmp13095 : tmp13098;
  assign tmp13085 = s4 ? tmp13086 : tmp13094;
  assign tmp13105 = s0 ? tmp13071 : 1;
  assign tmp13104 = s1 ? tmp13105 : 1;
  assign tmp13103 = s2 ? tmp13104 : tmp13071;
  assign tmp13106 = s2 ? tmp12938 : tmp12947;
  assign tmp13102 = s3 ? tmp13103 : tmp13106;
  assign tmp13109 = s1 ? tmp13083 : tmp13071;
  assign tmp13108 = s2 ? tmp12903 : tmp13109;
  assign tmp13107 = s3 ? tmp13108 : tmp12946;
  assign tmp13101 = s4 ? tmp13102 : tmp13107;
  assign tmp13084 = s5 ? tmp13085 : tmp13101;
  assign tmp13067 = s6 ? tmp13068 : tmp13084;
  assign tmp13114 = s1 ? 1 : 0;
  assign tmp13113 = ~(s2 ? tmp13114 : tmp13082);
  assign tmp13112 = s3 ? tmp13078 : tmp13113;
  assign tmp13111 = s4 ? tmp13069 : tmp13112;
  assign tmp13119 = s1 ? tmp13071 : tmp13076;
  assign tmp13118 = s2 ? tmp13075 : tmp13119;
  assign tmp13121 = s1 ? 1 : tmp13071;
  assign tmp13120 = s2 ? tmp13071 : tmp13121;
  assign tmp13117 = s3 ? tmp13118 : tmp13120;
  assign tmp13123 = s2 ? tmp13096 : tmp13071;
  assign tmp13125 = s1 ? tmp13071 : tmp12903;
  assign tmp13124 = s2 ? tmp13125 : 1;
  assign tmp13122 = s3 ? tmp13123 : tmp13124;
  assign tmp13116 = s4 ? tmp13117 : tmp13122;
  assign tmp13128 = s2 ? tmp13104 : tmp12927;
  assign tmp13127 = s3 ? tmp13103 : tmp13128;
  assign tmp13130 = s2 ? 1 : tmp13071;
  assign tmp13129 = s3 ? tmp13130 : tmp12903;
  assign tmp13126 = s4 ? tmp13127 : tmp13129;
  assign tmp13115 = s5 ? tmp13116 : tmp13126;
  assign tmp13110 = s6 ? tmp13111 : tmp13115;
  assign tmp13066 = s7 ? tmp13067 : tmp13110;
  assign tmp13137 = ~(l3 ? 1 : 0);
  assign tmp13136 = l1 ? tmp12903 : tmp13137;
  assign tmp13140 = l3 ? 1 : 0;
  assign tmp13139 = l1 ? 1 : tmp13140;
  assign tmp13141 = ~(l1 ? tmp12903 : tmp13137);
  assign tmp13138 = ~(s0 ? tmp13139 : tmp13141);
  assign tmp13135 = s1 ? tmp13136 : tmp13138;
  assign tmp13144 = s0 ? tmp13136 : tmp13137;
  assign tmp13143 = s1 ? tmp13144 : tmp13136;
  assign tmp13142 = s2 ? tmp13136 : tmp13143;
  assign tmp13134 = s3 ? tmp13135 : tmp13142;
  assign tmp13148 = s0 ? tmp13136 : 0;
  assign tmp13147 = s1 ? tmp13148 : tmp13136;
  assign tmp13150 = ~(s0 ? tmp13139 : 1);
  assign tmp13149 = s1 ? tmp13148 : tmp13150;
  assign tmp13146 = s2 ? tmp13147 : tmp13149;
  assign tmp13152 = s1 ? tmp13139 : tmp12916;
  assign tmp13154 = s0 ? 1 : tmp13136;
  assign tmp13153 = ~(s1 ? tmp13136 : tmp13154);
  assign tmp13151 = ~(s2 ? tmp13152 : tmp13153);
  assign tmp13145 = s3 ? tmp13146 : tmp13151;
  assign tmp13133 = s4 ? tmp13134 : tmp13145;
  assign tmp13160 = ~(s0 ? 1 : tmp13141);
  assign tmp13159 = s1 ? tmp13148 : tmp13160;
  assign tmp13162 = s0 ? 1 : tmp13141;
  assign tmp13163 = ~(s0 ? tmp13136 : tmp13137);
  assign tmp13161 = ~(s1 ? tmp13162 : tmp13163);
  assign tmp13158 = s2 ? tmp13159 : tmp13161;
  assign tmp13165 = s0 ? tmp13140 : tmp13141;
  assign tmp13166 = ~(s1 ? 1 : tmp13136);
  assign tmp13164 = ~(s2 ? tmp13165 : tmp13166);
  assign tmp13157 = s3 ? tmp13158 : tmp13164;
  assign tmp13170 = ~(s0 ? 1 : tmp12905);
  assign tmp13169 = s1 ? tmp13154 : tmp13170;
  assign tmp13172 = ~(s0 ? tmp13136 : 0);
  assign tmp13171 = ~(s1 ? tmp13006 : tmp13172);
  assign tmp13168 = s2 ? tmp13169 : tmp13171;
  assign tmp13174 = s1 ? tmp13136 : tmp12904;
  assign tmp13173 = s2 ? tmp13174 : 1;
  assign tmp13167 = s3 ? tmp13168 : tmp13173;
  assign tmp13156 = s4 ? tmp13157 : tmp13167;
  assign tmp13179 = s0 ? tmp13136 : 1;
  assign tmp13178 = s1 ? tmp13179 : 1;
  assign tmp13181 = s0 ? tmp12903 : tmp13136;
  assign tmp13180 = s1 ? tmp13154 : tmp13181;
  assign tmp13177 = s2 ? tmp13178 : tmp13180;
  assign tmp13176 = s3 ? tmp13177 : tmp13106;
  assign tmp13184 = s1 ? tmp12903 : 1;
  assign tmp13186 = s0 ? tmp13136 : tmp12903;
  assign tmp13185 = s1 ? tmp13154 : tmp13186;
  assign tmp13183 = s2 ? tmp13184 : tmp13185;
  assign tmp13182 = s3 ? tmp13183 : tmp12946;
  assign tmp13175 = s4 ? tmp13176 : tmp13182;
  assign tmp13155 = s5 ? tmp13156 : tmp13175;
  assign tmp13132 = s6 ? tmp13133 : tmp13155;
  assign tmp13192 = ~(l1 ? 1 : tmp13140);
  assign tmp13191 = s1 ? tmp13148 : tmp13192;
  assign tmp13190 = s2 ? tmp13147 : tmp13191;
  assign tmp13194 = s1 ? tmp13139 : 0;
  assign tmp13193 = ~(s2 ? tmp13194 : tmp13153);
  assign tmp13189 = s3 ? tmp13190 : tmp13193;
  assign tmp13188 = s4 ? tmp13134 : tmp13189;
  assign tmp13199 = s1 ? tmp13136 : tmp13144;
  assign tmp13198 = s2 ? tmp13147 : tmp13199;
  assign tmp13201 = s1 ? 1 : tmp13136;
  assign tmp13200 = s2 ? tmp13136 : tmp13201;
  assign tmp13197 = s3 ? tmp13198 : tmp13200;
  assign tmp13203 = s2 ? tmp13169 : tmp13136;
  assign tmp13205 = s1 ? tmp13136 : tmp12903;
  assign tmp13204 = s2 ? tmp13205 : 1;
  assign tmp13202 = s3 ? tmp13203 : tmp13204;
  assign tmp13196 = s4 ? tmp13197 : tmp13202;
  assign tmp13208 = s2 ? tmp13178 : tmp13205;
  assign tmp13207 = s3 ? tmp13208 : tmp13128;
  assign tmp13211 = s1 ? tmp13136 : tmp13071;
  assign tmp13210 = s2 ? 1 : tmp13211;
  assign tmp13209 = s3 ? tmp13210 : tmp12903;
  assign tmp13206 = s4 ? tmp13207 : tmp13209;
  assign tmp13195 = s5 ? tmp13196 : tmp13206;
  assign tmp13187 = s6 ? tmp13188 : tmp13195;
  assign tmp13131 = s7 ? tmp13132 : tmp13187;
  assign tmp13065 = s8 ? tmp13066 : tmp13131;
  assign tmp13220 = s0 ? tmp12903 : tmp13071;
  assign tmp13219 = s1 ? tmp13220 : tmp13071;
  assign tmp13218 = s2 ? tmp13104 : tmp13219;
  assign tmp13217 = s3 ? tmp13218 : tmp13106;
  assign tmp13216 = s4 ? tmp13217 : tmp13107;
  assign tmp13215 = s5 ? tmp13085 : tmp13216;
  assign tmp13214 = s6 ? tmp13068 : tmp13215;
  assign tmp13225 = s2 ? tmp13104 : tmp13125;
  assign tmp13226 = s2 ? tmp12938 : tmp12927;
  assign tmp13224 = s3 ? tmp13225 : tmp13226;
  assign tmp13223 = s4 ? tmp13224 : tmp13129;
  assign tmp13222 = s5 ? tmp13116 : tmp13223;
  assign tmp13221 = s6 ? tmp13111 : tmp13222;
  assign tmp13213 = s7 ? tmp13214 : tmp13221;
  assign tmp13212 = s8 ? tmp13131 : tmp13213;
  assign tmp13064 = s9 ? tmp13065 : tmp13212;
  assign tmp13233 = s3 ? tmp13225 : tmp13128;
  assign tmp13232 = s4 ? tmp13233 : tmp13129;
  assign tmp13231 = s5 ? tmp13116 : tmp13232;
  assign tmp13230 = s6 ? tmp13111 : tmp13231;
  assign tmp13229 = s7 ? tmp13067 : tmp13230;
  assign tmp13228 = s8 ? tmp13229 : tmp13067;
  assign tmp13235 = s7 ? tmp13110 : tmp13221;
  assign tmp13241 = s2 ? 1 : tmp13136;
  assign tmp13240 = s3 ? tmp13241 : tmp12903;
  assign tmp13239 = s4 ? tmp13207 : tmp13240;
  assign tmp13238 = s5 ? tmp13196 : tmp13239;
  assign tmp13237 = s6 ? tmp13188 : tmp13238;
  assign tmp13236 = s7 ? tmp13237 : tmp13230;
  assign tmp13234 = s8 ? tmp13235 : tmp13236;
  assign tmp13227 = s9 ? tmp13228 : tmp13234;
  assign tmp13063 = s10 ? tmp13064 : tmp13227;
  assign tmp13245 = s7 ? tmp13187 : tmp13230;
  assign tmp13244 = s8 ? tmp13235 : tmp13245;
  assign tmp13243 = s9 ? tmp13228 : tmp13244;
  assign tmp13242 = s10 ? tmp13064 : tmp13243;
  assign tmp13062 = s11 ? tmp13063 : tmp13242;
  assign tmp13254 = s1 ? tmp12903 : tmp13100;
  assign tmp13253 = s3 ? tmp13254 : tmp12907;
  assign tmp13256 = s2 ? tmp12908 : tmp12923;
  assign tmp13257 = ~(s2 ? tmp13081 : tmp12906);
  assign tmp13255 = s3 ? tmp13256 : tmp13257;
  assign tmp13252 = s4 ? tmp13253 : tmp13255;
  assign tmp13262 = s1 ? tmp12909 : tmp13100;
  assign tmp13261 = s2 ? tmp13262 : tmp12975;
  assign tmp13260 = s3 ? tmp13261 : tmp12976;
  assign tmp13265 = ~(s1 ? 1 : tmp12933);
  assign tmp13264 = s2 ? tmp12945 : tmp13265;
  assign tmp13266 = s2 ? tmp13254 : 1;
  assign tmp13263 = s3 ? tmp13264 : tmp13266;
  assign tmp13259 = s4 ? tmp13260 : tmp13263;
  assign tmp13269 = s2 ? tmp12938 : tmp12903;
  assign tmp13268 = s3 ? tmp13269 : tmp13106;
  assign tmp13272 = s1 ? tmp12918 : tmp12903;
  assign tmp13271 = s2 ? tmp12903 : tmp13272;
  assign tmp13270 = s3 ? tmp13271 : tmp12946;
  assign tmp13267 = s4 ? tmp13268 : tmp13270;
  assign tmp13258 = s5 ? tmp13259 : tmp13267;
  assign tmp13251 = s6 ? tmp13252 : tmp13258;
  assign tmp13276 = ~(s2 ? tmp13114 : tmp12906);
  assign tmp13275 = s3 ? tmp13256 : tmp13276;
  assign tmp13274 = s4 ? tmp13253 : tmp13275;
  assign tmp13280 = s2 ? tmp12908 : tmp12983;
  assign tmp13279 = s3 ? tmp13280 : tmp12926;
  assign tmp13282 = s2 ? tmp12945 : tmp12903;
  assign tmp13281 = s3 ? tmp13282 : tmp12986;
  assign tmp13278 = s4 ? tmp13279 : tmp13281;
  assign tmp13284 = s3 ? tmp13269 : tmp13128;
  assign tmp13285 = s3 ? tmp13071 : tmp12903;
  assign tmp13283 = s4 ? tmp13284 : tmp13285;
  assign tmp13277 = s5 ? tmp13278 : tmp13283;
  assign tmp13273 = s6 ? tmp13274 : tmp13277;
  assign tmp13250 = s7 ? tmp13251 : tmp13273;
  assign tmp13291 = l1 ? tmp12903 : 1;
  assign tmp13293 = ~(l1 ? tmp12903 : 1);
  assign tmp13292 = ~(s0 ? tmp12905 : tmp13293);
  assign tmp13290 = s1 ? tmp13291 : tmp13292;
  assign tmp13296 = s0 ? tmp13291 : 1;
  assign tmp13295 = s1 ? tmp13296 : tmp13291;
  assign tmp13294 = s2 ? tmp13291 : tmp13295;
  assign tmp13289 = s3 ? tmp13290 : tmp13294;
  assign tmp13300 = s0 ? tmp13291 : 0;
  assign tmp13299 = s1 ? tmp13300 : tmp13291;
  assign tmp13301 = s1 ? tmp13300 : tmp12913;
  assign tmp13298 = s2 ? tmp13299 : tmp13301;
  assign tmp13302 = ~(s2 ? tmp12915 : tmp13293);
  assign tmp13297 = s3 ? tmp13298 : tmp13302;
  assign tmp13288 = s4 ? tmp13289 : tmp13297;
  assign tmp13308 = ~(s0 ? 1 : tmp13293);
  assign tmp13307 = s1 ? tmp13300 : tmp13308;
  assign tmp13310 = s0 ? 1 : tmp13293;
  assign tmp13311 = ~(s0 ? tmp13291 : 1);
  assign tmp13309 = ~(s1 ? tmp13310 : tmp13311);
  assign tmp13306 = s2 ? tmp13307 : tmp13309;
  assign tmp13313 = s0 ? 1 : tmp13291;
  assign tmp13314 = s1 ? 1 : tmp13291;
  assign tmp13312 = s2 ? tmp13313 : tmp13314;
  assign tmp13305 = s3 ? tmp13306 : tmp13312;
  assign tmp13317 = s1 ? tmp13313 : tmp13170;
  assign tmp13319 = ~(s0 ? tmp13291 : 0);
  assign tmp13318 = ~(s1 ? tmp13006 : tmp13319);
  assign tmp13316 = s2 ? tmp13317 : tmp13318;
  assign tmp13321 = s1 ? tmp13291 : tmp12904;
  assign tmp13320 = s2 ? tmp13321 : 1;
  assign tmp13315 = s3 ? tmp13316 : tmp13320;
  assign tmp13304 = s4 ? tmp13305 : tmp13315;
  assign tmp13325 = s1 ? tmp13296 : 1;
  assign tmp13327 = s0 ? tmp12903 : tmp13291;
  assign tmp13326 = s1 ? tmp13291 : tmp13327;
  assign tmp13324 = s2 ? tmp13325 : tmp13326;
  assign tmp13323 = s3 ? tmp13324 : tmp13106;
  assign tmp13331 = s0 ? tmp13291 : tmp12903;
  assign tmp13330 = s1 ? tmp13313 : tmp13331;
  assign tmp13329 = s2 ? tmp13184 : tmp13330;
  assign tmp13328 = s3 ? tmp13329 : tmp12946;
  assign tmp13322 = s4 ? tmp13323 : tmp13328;
  assign tmp13303 = s5 ? tmp13304 : tmp13322;
  assign tmp13287 = s6 ? tmp13288 : tmp13303;
  assign tmp13336 = s1 ? tmp13300 : tmp12931;
  assign tmp13335 = s2 ? tmp13299 : tmp13336;
  assign tmp13337 = ~(s2 ? tmp12955 : tmp13293);
  assign tmp13334 = s3 ? tmp13335 : tmp13337;
  assign tmp13333 = s4 ? tmp13289 : tmp13334;
  assign tmp13342 = s1 ? tmp13291 : tmp13296;
  assign tmp13341 = s2 ? tmp13299 : tmp13342;
  assign tmp13343 = s2 ? tmp13291 : tmp13314;
  assign tmp13340 = s3 ? tmp13341 : tmp13343;
  assign tmp13345 = s2 ? tmp13317 : tmp13291;
  assign tmp13347 = s1 ? tmp13291 : tmp12903;
  assign tmp13346 = s2 ? tmp13347 : 1;
  assign tmp13344 = s3 ? tmp13345 : tmp13346;
  assign tmp13339 = s4 ? tmp13340 : tmp13344;
  assign tmp13350 = s2 ? tmp13325 : tmp13347;
  assign tmp13349 = s3 ? tmp13350 : tmp13128;
  assign tmp13353 = s1 ? tmp13291 : tmp13071;
  assign tmp13352 = s2 ? 1 : tmp13353;
  assign tmp13351 = s3 ? tmp13352 : tmp12903;
  assign tmp13348 = s4 ? tmp13349 : tmp13351;
  assign tmp13338 = s5 ? tmp13339 : tmp13348;
  assign tmp13332 = s6 ? tmp13333 : tmp13338;
  assign tmp13286 = s7 ? tmp13287 : tmp13332;
  assign tmp13249 = s8 ? tmp13250 : tmp13286;
  assign tmp13360 = s2 ? tmp13262 : tmp12924;
  assign tmp13359 = s3 ? tmp13360 : tmp12926;
  assign tmp13358 = s4 ? tmp13359 : tmp13263;
  assign tmp13357 = s5 ? tmp13358 : tmp13267;
  assign tmp13356 = s6 ? tmp13252 : tmp13357;
  assign tmp13365 = s2 ? tmp12908 : tmp12903;
  assign tmp13364 = s3 ? tmp13365 : tmp12926;
  assign tmp13363 = s4 ? tmp13364 : tmp13281;
  assign tmp13367 = s3 ? tmp13269 : tmp13226;
  assign tmp13366 = s4 ? tmp13367 : tmp12903;
  assign tmp13362 = s5 ? tmp13363 : tmp13366;
  assign tmp13361 = s6 ? tmp13274 : tmp13362;
  assign tmp13355 = s7 ? tmp13356 : tmp13361;
  assign tmp13354 = s8 ? tmp13286 : tmp13355;
  assign tmp13248 = s9 ? tmp13249 : tmp13354;
  assign tmp13372 = s5 ? tmp13363 : tmp13283;
  assign tmp13371 = s6 ? tmp13274 : tmp13372;
  assign tmp13370 = s7 ? tmp13356 : tmp13371;
  assign tmp13369 = s8 ? tmp13370 : tmp13356;
  assign tmp13377 = s3 ? tmp12968 : tmp12903;
  assign tmp13376 = s4 ? tmp13284 : tmp13377;
  assign tmp13375 = s5 ? tmp13278 : tmp13376;
  assign tmp13374 = s6 ? tmp13274 : tmp13375;
  assign tmp13383 = s2 ? 1 : tmp13291;
  assign tmp13382 = s3 ? tmp13383 : tmp12903;
  assign tmp13381 = s4 ? tmp13349 : tmp13382;
  assign tmp13380 = s5 ? tmp13339 : tmp13381;
  assign tmp13379 = s6 ? tmp13333 : tmp13380;
  assign tmp13385 = s5 ? tmp13363 : tmp13376;
  assign tmp13384 = s6 ? tmp13274 : tmp13385;
  assign tmp13378 = s7 ? tmp13379 : tmp13384;
  assign tmp13373 = s8 ? tmp13374 : tmp13378;
  assign tmp13368 = s9 ? tmp13369 : tmp13373;
  assign tmp13247 = s10 ? tmp13248 : tmp13368;
  assign tmp13389 = s7 ? tmp13332 : tmp13371;
  assign tmp13388 = s8 ? tmp13273 : tmp13389;
  assign tmp13387 = s9 ? tmp13369 : tmp13388;
  assign tmp13386 = s10 ? tmp13248 : tmp13387;
  assign tmp13246 = s11 ? tmp13247 : tmp13386;
  assign tmp13061 = ~(s12 ? tmp13062 : tmp13246);
  assign tmp12892 = s13 ? tmp12893 : tmp13061;
  assign tmp12891 = s14 ? 1 : tmp12892;
  assign tmp13404 = ~(l4 ? 1 : 0);
  assign tmp13403 = l2 ? 1 : tmp13404;
  assign tmp13402 = l1 ? tmp12903 : tmp13403;
  assign tmp13406 = ~(l1 ? tmp12903 : tmp13403);
  assign tmp13405 = ~(s0 ? tmp12905 : tmp13406);
  assign tmp13401 = s1 ? tmp13402 : tmp13405;
  assign tmp13408 = s1 ? tmp12909 : tmp13402;
  assign tmp13407 = s2 ? tmp13402 : tmp13408;
  assign tmp13400 = s3 ? tmp13401 : tmp13407;
  assign tmp13412 = s0 ? tmp13402 : 0;
  assign tmp13411 = s1 ? tmp13412 : tmp13402;
  assign tmp13413 = s1 ? tmp13412 : tmp12913;
  assign tmp13410 = s2 ? tmp13411 : tmp13413;
  assign tmp13416 = s0 ? tmp13291 : tmp13402;
  assign tmp13415 = ~(s1 ? tmp13402 : tmp13416);
  assign tmp13414 = ~(s2 ? tmp12915 : tmp13415);
  assign tmp13409 = s3 ? tmp13410 : tmp13414;
  assign tmp13399 = s4 ? tmp13400 : tmp13409;
  assign tmp13421 = s1 ? tmp13412 : tmp13100;
  assign tmp13423 = s0 ? 1 : tmp13406;
  assign tmp13424 = ~(s0 ? tmp13402 : 0);
  assign tmp13422 = ~(s1 ? tmp13423 : tmp13424);
  assign tmp13420 = s2 ? tmp13421 : tmp13422;
  assign tmp13426 = ~(s1 ? tmp13296 : tmp13402);
  assign tmp13425 = ~(s2 ? tmp13423 : tmp13426);
  assign tmp13419 = s3 ? tmp13420 : tmp13425;
  assign tmp13430 = s0 ? 1 : tmp13402;
  assign tmp13429 = s1 ? tmp13430 : tmp12931;
  assign tmp13431 = ~(s1 ? tmp12905 : tmp13424);
  assign tmp13428 = s2 ? tmp13429 : tmp13431;
  assign tmp13432 = s2 ? tmp13401 : 1;
  assign tmp13427 = s3 ? tmp13428 : tmp13432;
  assign tmp13418 = s4 ? tmp13419 : tmp13427;
  assign tmp13437 = s0 ? tmp13402 : 1;
  assign tmp13436 = s1 ? tmp13437 : 1;
  assign tmp13435 = s2 ? tmp13436 : tmp13272;
  assign tmp13439 = s1 ? 1 : tmp13430;
  assign tmp13438 = s2 ? tmp12938 : tmp13439;
  assign tmp13434 = s3 ? tmp13435 : tmp13438;
  assign tmp13442 = s1 ? tmp13437 : tmp13313;
  assign tmp13443 = s1 ? tmp13430 : tmp12903;
  assign tmp13441 = s2 ? tmp13442 : tmp13443;
  assign tmp13445 = s1 ? tmp13430 : 1;
  assign tmp13444 = s2 ? tmp13439 : tmp13445;
  assign tmp13440 = s3 ? tmp13441 : tmp13444;
  assign tmp13433 = s4 ? tmp13434 : tmp13440;
  assign tmp13417 = s5 ? tmp13418 : tmp13433;
  assign tmp13398 = s6 ? tmp13399 : tmp13417;
  assign tmp13450 = s1 ? tmp13412 : tmp12931;
  assign tmp13449 = s2 ? tmp13411 : tmp13450;
  assign tmp13451 = ~(s2 ? tmp12955 : tmp13415);
  assign tmp13448 = s3 ? tmp13449 : tmp13451;
  assign tmp13447 = s4 ? tmp13400 : tmp13448;
  assign tmp13456 = s1 ? tmp13412 : tmp12903;
  assign tmp13457 = s1 ? tmp13402 : tmp13412;
  assign tmp13455 = s2 ? tmp13456 : tmp13457;
  assign tmp13459 = s1 ? tmp13296 : tmp13402;
  assign tmp13458 = s2 ? tmp13402 : tmp13459;
  assign tmp13454 = s3 ? tmp13455 : tmp13458;
  assign tmp13462 = ~(s1 ? tmp12905 : tmp13406);
  assign tmp13461 = s2 ? tmp13429 : tmp13462;
  assign tmp13460 = s3 ? tmp13461 : tmp13432;
  assign tmp13453 = s4 ? tmp13454 : tmp13460;
  assign tmp13465 = s2 ? tmp13436 : tmp12903;
  assign tmp13467 = s1 ? 1 : tmp13402;
  assign tmp13466 = s2 ? tmp13104 : tmp13467;
  assign tmp13464 = s3 ? tmp13465 : tmp13466;
  assign tmp13470 = s1 ? tmp13437 : tmp13291;
  assign tmp13469 = s2 ? tmp13470 : tmp13402;
  assign tmp13471 = s2 ? tmp13467 : tmp13402;
  assign tmp13468 = s3 ? tmp13469 : tmp13471;
  assign tmp13463 = s4 ? tmp13464 : tmp13468;
  assign tmp13452 = s5 ? tmp13453 : tmp13463;
  assign tmp13446 = s6 ? tmp13447 : tmp13452;
  assign tmp13397 = s7 ? tmp13398 : tmp13446;
  assign tmp13475 = s3 ? tmp13401 : tmp13458;
  assign tmp13474 = s4 ? tmp13475 : tmp13409;
  assign tmp13480 = s1 ? tmp13412 : tmp13308;
  assign tmp13482 = ~(s0 ? tmp13402 : 1);
  assign tmp13481 = ~(s1 ? tmp13423 : tmp13482);
  assign tmp13479 = s2 ? tmp13480 : tmp13481;
  assign tmp13483 = s2 ? tmp13430 : tmp13467;
  assign tmp13478 = s3 ? tmp13479 : tmp13483;
  assign tmp13486 = s1 ? tmp13430 : tmp13170;
  assign tmp13487 = ~(s1 ? tmp13006 : tmp13424);
  assign tmp13485 = s2 ? tmp13486 : tmp13487;
  assign tmp13484 = s3 ? tmp13485 : tmp13432;
  assign tmp13477 = s4 ? tmp13478 : tmp13484;
  assign tmp13491 = s1 ? tmp13313 : tmp13327;
  assign tmp13490 = s2 ? tmp13436 : tmp13491;
  assign tmp13489 = s3 ? tmp13490 : tmp13438;
  assign tmp13494 = s1 ? tmp13430 : tmp13331;
  assign tmp13493 = s2 ? tmp13436 : tmp13494;
  assign tmp13492 = s3 ? tmp13493 : tmp13444;
  assign tmp13488 = s4 ? tmp13489 : tmp13492;
  assign tmp13476 = s5 ? tmp13477 : tmp13488;
  assign tmp13473 = s6 ? tmp13474 : tmp13476;
  assign tmp13496 = s4 ? tmp13475 : tmp13448;
  assign tmp13501 = s1 ? tmp13412 : tmp13291;
  assign tmp13502 = s1 ? tmp13402 : tmp13437;
  assign tmp13500 = s2 ? tmp13501 : tmp13502;
  assign tmp13503 = s2 ? tmp13402 : tmp13467;
  assign tmp13499 = s3 ? tmp13500 : tmp13503;
  assign tmp13505 = s2 ? tmp13486 : tmp13402;
  assign tmp13506 = s2 ? tmp13402 : 1;
  assign tmp13504 = s3 ? tmp13505 : tmp13506;
  assign tmp13498 = s4 ? tmp13499 : tmp13504;
  assign tmp13509 = s2 ? tmp13436 : tmp13347;
  assign tmp13508 = s3 ? tmp13509 : tmp13466;
  assign tmp13511 = s2 ? tmp13436 : tmp13402;
  assign tmp13510 = s3 ? tmp13511 : tmp13471;
  assign tmp13507 = s4 ? tmp13508 : tmp13510;
  assign tmp13497 = s5 ? tmp13498 : tmp13507;
  assign tmp13495 = s6 ? tmp13496 : tmp13497;
  assign tmp13472 = s7 ? tmp13473 : tmp13495;
  assign tmp13396 = s8 ? tmp13397 : tmp13472;
  assign tmp13517 = s2 ? tmp13291 : tmp13299;
  assign tmp13516 = s3 ? tmp13290 : tmp13517;
  assign tmp13515 = s4 ? tmp13516 : tmp13297;
  assign tmp13522 = s1 ? tmp13300 : tmp13100;
  assign tmp13524 = ~(s0 ? tmp13291 : tmp12903);
  assign tmp13523 = ~(s1 ? tmp13310 : tmp13524);
  assign tmp13521 = s2 ? tmp13522 : tmp13523;
  assign tmp13525 = s2 ? tmp13327 : tmp13295;
  assign tmp13520 = s3 ? tmp13521 : tmp13525;
  assign tmp13528 = s1 ? tmp13313 : tmp12931;
  assign tmp13529 = ~(s1 ? tmp12905 : tmp13319);
  assign tmp13527 = s2 ? tmp13528 : tmp13529;
  assign tmp13530 = s2 ? tmp13290 : 1;
  assign tmp13526 = s3 ? tmp13527 : tmp13530;
  assign tmp13519 = s4 ? tmp13520 : tmp13526;
  assign tmp13533 = s2 ? tmp13325 : tmp13272;
  assign tmp13535 = s1 ? 1 : tmp13313;
  assign tmp13534 = s2 ? tmp12938 : tmp13535;
  assign tmp13532 = s3 ? tmp13533 : tmp13534;
  assign tmp13538 = s1 ? tmp13296 : tmp13313;
  assign tmp13539 = s1 ? tmp13313 : tmp12903;
  assign tmp13537 = s2 ? tmp13538 : tmp13539;
  assign tmp13541 = s1 ? tmp13313 : 1;
  assign tmp13540 = s2 ? tmp13535 : tmp13541;
  assign tmp13536 = s3 ? tmp13537 : tmp13540;
  assign tmp13531 = s4 ? tmp13532 : tmp13536;
  assign tmp13518 = s5 ? tmp13519 : tmp13531;
  assign tmp13514 = s6 ? tmp13515 : tmp13518;
  assign tmp13543 = s4 ? tmp13516 : tmp13334;
  assign tmp13548 = s1 ? tmp13300 : tmp12903;
  assign tmp13549 = s1 ? tmp13291 : tmp13331;
  assign tmp13547 = s2 ? tmp13548 : tmp13549;
  assign tmp13546 = s3 ? tmp13547 : tmp13294;
  assign tmp13551 = s2 ? tmp13528 : tmp13291;
  assign tmp13552 = s2 ? tmp13291 : 1;
  assign tmp13550 = s3 ? tmp13551 : tmp13552;
  assign tmp13545 = s4 ? tmp13546 : tmp13550;
  assign tmp13555 = s2 ? tmp13325 : tmp12903;
  assign tmp13556 = s2 ? tmp12938 : tmp13314;
  assign tmp13554 = s3 ? tmp13555 : tmp13556;
  assign tmp13558 = s2 ? tmp13295 : tmp13291;
  assign tmp13559 = s2 ? tmp13314 : tmp13291;
  assign tmp13557 = s3 ? tmp13558 : tmp13559;
  assign tmp13553 = s4 ? tmp13554 : tmp13557;
  assign tmp13544 = s5 ? tmp13545 : tmp13553;
  assign tmp13542 = s6 ? tmp13543 : tmp13544;
  assign tmp13513 = s7 ? tmp13514 : tmp13542;
  assign tmp13512 = s8 ? tmp13472 : tmp13513;
  assign tmp13395 = s9 ? tmp13396 : tmp13512;
  assign tmp13569 = ~(s0 ? tmp13402 : tmp12903);
  assign tmp13568 = ~(s1 ? tmp13423 : tmp13569);
  assign tmp13567 = s2 ? tmp13421 : tmp13568;
  assign tmp13571 = s0 ? tmp12903 : tmp13402;
  assign tmp13570 = s2 ? tmp13571 : tmp13459;
  assign tmp13566 = s3 ? tmp13567 : tmp13570;
  assign tmp13565 = s4 ? tmp13566 : tmp13427;
  assign tmp13564 = s5 ? tmp13565 : tmp13433;
  assign tmp13563 = s6 ? tmp13399 : tmp13564;
  assign tmp13578 = s0 ? tmp13402 : tmp12903;
  assign tmp13577 = s1 ? tmp13402 : tmp13578;
  assign tmp13576 = s2 ? tmp13456 : tmp13577;
  assign tmp13575 = s3 ? tmp13576 : tmp13458;
  assign tmp13580 = s2 ? tmp13429 : tmp13402;
  assign tmp13579 = s3 ? tmp13580 : tmp13506;
  assign tmp13574 = s4 ? tmp13575 : tmp13579;
  assign tmp13573 = s5 ? tmp13574 : tmp13463;
  assign tmp13572 = s6 ? tmp13447 : tmp13573;
  assign tmp13562 = s7 ? tmp13563 : tmp13572;
  assign tmp13561 = s8 ? tmp13562 : tmp13563;
  assign tmp13586 = s3 ? tmp13461 : tmp13506;
  assign tmp13585 = s4 ? tmp13454 : tmp13586;
  assign tmp13588 = s3 ? tmp13469 : tmp13467;
  assign tmp13587 = s4 ? tmp13464 : tmp13588;
  assign tmp13584 = s5 ? tmp13585 : tmp13587;
  assign tmp13583 = s6 ? tmp13447 : tmp13584;
  assign tmp13592 = s3 ? tmp13558 : tmp13314;
  assign tmp13591 = s4 ? tmp13554 : tmp13592;
  assign tmp13590 = s5 ? tmp13545 : tmp13591;
  assign tmp13589 = s6 ? tmp13543 : tmp13590;
  assign tmp13582 = s7 ? tmp13583 : tmp13589;
  assign tmp13597 = s3 ? tmp13511 : tmp13467;
  assign tmp13596 = s4 ? tmp13508 : tmp13597;
  assign tmp13595 = s5 ? tmp13498 : tmp13596;
  assign tmp13594 = s6 ? tmp13496 : tmp13595;
  assign tmp13599 = s5 ? tmp13574 : tmp13587;
  assign tmp13598 = s6 ? tmp13447 : tmp13599;
  assign tmp13593 = s7 ? tmp13594 : tmp13598;
  assign tmp13581 = s8 ? tmp13582 : tmp13593;
  assign tmp13560 = s9 ? tmp13561 : tmp13581;
  assign tmp13394 = s10 ? tmp13395 : tmp13560;
  assign tmp13603 = s7 ? tmp13446 : tmp13542;
  assign tmp13604 = s7 ? tmp13495 : tmp13572;
  assign tmp13602 = s8 ? tmp13603 : tmp13604;
  assign tmp13601 = s9 ? tmp13561 : tmp13602;
  assign tmp13600 = s10 ? tmp13395 : tmp13601;
  assign tmp13393 = s11 ? tmp13394 : tmp13600;
  assign tmp13392 = s12 ? tmp13393 : 1;
  assign tmp13391 = s13 ? tmp13392 : 1;
  assign tmp13390 = ~(s14 ? 1 : tmp13391);
  assign tmp12890 = s15 ? tmp12891 : tmp13390;
  assign tmp13616 = s4 ? tmp12981 : tmp12960;
  assign tmp13615 = s5 ? tmp13616 : tmp12963;
  assign tmp13614 = s6 ? tmp12950 : tmp13615;
  assign tmp13613 = s7 ? tmp12970 : tmp13614;
  assign tmp13624 = l4 ? 1 : 0;
  assign tmp13623 = l2 ? tmp13624 : 1;
  assign tmp13622 = l1 ? 1 : tmp13623;
  assign tmp13626 = l1 ? 1 : tmp13624;
  assign tmp13625 = s0 ? tmp13626 : tmp13622;
  assign tmp13621 = s1 ? tmp13622 : tmp13625;
  assign tmp13629 = s0 ? tmp13622 : 1;
  assign tmp13628 = s1 ? tmp13629 : tmp13622;
  assign tmp13627 = s2 ? tmp13622 : tmp13628;
  assign tmp13620 = s3 ? tmp13621 : tmp13627;
  assign tmp13633 = s0 ? tmp13626 : 1;
  assign tmp13632 = s1 ? tmp13629 : tmp13633;
  assign tmp13631 = s2 ? tmp13628 : tmp13632;
  assign tmp13635 = s1 ? tmp13626 : tmp12916;
  assign tmp13637 = s0 ? tmp13624 : tmp13622;
  assign tmp13636 = s1 ? tmp13622 : tmp13637;
  assign tmp13634 = s2 ? tmp13635 : tmp13636;
  assign tmp13630 = s3 ? tmp13631 : tmp13634;
  assign tmp13619 = s4 ? tmp13620 : tmp13630;
  assign tmp13642 = s1 ? tmp13629 : 1;
  assign tmp13644 = s0 ? 1 : tmp13622;
  assign tmp13643 = s1 ? tmp13644 : tmp13629;
  assign tmp13641 = s2 ? tmp13642 : tmp13643;
  assign tmp13647 = s0 ? tmp13624 : 0;
  assign tmp13646 = s1 ? tmp13647 : tmp13622;
  assign tmp13645 = s2 ? tmp13644 : tmp13646;
  assign tmp13640 = s3 ? tmp13641 : tmp13645;
  assign tmp13652 = ~(l1 ? 1 : tmp13623);
  assign tmp13651 = s0 ? 1 : tmp13652;
  assign tmp13653 = ~(s0 ? 1 : tmp13626);
  assign tmp13650 = s1 ? tmp13651 : tmp13653;
  assign tmp13655 = s0 ? 1 : tmp13626;
  assign tmp13654 = ~(s1 ? tmp13655 : tmp13629);
  assign tmp13649 = s2 ? tmp13650 : tmp13654;
  assign tmp13658 = s0 ? tmp13626 : tmp12906;
  assign tmp13657 = s1 ? tmp13622 : tmp13658;
  assign tmp13656 = ~(s2 ? tmp13657 : 0);
  assign tmp13648 = ~(s3 ? tmp13649 : tmp13656);
  assign tmp13639 = s4 ? tmp13640 : tmp13648;
  assign tmp13663 = s0 ? tmp13622 : 0;
  assign tmp13664 = ~(s0 ? 1 : tmp13404);
  assign tmp13662 = s1 ? tmp13663 : tmp13664;
  assign tmp13666 = s0 ? tmp13624 : 1;
  assign tmp13665 = s1 ? tmp13666 : 1;
  assign tmp13661 = s2 ? tmp13662 : tmp13665;
  assign tmp13667 = s2 ? tmp12940 : tmp12942;
  assign tmp13660 = s3 ? tmp13661 : tmp13667;
  assign tmp13671 = s0 ? 1 : tmp13404;
  assign tmp13670 = s1 ? tmp12939 : tmp13671;
  assign tmp13672 = s1 ? tmp13651 : 0;
  assign tmp13669 = s2 ? tmp13670 : tmp13672;
  assign tmp13675 = ~(s0 ? 1 : tmp12903);
  assign tmp13674 = s1 ? tmp13647 : tmp13675;
  assign tmp13676 = ~(s1 ? tmp12918 : 1);
  assign tmp13673 = ~(s2 ? tmp13674 : tmp13676);
  assign tmp13668 = ~(s3 ? tmp13669 : tmp13673);
  assign tmp13659 = s4 ? tmp13660 : tmp13668;
  assign tmp13638 = s5 ? tmp13639 : tmp13659;
  assign tmp13618 = s6 ? tmp13619 : tmp13638;
  assign tmp13681 = s1 ? tmp13629 : tmp13626;
  assign tmp13680 = s2 ? tmp13628 : tmp13681;
  assign tmp13683 = s1 ? tmp13626 : 0;
  assign tmp13682 = s2 ? tmp13683 : tmp13636;
  assign tmp13679 = s3 ? tmp13680 : tmp13682;
  assign tmp13678 = s4 ? tmp13620 : tmp13679;
  assign tmp13688 = s1 ? tmp13622 : tmp13629;
  assign tmp13687 = s2 ? tmp13642 : tmp13688;
  assign tmp13689 = s2 ? tmp13622 : tmp13646;
  assign tmp13686 = s3 ? tmp13687 : tmp13689;
  assign tmp13692 = ~(s1 ? tmp13626 : tmp13622);
  assign tmp13691 = s2 ? tmp13650 : tmp13692;
  assign tmp13690 = ~(s3 ? tmp13691 : tmp13656);
  assign tmp13685 = s4 ? tmp13686 : tmp13690;
  assign tmp13696 = s1 ? tmp13663 : tmp13624;
  assign tmp13695 = s2 ? tmp13696 : 1;
  assign tmp13697 = ~(s2 ? 1 : tmp12927);
  assign tmp13694 = s3 ? tmp13695 : tmp13697;
  assign tmp13700 = s1 ? 1 : tmp13404;
  assign tmp13699 = s2 ? tmp13700 : tmp13652;
  assign tmp13698 = ~(s3 ? tmp13699 : tmp12927);
  assign tmp13693 = s4 ? tmp13694 : tmp13698;
  assign tmp13684 = s5 ? tmp13685 : tmp13693;
  assign tmp13677 = s6 ? tmp13678 : tmp13684;
  assign tmp13617 = ~(s7 ? tmp13618 : tmp13677);
  assign tmp13612 = s8 ? tmp13613 : tmp13617;
  assign tmp13702 = s7 ? tmp13618 : tmp13677;
  assign tmp13708 = s1 ? tmp13633 : tmp13626;
  assign tmp13707 = s2 ? tmp13708 : tmp13633;
  assign tmp13711 = s0 ? tmp13624 : tmp13626;
  assign tmp13710 = s1 ? tmp13626 : tmp13711;
  assign tmp13709 = s2 ? tmp13635 : tmp13710;
  assign tmp13706 = s3 ? tmp13707 : tmp13709;
  assign tmp13705 = s4 ? tmp13626 : tmp13706;
  assign tmp13716 = s1 ? tmp13633 : 1;
  assign tmp13717 = s1 ? tmp13655 : tmp13626;
  assign tmp13715 = s2 ? tmp13716 : tmp13717;
  assign tmp13719 = s1 ? tmp13647 : tmp13626;
  assign tmp13718 = s2 ? tmp13626 : tmp13719;
  assign tmp13714 = s3 ? tmp13715 : tmp13718;
  assign tmp13724 = ~(l1 ? 1 : tmp13624);
  assign tmp13723 = s0 ? 1 : tmp13724;
  assign tmp13722 = s1 ? tmp13723 : tmp13653;
  assign tmp13725 = ~(s1 ? tmp13655 : tmp13633);
  assign tmp13721 = s2 ? tmp13722 : tmp13725;
  assign tmp13728 = s0 ? tmp13626 : tmp12905;
  assign tmp13727 = s1 ? tmp13626 : tmp13728;
  assign tmp13726 = ~(s2 ? tmp13727 : 0);
  assign tmp13720 = ~(s3 ? tmp13721 : tmp13726);
  assign tmp13713 = s4 ? tmp13714 : tmp13720;
  assign tmp13733 = s0 ? tmp13626 : 0;
  assign tmp13732 = s1 ? tmp13733 : tmp13664;
  assign tmp13731 = s2 ? tmp13732 : tmp13665;
  assign tmp13730 = s3 ? tmp13731 : tmp13020;
  assign tmp13736 = s1 ? tmp13018 : tmp13664;
  assign tmp13737 = ~(s1 ? tmp13723 : 0);
  assign tmp13735 = s2 ? tmp13736 : tmp13737;
  assign tmp13739 = s1 ? tmp13647 : tmp12999;
  assign tmp13740 = ~(s1 ? tmp13012 : 1);
  assign tmp13738 = s2 ? tmp13739 : tmp13740;
  assign tmp13734 = s3 ? tmp13735 : tmp13738;
  assign tmp13729 = s4 ? tmp13730 : tmp13734;
  assign tmp13712 = s5 ? tmp13713 : tmp13729;
  assign tmp13704 = s6 ? tmp13705 : tmp13712;
  assign tmp13744 = s2 ? tmp13683 : tmp13710;
  assign tmp13743 = s3 ? tmp13708 : tmp13744;
  assign tmp13742 = s4 ? tmp13626 : tmp13743;
  assign tmp13748 = s2 ? tmp13716 : tmp13626;
  assign tmp13747 = s3 ? tmp13748 : tmp13718;
  assign tmp13750 = s2 ? tmp13722 : tmp13724;
  assign tmp13749 = ~(s3 ? tmp13750 : tmp13726);
  assign tmp13746 = s4 ? tmp13747 : tmp13749;
  assign tmp13754 = s1 ? tmp13733 : tmp13624;
  assign tmp13753 = s2 ? tmp13754 : 1;
  assign tmp13752 = s3 ? tmp13753 : tmp13039;
  assign tmp13756 = s2 ? tmp13700 : tmp13724;
  assign tmp13755 = ~(s3 ? tmp13756 : tmp13040);
  assign tmp13751 = s4 ? tmp13752 : tmp13755;
  assign tmp13745 = s5 ? tmp13746 : tmp13751;
  assign tmp13741 = s6 ? tmp13742 : tmp13745;
  assign tmp13703 = s7 ? tmp13704 : tmp13741;
  assign tmp13701 = ~(s8 ? tmp13702 : tmp13703);
  assign tmp13611 = s9 ? tmp13612 : tmp13701;
  assign tmp13758 = s8 ? tmp13702 : tmp13618;
  assign tmp13763 = s4 ? tmp12981 : tmp13054;
  assign tmp13762 = s5 ? tmp13763 : tmp12963;
  assign tmp13761 = s6 ? tmp12950 : tmp13762;
  assign tmp13769 = s1 ? tmp13626 : tmp12905;
  assign tmp13768 = ~(s2 ? tmp13769 : 0);
  assign tmp13767 = ~(s3 ? tmp13750 : tmp13768);
  assign tmp13766 = s4 ? tmp13747 : tmp13767;
  assign tmp13765 = s5 ? tmp13766 : tmp13751;
  assign tmp13764 = ~(s6 ? tmp13742 : tmp13765);
  assign tmp13760 = s7 ? tmp13761 : tmp13764;
  assign tmp13775 = s1 ? tmp13622 : tmp12906;
  assign tmp13774 = ~(s2 ? tmp13775 : 0);
  assign tmp13773 = ~(s3 ? tmp13691 : tmp13774);
  assign tmp13772 = s4 ? tmp13686 : tmp13773;
  assign tmp13771 = s5 ? tmp13772 : tmp13693;
  assign tmp13770 = ~(s6 ? tmp13678 : tmp13771);
  assign tmp13759 = ~(s8 ? tmp13760 : tmp13770);
  assign tmp13757 = ~(s9 ? tmp13758 : tmp13759);
  assign tmp13610 = s10 ? tmp13611 : tmp13757;
  assign tmp13780 = ~(s6 ? tmp13742 : tmp13745);
  assign tmp13779 = s7 ? tmp13614 : tmp13780;
  assign tmp13781 = ~(s6 ? tmp13678 : tmp13684);
  assign tmp13778 = ~(s8 ? tmp13779 : tmp13781);
  assign tmp13777 = ~(s9 ? tmp13758 : tmp13778);
  assign tmp13776 = s10 ? tmp13611 : tmp13777;
  assign tmp13609 = ~(s11 ? tmp13610 : tmp13776);
  assign tmp13608 = s12 ? 1 : tmp13609;
  assign tmp13791 = l1 ? tmp12903 : tmp12906;
  assign tmp13793 = ~(l1 ? tmp12903 : tmp12906);
  assign tmp13792 = ~(s0 ? 1 : tmp13793);
  assign tmp13790 = s1 ? tmp13791 : tmp13792;
  assign tmp13796 = s0 ? tmp13791 : 0;
  assign tmp13795 = s1 ? tmp13796 : tmp13791;
  assign tmp13794 = s2 ? tmp13791 : tmp13795;
  assign tmp13789 = s3 ? tmp13790 : tmp13794;
  assign tmp13799 = s1 ? tmp13796 : 0;
  assign tmp13798 = s2 ? tmp13795 : tmp13799;
  assign tmp13802 = s0 ? 1 : tmp13791;
  assign tmp13801 = ~(s1 ? tmp13791 : tmp13802);
  assign tmp13800 = ~(s2 ? tmp13081 : tmp13801);
  assign tmp13797 = s3 ? tmp13798 : tmp13800;
  assign tmp13788 = s4 ? tmp13789 : tmp13797;
  assign tmp13807 = s1 ? tmp13796 : tmp13792;
  assign tmp13809 = s0 ? 1 : tmp13793;
  assign tmp13810 = ~(s0 ? tmp13791 : 0);
  assign tmp13808 = ~(s1 ? tmp13809 : tmp13810);
  assign tmp13806 = s2 ? tmp13807 : tmp13808;
  assign tmp13812 = ~(s1 ? 1 : tmp13791);
  assign tmp13811 = ~(s2 ? tmp13809 : tmp13812);
  assign tmp13805 = s3 ? tmp13806 : tmp13811;
  assign tmp13815 = s1 ? tmp13802 : 0;
  assign tmp13816 = ~(s1 ? 1 : tmp13810);
  assign tmp13814 = s2 ? tmp13815 : tmp13816;
  assign tmp13818 = s1 ? tmp13791 : tmp13100;
  assign tmp13817 = s2 ? tmp13818 : 1;
  assign tmp13813 = s3 ? tmp13814 : tmp13817;
  assign tmp13804 = s4 ? tmp13805 : tmp13813;
  assign tmp13824 = l1 ? 1 : tmp12906;
  assign tmp13823 = s0 ? tmp13791 : tmp13824;
  assign tmp13822 = s1 ? tmp13823 : 1;
  assign tmp13825 = s1 ? tmp13802 : tmp13791;
  assign tmp13821 = s2 ? tmp13822 : tmp13825;
  assign tmp13820 = s3 ? tmp13821 : tmp13106;
  assign tmp13829 = s0 ? tmp13824 : tmp13791;
  assign tmp13828 = s1 ? tmp13829 : tmp13791;
  assign tmp13827 = s2 ? tmp12903 : tmp13828;
  assign tmp13826 = s3 ? tmp13827 : tmp12946;
  assign tmp13819 = s4 ? tmp13820 : tmp13826;
  assign tmp13803 = s5 ? tmp13804 : tmp13819;
  assign tmp13787 = s6 ? tmp13788 : tmp13803;
  assign tmp13833 = ~(s2 ? tmp13114 : tmp13801);
  assign tmp13832 = s3 ? tmp13798 : tmp13833;
  assign tmp13831 = s4 ? tmp13789 : tmp13832;
  assign tmp13838 = s1 ? tmp13791 : tmp13796;
  assign tmp13837 = s2 ? tmp13795 : tmp13838;
  assign tmp13840 = s1 ? 1 : tmp13791;
  assign tmp13839 = s2 ? tmp13791 : tmp13840;
  assign tmp13836 = s3 ? tmp13837 : tmp13839;
  assign tmp13842 = s2 ? tmp13815 : tmp13791;
  assign tmp13844 = s1 ? tmp13791 : tmp12903;
  assign tmp13843 = s2 ? tmp13844 : 1;
  assign tmp13841 = s3 ? tmp13842 : tmp13843;
  assign tmp13835 = s4 ? tmp13836 : tmp13841;
  assign tmp13847 = s2 ? tmp13822 : tmp13844;
  assign tmp13846 = s3 ? tmp13847 : tmp12966;
  assign tmp13849 = s2 ? 1 : tmp13791;
  assign tmp13848 = s3 ? tmp13849 : tmp12903;
  assign tmp13845 = s4 ? tmp13846 : tmp13848;
  assign tmp13834 = s5 ? tmp13835 : tmp13845;
  assign tmp13830 = s6 ? tmp13831 : tmp13834;
  assign tmp13786 = s7 ? tmp13787 : tmp13830;
  assign tmp13856 = s1 ? tmp13791 : tmp12904;
  assign tmp13855 = s2 ? tmp13856 : 1;
  assign tmp13854 = s3 ? tmp13814 : tmp13855;
  assign tmp13853 = s4 ? tmp13805 : tmp13854;
  assign tmp13859 = s2 ? tmp13184 : tmp13828;
  assign tmp13858 = s3 ? tmp13859 : tmp12946;
  assign tmp13857 = s4 ? tmp13820 : tmp13858;
  assign tmp13852 = s5 ? tmp13853 : tmp13857;
  assign tmp13851 = s6 ? tmp13788 : tmp13852;
  assign tmp13850 = s7 ? tmp13851 : tmp13830;
  assign tmp13785 = s8 ? tmp13786 : tmp13850;
  assign tmp13865 = ~(s2 ? tmp13081 : tmp13073);
  assign tmp13864 = s3 ? tmp13078 : tmp13865;
  assign tmp13863 = s4 ? tmp13069 : tmp13864;
  assign tmp13870 = ~(s1 ? tmp12994 : tmp13071);
  assign tmp13869 = ~(s2 ? tmp13090 : tmp13870);
  assign tmp13868 = s3 ? tmp13087 : tmp13869;
  assign tmp13867 = s4 ? tmp13868 : tmp13094;
  assign tmp13875 = s0 ? tmp13071 : tmp12905;
  assign tmp13874 = s1 ? tmp13875 : tmp12905;
  assign tmp13873 = s2 ? tmp13874 : tmp13071;
  assign tmp13872 = s3 ? tmp13873 : tmp13106;
  assign tmp13878 = s1 ? tmp12903 : tmp12905;
  assign tmp13880 = s0 ? tmp12905 : tmp13071;
  assign tmp13879 = s1 ? tmp13880 : tmp13071;
  assign tmp13877 = s2 ? tmp13878 : tmp13879;
  assign tmp13882 = s1 ? tmp12905 : tmp12918;
  assign tmp13881 = s2 ? tmp13882 : tmp12948;
  assign tmp13876 = s3 ? tmp13877 : tmp13881;
  assign tmp13871 = s4 ? tmp13872 : tmp13876;
  assign tmp13866 = s5 ? tmp13867 : tmp13871;
  assign tmp13862 = s6 ? tmp13863 : tmp13866;
  assign tmp13886 = ~(s2 ? tmp13114 : tmp13073);
  assign tmp13885 = s3 ? tmp13078 : tmp13886;
  assign tmp13884 = s4 ? tmp13069 : tmp13885;
  assign tmp13891 = s1 ? tmp12994 : tmp13071;
  assign tmp13890 = s2 ? tmp13071 : tmp13891;
  assign tmp13889 = s3 ? tmp13118 : tmp13890;
  assign tmp13888 = s4 ? tmp13889 : tmp13122;
  assign tmp13893 = s3 ? tmp13873 : tmp13226;
  assign tmp13895 = s2 ? tmp12905 : tmp13071;
  assign tmp13894 = s3 ? tmp13895 : tmp12903;
  assign tmp13892 = s4 ? tmp13893 : tmp13894;
  assign tmp13887 = s5 ? tmp13888 : tmp13892;
  assign tmp13883 = s6 ? tmp13884 : tmp13887;
  assign tmp13861 = s7 ? tmp13862 : tmp13883;
  assign tmp13860 = s8 ? tmp13850 : tmp13861;
  assign tmp13784 = s9 ? tmp13785 : tmp13860;
  assign tmp13904 = s0 ? tmp12905 : tmp13791;
  assign tmp13903 = ~(s1 ? tmp13791 : tmp13904);
  assign tmp13902 = ~(s2 ? tmp13081 : tmp13903);
  assign tmp13901 = s3 ? tmp13798 : tmp13902;
  assign tmp13900 = s4 ? tmp13789 : tmp13901;
  assign tmp13909 = ~(s1 ? tmp12994 : tmp13791);
  assign tmp13908 = ~(s2 ? tmp13809 : tmp13909);
  assign tmp13907 = s3 ? tmp13806 : tmp13908;
  assign tmp13906 = s4 ? tmp13907 : tmp13813;
  assign tmp13913 = s1 ? tmp13823 : tmp12905;
  assign tmp13914 = s1 ? tmp13904 : tmp13791;
  assign tmp13912 = s2 ? tmp13913 : tmp13914;
  assign tmp13911 = s3 ? tmp13912 : tmp13106;
  assign tmp13916 = s2 ? tmp13878 : tmp13828;
  assign tmp13915 = s3 ? tmp13916 : tmp13881;
  assign tmp13910 = s4 ? tmp13911 : tmp13915;
  assign tmp13905 = s5 ? tmp13906 : tmp13910;
  assign tmp13899 = s6 ? tmp13900 : tmp13905;
  assign tmp13920 = ~(s2 ? tmp13114 : tmp13903);
  assign tmp13919 = s3 ? tmp13798 : tmp13920;
  assign tmp13918 = s4 ? tmp13789 : tmp13919;
  assign tmp13925 = s1 ? tmp12994 : tmp13791;
  assign tmp13924 = s2 ? tmp13791 : tmp13925;
  assign tmp13923 = s3 ? tmp13837 : tmp13924;
  assign tmp13922 = s4 ? tmp13923 : tmp13841;
  assign tmp13928 = s2 ? tmp13913 : tmp13844;
  assign tmp13927 = s3 ? tmp13928 : tmp12966;
  assign tmp13930 = s2 ? tmp12905 : tmp13791;
  assign tmp13929 = s3 ? tmp13930 : tmp12903;
  assign tmp13926 = s4 ? tmp13927 : tmp13929;
  assign tmp13921 = s5 ? tmp13922 : tmp13926;
  assign tmp13917 = s6 ? tmp13918 : tmp13921;
  assign tmp13898 = s7 ? tmp13899 : tmp13917;
  assign tmp13897 = s8 ? tmp13898 : tmp13899;
  assign tmp13932 = s7 ? tmp13830 : tmp13883;
  assign tmp13931 = s8 ? tmp13932 : tmp13917;
  assign tmp13896 = s9 ? tmp13897 : tmp13931;
  assign tmp13783 = s10 ? tmp13784 : tmp13896;
  assign tmp13941 = s3 ? tmp13269 : tmp12966;
  assign tmp13940 = s4 ? tmp13941 : tmp13377;
  assign tmp13939 = s5 ? tmp13278 : tmp13940;
  assign tmp13938 = s6 ? tmp13274 : tmp13939;
  assign tmp13937 = s7 ? tmp13251 : tmp13938;
  assign tmp13946 = s3 ? tmp13350 : tmp12966;
  assign tmp13945 = s4 ? tmp13946 : tmp13382;
  assign tmp13944 = s5 ? tmp13339 : tmp13945;
  assign tmp13943 = s6 ? tmp13333 : tmp13944;
  assign tmp13942 = s7 ? tmp13287 : tmp13943;
  assign tmp13936 = s8 ? tmp13937 : tmp13942;
  assign tmp13947 = s8 ? tmp13942 : tmp13355;
  assign tmp13935 = s9 ? tmp13936 : tmp13947;
  assign tmp13952 = s5 ? tmp13363 : tmp13940;
  assign tmp13951 = s6 ? tmp13274 : tmp13952;
  assign tmp13950 = s7 ? tmp13356 : tmp13951;
  assign tmp13949 = s8 ? tmp13950 : tmp13356;
  assign tmp13957 = s4 ? tmp13367 : tmp13377;
  assign tmp13956 = s5 ? tmp13363 : tmp13957;
  assign tmp13955 = s6 ? tmp13274 : tmp13956;
  assign tmp13954 = s7 ? tmp13938 : tmp13955;
  assign tmp13958 = s7 ? tmp13943 : tmp13951;
  assign tmp13953 = s8 ? tmp13954 : tmp13958;
  assign tmp13948 = s9 ? tmp13949 : tmp13953;
  assign tmp13934 = s10 ? tmp13935 : tmp13948;
  assign tmp13962 = s7 ? tmp13938 : tmp13361;
  assign tmp13961 = s8 ? tmp13962 : tmp13958;
  assign tmp13960 = s9 ? tmp13949 : tmp13961;
  assign tmp13959 = s10 ? tmp13935 : tmp13960;
  assign tmp13933 = s11 ? tmp13934 : tmp13959;
  assign tmp13782 = ~(s12 ? tmp13783 : tmp13933);
  assign tmp13607 = s13 ? tmp13608 : tmp13782;
  assign tmp13606 = s14 ? 1 : tmp13607;
  assign tmp13977 = ~(s0 ? tmp13402 : tmp12931);
  assign tmp13976 = ~(s1 ? tmp13423 : tmp13977);
  assign tmp13975 = s2 ? tmp13421 : tmp13976;
  assign tmp13979 = s0 ? tmp12905 : tmp13406;
  assign tmp13978 = ~(s2 ? tmp13979 : tmp13426);
  assign tmp13974 = s3 ? tmp13975 : tmp13978;
  assign tmp13973 = s4 ? tmp13974 : tmp13427;
  assign tmp13972 = s5 ? tmp13973 : tmp13433;
  assign tmp13971 = s6 ? tmp13399 : tmp13972;
  assign tmp13986 = s0 ? tmp13402 : tmp12931;
  assign tmp13985 = s1 ? tmp13402 : tmp13986;
  assign tmp13984 = s2 ? tmp13456 : tmp13985;
  assign tmp13983 = s3 ? tmp13984 : tmp13458;
  assign tmp13982 = s4 ? tmp13983 : tmp13460;
  assign tmp13989 = s2 ? 1 : tmp13467;
  assign tmp13988 = s3 ? tmp13465 : tmp13989;
  assign tmp13991 = s2 ? tmp13314 : tmp13402;
  assign tmp13990 = s3 ? tmp13991 : tmp13467;
  assign tmp13987 = s4 ? tmp13988 : tmp13990;
  assign tmp13981 = s5 ? tmp13982 : tmp13987;
  assign tmp13980 = s6 ? tmp13447 : tmp13981;
  assign tmp13970 = s7 ? tmp13971 : tmp13980;
  assign tmp13997 = s1 ? tmp13416 : tmp13402;
  assign tmp13996 = s2 ? tmp13997 : tmp13459;
  assign tmp13995 = s3 ? tmp13401 : tmp13996;
  assign tmp13994 = s4 ? tmp13995 : tmp13409;
  assign tmp13993 = s6 ? tmp13994 : tmp13476;
  assign tmp13999 = s4 ? tmp13995 : tmp13448;
  assign tmp14002 = s3 ? tmp13509 : tmp13989;
  assign tmp14004 = s2 ? 1 : tmp13402;
  assign tmp14003 = s3 ? tmp14004 : tmp13467;
  assign tmp14001 = s4 ? tmp14002 : tmp14003;
  assign tmp14000 = s5 ? tmp13498 : tmp14001;
  assign tmp13998 = s6 ? tmp13999 : tmp14000;
  assign tmp13992 = s7 ? tmp13993 : tmp13998;
  assign tmp13969 = s8 ? tmp13970 : tmp13992;
  assign tmp14011 = s2 ? tmp13522 : tmp13309;
  assign tmp14012 = s2 ? tmp13313 : tmp13295;
  assign tmp14010 = s3 ? tmp14011 : tmp14012;
  assign tmp14009 = s4 ? tmp14010 : tmp13526;
  assign tmp14008 = s5 ? tmp14009 : tmp13531;
  assign tmp14007 = s6 ? tmp13515 : tmp14008;
  assign tmp14017 = s2 ? tmp13548 : tmp13342;
  assign tmp14016 = s3 ? tmp14017 : tmp13294;
  assign tmp14015 = s4 ? tmp14016 : tmp13550;
  assign tmp14014 = s5 ? tmp14015 : tmp13553;
  assign tmp14013 = s6 ? tmp13543 : tmp14014;
  assign tmp14006 = s7 ? tmp14007 : tmp14013;
  assign tmp14005 = s8 ? tmp13992 : tmp14006;
  assign tmp13968 = s9 ? tmp13969 : tmp14005;
  assign tmp14025 = s2 ? tmp13421 : tmp13481;
  assign tmp14026 = s2 ? tmp13430 : tmp13459;
  assign tmp14024 = s3 ? tmp14025 : tmp14026;
  assign tmp14023 = s4 ? tmp14024 : tmp13427;
  assign tmp14022 = s5 ? tmp14023 : tmp13433;
  assign tmp14021 = s6 ? tmp13399 : tmp14022;
  assign tmp14031 = s2 ? tmp13456 : tmp13502;
  assign tmp14030 = s3 ? tmp14031 : tmp13458;
  assign tmp14029 = s4 ? tmp14030 : tmp13579;
  assign tmp14028 = s5 ? tmp14029 : tmp13987;
  assign tmp14027 = s6 ? tmp13447 : tmp14028;
  assign tmp14020 = s7 ? tmp14021 : tmp14027;
  assign tmp14019 = s8 ? tmp14020 : tmp14021;
  assign tmp14036 = s4 ? tmp13983 : tmp13586;
  assign tmp14035 = s5 ? tmp14036 : tmp13987;
  assign tmp14034 = s6 ? tmp13447 : tmp14035;
  assign tmp14038 = s5 ? tmp14015 : tmp13591;
  assign tmp14037 = s6 ? tmp13543 : tmp14038;
  assign tmp14033 = s7 ? tmp14034 : tmp14037;
  assign tmp14039 = s7 ? tmp13998 : tmp14027;
  assign tmp14032 = s8 ? tmp14033 : tmp14039;
  assign tmp14018 = s9 ? tmp14019 : tmp14032;
  assign tmp13967 = s10 ? tmp13968 : tmp14018;
  assign tmp14043 = s7 ? tmp13980 : tmp14013;
  assign tmp14042 = s8 ? tmp14043 : tmp14039;
  assign tmp14041 = s9 ? tmp14019 : tmp14042;
  assign tmp14040 = s10 ? tmp13968 : tmp14041;
  assign tmp13966 = s11 ? tmp13967 : tmp14040;
  assign tmp14053 = s1 ? tmp13006 : 1;
  assign tmp14052 = s2 ? tmp14053 : 1;
  assign tmp14051 = s3 ? tmp14052 : 1;
  assign tmp14050 = s4 ? 1 : tmp14051;
  assign tmp14059 = s0 ? 1 : tmp13824;
  assign tmp14058 = s1 ? tmp14059 : 1;
  assign tmp14061 = s0 ? tmp13824 : 1;
  assign tmp14060 = s1 ? tmp14061 : 1;
  assign tmp14057 = s2 ? tmp14058 : tmp14060;
  assign tmp14056 = s3 ? tmp14057 : 1;
  assign tmp14064 = s1 ? 1 : tmp12994;
  assign tmp14065 = s1 ? tmp12994 : tmp13006;
  assign tmp14063 = s2 ? tmp14064 : tmp14065;
  assign tmp14062 = s3 ? tmp14063 : 1;
  assign tmp14055 = s4 ? tmp14056 : tmp14062;
  assign tmp14054 = s5 ? tmp14055 : 1;
  assign tmp14049 = s6 ? tmp14050 : tmp14054;
  assign tmp14070 = s2 ? tmp14058 : 1;
  assign tmp14069 = s3 ? tmp14070 : 1;
  assign tmp14072 = s2 ? tmp14064 : 1;
  assign tmp14071 = s3 ? tmp14072 : 1;
  assign tmp14068 = s4 ? tmp14069 : tmp14071;
  assign tmp14067 = s5 ? tmp14068 : 1;
  assign tmp14066 = s6 ? tmp14050 : tmp14067;
  assign tmp14048 = s7 ? tmp14049 : tmp14066;
  assign tmp14078 = ~(l2 ? tmp13624 : 0);
  assign tmp14077 = l1 ? 1 : tmp14078;
  assign tmp14081 = s0 ? 1 : tmp14077;
  assign tmp14080 = s1 ? tmp14081 : tmp14077;
  assign tmp14079 = s2 ? tmp14080 : tmp14077;
  assign tmp14076 = s3 ? tmp14077 : tmp14079;
  assign tmp14085 = s0 ? tmp14077 : 0;
  assign tmp14084 = s1 ? tmp14085 : tmp14077;
  assign tmp14086 = s0 ? tmp14077 : 1;
  assign tmp14083 = s2 ? tmp14084 : tmp14086;
  assign tmp14088 = s1 ? tmp13624 : 0;
  assign tmp14089 = ~(l1 ? 1 : tmp14078);
  assign tmp14087 = ~(s2 ? tmp14088 : tmp14089);
  assign tmp14082 = s3 ? tmp14083 : tmp14087;
  assign tmp14075 = s4 ? tmp14076 : tmp14082;
  assign tmp14095 = s0 ? tmp14077 : tmp13824;
  assign tmp14094 = s1 ? tmp14095 : 1;
  assign tmp14097 = s0 ? tmp13824 : tmp14077;
  assign tmp14096 = s1 ? tmp14097 : tmp14077;
  assign tmp14093 = s2 ? tmp14094 : tmp14096;
  assign tmp14101 = l1 ? 1 : tmp13404;
  assign tmp14100 = s0 ? tmp14101 : 1;
  assign tmp14099 = s1 ? tmp14100 : tmp14077;
  assign tmp14098 = s2 ? tmp14077 : tmp14099;
  assign tmp14092 = s3 ? tmp14093 : tmp14098;
  assign tmp14105 = ~(s0 ? 1 : tmp13624);
  assign tmp14104 = s1 ? tmp14081 : tmp14105;
  assign tmp14107 = s0 ? 1 : tmp13624;
  assign tmp14108 = ~(s0 ? tmp14077 : 0);
  assign tmp14106 = ~(s1 ? tmp14107 : tmp14108);
  assign tmp14103 = s2 ? tmp14104 : tmp14106;
  assign tmp14111 = ~(s0 ? tmp13624 : 0);
  assign tmp14110 = s1 ? tmp14077 : tmp14111;
  assign tmp14109 = s2 ? tmp14110 : 1;
  assign tmp14102 = s3 ? tmp14103 : tmp14109;
  assign tmp14091 = s4 ? tmp14092 : tmp14102;
  assign tmp14116 = s0 ? 1 : tmp14101;
  assign tmp14115 = s1 ? tmp14086 : tmp14116;
  assign tmp14117 = s1 ? tmp14100 : 1;
  assign tmp14114 = s2 ? tmp14115 : tmp14117;
  assign tmp14113 = s3 ? tmp14114 : 1;
  assign tmp14120 = s1 ? 1 : tmp14116;
  assign tmp14121 = s1 ? tmp14081 : 1;
  assign tmp14119 = s2 ? tmp14120 : tmp14121;
  assign tmp14122 = s2 ? tmp14117 : 1;
  assign tmp14118 = s3 ? tmp14119 : tmp14122;
  assign tmp14112 = s4 ? tmp14113 : tmp14118;
  assign tmp14090 = s5 ? tmp14091 : tmp14112;
  assign tmp14074 = s6 ? tmp14075 : tmp14090;
  assign tmp14127 = s2 ? tmp14094 : tmp14077;
  assign tmp14126 = s3 ? tmp14127 : tmp14098;
  assign tmp14129 = s2 ? tmp14104 : tmp14077;
  assign tmp14131 = s1 ? tmp14077 : 1;
  assign tmp14130 = s2 ? tmp14131 : 1;
  assign tmp14128 = s3 ? tmp14129 : tmp14130;
  assign tmp14125 = s4 ? tmp14126 : tmp14128;
  assign tmp14135 = s1 ? tmp14086 : tmp14101;
  assign tmp14134 = s2 ? tmp14135 : tmp14117;
  assign tmp14133 = s3 ? tmp14134 : 1;
  assign tmp14138 = s1 ? 1 : tmp14101;
  assign tmp14137 = s2 ? tmp14138 : tmp14077;
  assign tmp14136 = s3 ? tmp14137 : tmp14117;
  assign tmp14132 = s4 ? tmp14133 : tmp14136;
  assign tmp14124 = s5 ? tmp14125 : tmp14132;
  assign tmp14123 = s6 ? tmp14075 : tmp14124;
  assign tmp14073 = s7 ? tmp14074 : tmp14123;
  assign tmp14047 = s8 ? tmp14048 : tmp14073;
  assign tmp14145 = s1 ? tmp14095 : tmp14077;
  assign tmp14144 = s2 ? tmp14145 : tmp14086;
  assign tmp14143 = s3 ? tmp14144 : tmp14087;
  assign tmp14142 = s4 ? tmp14076 : tmp14143;
  assign tmp14151 = ~(s0 ? tmp14077 : tmp13824);
  assign tmp14150 = ~(s1 ? tmp14107 : tmp14151);
  assign tmp14149 = s2 ? tmp14104 : tmp14150;
  assign tmp14148 = s3 ? tmp14149 : tmp14109;
  assign tmp14147 = s4 ? tmp14092 : tmp14148;
  assign tmp14146 = s5 ? tmp14147 : tmp14112;
  assign tmp14141 = s6 ? tmp14142 : tmp14146;
  assign tmp14152 = s6 ? tmp14142 : tmp14124;
  assign tmp14140 = s7 ? tmp14141 : tmp14152;
  assign tmp14159 = s0 ? tmp14101 : tmp12905;
  assign tmp14158 = s1 ? tmp14159 : tmp14101;
  assign tmp14157 = s2 ? tmp14158 : tmp14100;
  assign tmp14161 = ~(l1 ? 1 : tmp13404);
  assign tmp14160 = ~(s2 ? tmp14088 : tmp14161);
  assign tmp14156 = s3 ? tmp14157 : tmp14160;
  assign tmp14155 = s4 ? tmp14101 : tmp14156;
  assign tmp14166 = s1 ? tmp14159 : tmp12905;
  assign tmp14168 = s0 ? tmp12905 : tmp14101;
  assign tmp14167 = s1 ? tmp14168 : tmp14101;
  assign tmp14165 = s2 ? tmp14166 : tmp14167;
  assign tmp14170 = s1 ? tmp14100 : tmp14101;
  assign tmp14169 = s2 ? tmp14101 : tmp14170;
  assign tmp14164 = s3 ? tmp14165 : tmp14169;
  assign tmp14173 = s1 ? tmp14116 : tmp14105;
  assign tmp14175 = ~(s0 ? tmp14101 : tmp12905);
  assign tmp14174 = ~(s1 ? tmp14107 : tmp14175);
  assign tmp14172 = s2 ? tmp14173 : tmp14174;
  assign tmp14177 = s1 ? tmp14101 : tmp14111;
  assign tmp14176 = s2 ? tmp14177 : 1;
  assign tmp14171 = s3 ? tmp14172 : tmp14176;
  assign tmp14163 = s4 ? tmp14164 : tmp14171;
  assign tmp14181 = s1 ? tmp14100 : tmp14116;
  assign tmp14182 = s1 ? tmp14101 : tmp13006;
  assign tmp14180 = s2 ? tmp14181 : tmp14182;
  assign tmp14179 = s3 ? tmp14180 : 1;
  assign tmp14185 = s1 ? tmp14116 : tmp12994;
  assign tmp14184 = s2 ? tmp14120 : tmp14185;
  assign tmp14183 = s3 ? tmp14184 : tmp14122;
  assign tmp14178 = s4 ? tmp14179 : tmp14183;
  assign tmp14162 = s5 ? tmp14163 : tmp14178;
  assign tmp14154 = s6 ? tmp14155 : tmp14162;
  assign tmp14190 = s2 ? tmp14166 : tmp14101;
  assign tmp14189 = s3 ? tmp14190 : tmp14169;
  assign tmp14192 = s2 ? tmp14173 : tmp14101;
  assign tmp14194 = s1 ? tmp14101 : 1;
  assign tmp14193 = s2 ? tmp14194 : 1;
  assign tmp14191 = s3 ? tmp14192 : tmp14193;
  assign tmp14188 = s4 ? tmp14189 : tmp14191;
  assign tmp14197 = s2 ? tmp14170 : tmp14194;
  assign tmp14196 = s3 ? tmp14197 : 1;
  assign tmp14199 = s2 ? tmp14138 : tmp14101;
  assign tmp14198 = s3 ? tmp14199 : tmp14117;
  assign tmp14195 = s4 ? tmp14196 : tmp14198;
  assign tmp14187 = s5 ? tmp14188 : tmp14195;
  assign tmp14186 = s6 ? tmp14155 : tmp14187;
  assign tmp14153 = s7 ? tmp14154 : tmp14186;
  assign tmp14139 = s8 ? tmp14140 : tmp14153;
  assign tmp14046 = s9 ? tmp14047 : tmp14139;
  assign tmp14204 = s4 ? tmp14077 : tmp14143;
  assign tmp14209 = s1 ? tmp14095 : tmp13824;
  assign tmp14208 = s2 ? tmp14209 : tmp14096;
  assign tmp14207 = s3 ? tmp14208 : tmp14098;
  assign tmp14206 = s4 ? tmp14207 : tmp14148;
  assign tmp14213 = s1 ? tmp14077 : tmp14059;
  assign tmp14212 = s2 ? tmp14115 : tmp14213;
  assign tmp14211 = s3 ? tmp14212 : 1;
  assign tmp14216 = s1 ? tmp14081 : tmp14061;
  assign tmp14215 = s2 ? tmp14120 : tmp14216;
  assign tmp14214 = s3 ? tmp14215 : tmp14122;
  assign tmp14210 = s4 ? tmp14211 : tmp14214;
  assign tmp14205 = s5 ? tmp14206 : tmp14210;
  assign tmp14203 = s6 ? tmp14204 : tmp14205;
  assign tmp14221 = s2 ? tmp14209 : tmp14077;
  assign tmp14220 = s3 ? tmp14221 : tmp14098;
  assign tmp14219 = s4 ? tmp14220 : tmp14128;
  assign tmp14224 = s2 ? tmp14135 : tmp14131;
  assign tmp14223 = s3 ? tmp14224 : 1;
  assign tmp14222 = s4 ? tmp14223 : tmp14136;
  assign tmp14218 = s5 ? tmp14219 : tmp14222;
  assign tmp14217 = s6 ? tmp14204 : tmp14218;
  assign tmp14202 = s7 ? tmp14203 : tmp14217;
  assign tmp14201 = s8 ? tmp14202 : tmp14203;
  assign tmp14230 = s3 ? tmp14199 : 1;
  assign tmp14229 = s4 ? tmp14196 : tmp14230;
  assign tmp14228 = s5 ? tmp14188 : tmp14229;
  assign tmp14227 = s6 ? tmp14155 : tmp14228;
  assign tmp14226 = s7 ? tmp14066 : tmp14227;
  assign tmp14234 = s3 ? tmp14137 : 1;
  assign tmp14233 = s4 ? tmp14223 : tmp14234;
  assign tmp14232 = s5 ? tmp14219 : tmp14233;
  assign tmp14231 = s6 ? tmp14204 : tmp14232;
  assign tmp14225 = s8 ? tmp14226 : tmp14231;
  assign tmp14200 = s9 ? tmp14201 : tmp14225;
  assign tmp14045 = s10 ? tmp14046 : tmp14200;
  assign tmp14238 = s7 ? tmp14066 : tmp14186;
  assign tmp14237 = s8 ? tmp14238 : tmp14217;
  assign tmp14236 = s9 ? tmp14201 : tmp14237;
  assign tmp14235 = s10 ? tmp14046 : tmp14236;
  assign tmp14044 = s11 ? tmp14045 : tmp14235;
  assign tmp13965 = s12 ? tmp13966 : tmp14044;
  assign tmp13964 = s13 ? tmp13965 : 1;
  assign tmp13963 = ~(s14 ? 1 : tmp13964);
  assign tmp13605 = s15 ? tmp13606 : tmp13963;
  assign tmp12889 = s16 ? tmp12890 : tmp13605;
  assign tmp14254 = s1 ? tmp13006 : tmp12994;
  assign tmp14253 = s2 ? tmp13004 : tmp14254;
  assign tmp14255 = s2 ? tmp13006 : tmp13008;
  assign tmp14252 = s3 ? tmp14253 : tmp14255;
  assign tmp14251 = s4 ? tmp14252 : tmp13009;
  assign tmp14250 = s5 ? tmp14251 : tmp13014;
  assign tmp14249 = s6 ? tmp12990 : tmp14250;
  assign tmp14261 = s1 ? tmp12905 : tmp12994;
  assign tmp14260 = s2 ? tmp13004 : tmp14261;
  assign tmp14259 = s3 ? tmp14260 : tmp13007;
  assign tmp14258 = s4 ? tmp14259 : tmp13009;
  assign tmp14257 = s5 ? tmp14258 : tmp13036;
  assign tmp14256 = s6 ? tmp13029 : tmp14257;
  assign tmp14248 = s7 ? tmp14249 : tmp14256;
  assign tmp14247 = ~(s8 ? tmp13702 : tmp14248);
  assign tmp14246 = s9 ? tmp13612 : tmp14247;
  assign tmp14263 = s8 ? tmp12969 : tmp12970;
  assign tmp14266 = ~(s6 ? tmp13029 : tmp14257);
  assign tmp14265 = s7 ? tmp13761 : tmp14266;
  assign tmp14268 = s6 ? tmp13678 : tmp13771;
  assign tmp14269 = ~(s6 ? tmp12950 : tmp12979);
  assign tmp14267 = ~(s7 ? tmp14268 : tmp14269);
  assign tmp14264 = s8 ? tmp14265 : tmp14267;
  assign tmp14262 = s9 ? tmp14263 : tmp14264;
  assign tmp14245 = s10 ? tmp14246 : tmp14262;
  assign tmp14273 = s7 ? tmp13614 : tmp14266;
  assign tmp14274 = ~(s7 ? tmp13677 : tmp14269);
  assign tmp14272 = s8 ? tmp14273 : tmp14274;
  assign tmp14271 = s9 ? tmp14263 : tmp14272;
  assign tmp14270 = s10 ? tmp14246 : tmp14271;
  assign tmp14244 = ~(s11 ? tmp14245 : tmp14270);
  assign tmp14243 = s12 ? 1 : tmp14244;
  assign tmp14285 = s1 ? tmp13880 : 0;
  assign tmp14284 = s2 ? tmp14285 : tmp13097;
  assign tmp14283 = s3 ? tmp14284 : tmp13098;
  assign tmp14282 = s4 ? tmp13086 : tmp14283;
  assign tmp14289 = s1 ? tmp13875 : 1;
  assign tmp14288 = s2 ? tmp14289 : tmp13071;
  assign tmp14287 = s3 ? tmp14288 : tmp13106;
  assign tmp14291 = s2 ? tmp12903 : tmp13879;
  assign tmp14290 = s3 ? tmp14291 : tmp12946;
  assign tmp14286 = s4 ? tmp14287 : tmp14290;
  assign tmp14281 = s5 ? tmp14282 : tmp14286;
  assign tmp14280 = s6 ? tmp13068 : tmp14281;
  assign tmp14296 = s2 ? tmp14285 : tmp13071;
  assign tmp14295 = s3 ? tmp14296 : tmp13124;
  assign tmp14294 = s4 ? tmp13117 : tmp14295;
  assign tmp14298 = s3 ? tmp14288 : tmp13128;
  assign tmp14297 = s4 ? tmp14298 : tmp13129;
  assign tmp14293 = s5 ? tmp14294 : tmp14297;
  assign tmp14292 = s6 ? tmp13111 : tmp14293;
  assign tmp14279 = s7 ? tmp14280 : tmp14292;
  assign tmp14305 = s1 ? tmp13071 : tmp12904;
  assign tmp14304 = s2 ? tmp14305 : 1;
  assign tmp14303 = s3 ? tmp14284 : tmp14304;
  assign tmp14302 = s4 ? tmp13086 : tmp14303;
  assign tmp14308 = s2 ? tmp14289 : tmp13109;
  assign tmp14307 = s3 ? tmp14308 : tmp13106;
  assign tmp14310 = s2 ? tmp13184 : tmp13879;
  assign tmp14309 = s3 ? tmp14310 : tmp12946;
  assign tmp14306 = s4 ? tmp14307 : tmp14309;
  assign tmp14301 = s5 ? tmp14302 : tmp14306;
  assign tmp14300 = s6 ? tmp13068 : tmp14301;
  assign tmp14299 = s7 ? tmp14300 : tmp14292;
  assign tmp14278 = s8 ? tmp14279 : tmp14299;
  assign tmp14317 = s2 ? tmp14289 : tmp13219;
  assign tmp14316 = s3 ? tmp14317 : tmp13106;
  assign tmp14315 = s4 ? tmp14316 : tmp14290;
  assign tmp14314 = s5 ? tmp14282 : tmp14315;
  assign tmp14313 = s6 ? tmp13068 : tmp14314;
  assign tmp14322 = s2 ? tmp14289 : tmp13125;
  assign tmp14321 = s3 ? tmp14322 : tmp13226;
  assign tmp14320 = s4 ? tmp14321 : tmp13129;
  assign tmp14319 = s5 ? tmp14294 : tmp14320;
  assign tmp14318 = s6 ? tmp13111 : tmp14319;
  assign tmp14312 = s7 ? tmp14313 : tmp14318;
  assign tmp14311 = s8 ? tmp14299 : tmp14312;
  assign tmp14277 = s9 ? tmp14278 : tmp14311;
  assign tmp14329 = s3 ? tmp14322 : tmp13128;
  assign tmp14328 = s4 ? tmp14329 : tmp13129;
  assign tmp14327 = s5 ? tmp14294 : tmp14328;
  assign tmp14326 = s6 ? tmp13111 : tmp14327;
  assign tmp14325 = s7 ? tmp14280 : tmp14326;
  assign tmp14324 = s8 ? tmp14325 : tmp14280;
  assign tmp14330 = s7 ? tmp14292 : tmp14326;
  assign tmp14323 = s9 ? tmp14324 : tmp14330;
  assign tmp14276 = s10 ? tmp14277 : tmp14323;
  assign tmp14275 = ~(s12 ? tmp14276 : tmp13246);
  assign tmp14242 = s13 ? tmp14243 : tmp14275;
  assign tmp14241 = s14 ? 1 : tmp14242;
  assign tmp14343 = s2 ? tmp14053 : tmp13004;
  assign tmp14342 = s3 ? tmp14343 : 1;
  assign tmp14341 = s4 ? tmp14342 : tmp14062;
  assign tmp14340 = s5 ? tmp14341 : 1;
  assign tmp14339 = s6 ? tmp14050 : tmp14340;
  assign tmp14346 = s4 ? tmp14051 : tmp14071;
  assign tmp14345 = s5 ? tmp14346 : 1;
  assign tmp14344 = s6 ? tmp14050 : tmp14345;
  assign tmp14338 = s7 ? tmp14339 : tmp14344;
  assign tmp14337 = s8 ? tmp14140 : tmp14338;
  assign tmp14336 = s9 ? tmp14047 : tmp14337;
  assign tmp14351 = s4 ? 1 : tmp14069;
  assign tmp14356 = s1 ? tmp12994 : tmp14059;
  assign tmp14355 = s2 ? tmp14064 : tmp14356;
  assign tmp14354 = s3 ? tmp14355 : 1;
  assign tmp14353 = s4 ? tmp14056 : tmp14354;
  assign tmp14352 = s5 ? tmp14353 : 1;
  assign tmp14350 = s6 ? tmp14351 : tmp14352;
  assign tmp14357 = s6 ? tmp14351 : tmp14067;
  assign tmp14349 = s7 ? tmp14350 : tmp14357;
  assign tmp14348 = s8 ? tmp14349 : tmp14350;
  assign tmp14359 = s7 ? tmp14066 : tmp14344;
  assign tmp14363 = s4 ? tmp14133 : tmp14234;
  assign tmp14362 = s5 ? tmp14125 : tmp14363;
  assign tmp14361 = s6 ? tmp14142 : tmp14362;
  assign tmp14360 = s7 ? tmp14361 : tmp14357;
  assign tmp14358 = s8 ? tmp14359 : tmp14360;
  assign tmp14347 = s9 ? tmp14348 : tmp14358;
  assign tmp14335 = s10 ? tmp14336 : tmp14347;
  assign tmp14367 = s7 ? tmp14152 : tmp14357;
  assign tmp14366 = s8 ? tmp14359 : tmp14367;
  assign tmp14365 = s9 ? tmp14348 : tmp14366;
  assign tmp14364 = s10 ? tmp14336 : tmp14365;
  assign tmp14334 = s11 ? tmp14335 : tmp14364;
  assign tmp14333 = s12 ? tmp13393 : tmp14334;
  assign tmp14332 = s13 ? tmp14333 : 1;
  assign tmp14331 = ~(s14 ? 1 : tmp14332);
  assign tmp14240 = s15 ? tmp14241 : tmp14331;
  assign tmp14380 = ~(s1 ? tmp13071 : tmp13880);
  assign tmp14379 = ~(s2 ? tmp13081 : tmp14380);
  assign tmp14378 = s3 ? tmp13078 : tmp14379;
  assign tmp14377 = s4 ? tmp13069 : tmp14378;
  assign tmp14382 = s4 ? tmp13868 : tmp14283;
  assign tmp14386 = s1 ? tmp12903 : tmp13071;
  assign tmp14385 = s2 ? tmp14386 : tmp13879;
  assign tmp14384 = s3 ? tmp14385 : tmp13881;
  assign tmp14383 = s4 ? tmp13872 : tmp14384;
  assign tmp14381 = s5 ? tmp14382 : tmp14383;
  assign tmp14376 = s6 ? tmp14377 : tmp14381;
  assign tmp14390 = ~(s2 ? tmp13114 : tmp14380);
  assign tmp14389 = s3 ? tmp13078 : tmp14390;
  assign tmp14388 = s4 ? tmp13069 : tmp14389;
  assign tmp14392 = s4 ? tmp13889 : tmp14295;
  assign tmp14394 = s3 ? tmp13873 : tmp13128;
  assign tmp14393 = s4 ? tmp14394 : tmp13894;
  assign tmp14391 = s5 ? tmp14392 : tmp14393;
  assign tmp14387 = s6 ? tmp14388 : tmp14391;
  assign tmp14375 = s7 ? tmp14376 : tmp14387;
  assign tmp14400 = s2 ? tmp13874 : tmp13879;
  assign tmp14399 = s3 ? tmp14400 : tmp13106;
  assign tmp14398 = s4 ? tmp14399 : tmp13876;
  assign tmp14397 = s5 ? tmp14382 : tmp14398;
  assign tmp14396 = s6 ? tmp14377 : tmp14397;
  assign tmp14395 = s7 ? tmp14396 : tmp14387;
  assign tmp14374 = s8 ? tmp14375 : tmp14395;
  assign tmp14373 = s9 ? tmp14374 : tmp14395;
  assign tmp14402 = s8 ? tmp14395 : tmp14396;
  assign tmp14401 = s9 ? tmp14402 : tmp14387;
  assign tmp14372 = s10 ? tmp14373 : tmp14401;
  assign tmp14371 = ~(s12 ? tmp14372 : tmp13246);
  assign tmp14370 = s13 ? tmp13608 : tmp14371;
  assign tmp14369 = s14 ? 1 : tmp14370;
  assign tmp14405 = s12 ? tmp13393 : tmp14044;
  assign tmp14404 = s13 ? tmp14405 : 1;
  assign tmp14403 = ~(s14 ? 1 : tmp14404);
  assign tmp14368 = s15 ? tmp14369 : tmp14403;
  assign tmp14239 = s16 ? tmp14240 : tmp14368;
  assign tmp12888 = s17 ? tmp12889 : tmp14239;
  assign l4__1 = tmp12888;

  assign s18n = 0;

  assign tmp14422 = l2 ? 1 : 0;
  assign tmp14421 = l1 ? 1 : tmp14422;
  assign tmp14420 = s0 ? 1 : tmp14421;
  assign tmp14425 = s0 ? tmp14421 : 1;
  assign tmp14424 = s1 ? tmp14425 : tmp14421;
  assign tmp14423 = s2 ? tmp14421 : tmp14424;
  assign tmp14419 = s3 ? tmp14420 : tmp14423;
  assign tmp14428 = s1 ? tmp14425 : 1;
  assign tmp14427 = s2 ? tmp14424 : tmp14428;
  assign tmp14430 = s1 ? tmp14421 : tmp14420;
  assign tmp14429 = s2 ? 1 : tmp14430;
  assign tmp14426 = s3 ? tmp14427 : tmp14429;
  assign tmp14418 = s4 ? tmp14419 : tmp14426;
  assign tmp14435 = s1 ? tmp14425 : tmp14420;
  assign tmp14436 = s1 ? tmp14420 : tmp14425;
  assign tmp14434 = s2 ? tmp14435 : tmp14436;
  assign tmp14440 = l1 ? 1 : 0;
  assign tmp14439 = s0 ? tmp14421 : tmp14440;
  assign tmp14438 = s1 ? 1 : tmp14439;
  assign tmp14437 = s2 ? tmp14420 : tmp14438;
  assign tmp14433 = s3 ? tmp14434 : tmp14437;
  assign tmp14444 = s0 ? 1 : tmp14440;
  assign tmp14443 = s1 ? tmp14420 : tmp14444;
  assign tmp14445 = s1 ? tmp14444 : tmp14425;
  assign tmp14442 = s2 ? tmp14443 : tmp14445;
  assign tmp14447 = s1 ? tmp14439 : 1;
  assign tmp14446 = s2 ? tmp14447 : 1;
  assign tmp14441 = s3 ? tmp14442 : tmp14446;
  assign tmp14432 = s4 ? tmp14433 : tmp14441;
  assign tmp14452 = s0 ? tmp14440 : tmp14421;
  assign tmp14451 = s1 ? tmp14420 : tmp14452;
  assign tmp14450 = s2 ? tmp14428 : tmp14451;
  assign tmp14449 = s3 ? tmp14450 : 1;
  assign tmp14455 = s1 ? tmp14420 : tmp14439;
  assign tmp14454 = s2 ? 1 : tmp14455;
  assign tmp14453 = s3 ? tmp14454 : 1;
  assign tmp14448 = s4 ? tmp14449 : tmp14453;
  assign tmp14431 = s5 ? tmp14432 : tmp14448;
  assign tmp14417 = s6 ? tmp14418 : tmp14431;
  assign tmp14461 = s1 ? tmp14421 : tmp14425;
  assign tmp14460 = s2 ? tmp14424 : tmp14461;
  assign tmp14462 = s2 ? tmp14421 : tmp14438;
  assign tmp14459 = s3 ? tmp14460 : tmp14462;
  assign tmp14464 = s2 ? tmp14443 : tmp14421;
  assign tmp14463 = s3 ? tmp14464 : tmp14446;
  assign tmp14458 = s4 ? tmp14459 : tmp14463;
  assign tmp14468 = s1 ? tmp14421 : tmp14452;
  assign tmp14467 = s2 ? tmp14428 : tmp14468;
  assign tmp14471 = s0 ? tmp14440 : 1;
  assign tmp14470 = s1 ? tmp14471 : 1;
  assign tmp14469 = s2 ? tmp14470 : 1;
  assign tmp14466 = s3 ? tmp14467 : tmp14469;
  assign tmp14474 = s1 ? tmp14421 : tmp14439;
  assign tmp14473 = s2 ? 1 : tmp14474;
  assign tmp14472 = s3 ? tmp14473 : 1;
  assign tmp14465 = s4 ? tmp14466 : tmp14472;
  assign tmp14457 = s5 ? tmp14458 : tmp14465;
  assign tmp14456 = s6 ? tmp14418 : tmp14457;
  assign tmp14416 = s7 ? tmp14417 : tmp14456;
  assign tmp14479 = s3 ? 1 : tmp14469;
  assign tmp14482 = s1 ? 1 : tmp14440;
  assign tmp14481 = s2 ? 1 : tmp14482;
  assign tmp14480 = s3 ? tmp14481 : 1;
  assign tmp14478 = s4 ? tmp14479 : tmp14480;
  assign tmp14477 = s5 ? 1 : tmp14478;
  assign tmp14476 = s6 ? 1 : tmp14477;
  assign tmp14475 = s7 ? 1 : tmp14476;
  assign tmp14415 = s8 ? tmp14416 : tmp14475;
  assign tmp14490 = s1 ? 1 : tmp14420;
  assign tmp14489 = s2 ? 1 : tmp14490;
  assign tmp14488 = s3 ? 1 : tmp14489;
  assign tmp14493 = s1 ? 1 : tmp14444;
  assign tmp14494 = s1 ? tmp14444 : 1;
  assign tmp14492 = s2 ? tmp14493 : tmp14494;
  assign tmp14496 = s1 ? tmp14420 : 1;
  assign tmp14495 = s2 ? tmp14496 : 1;
  assign tmp14491 = s3 ? tmp14492 : tmp14495;
  assign tmp14487 = s4 ? tmp14488 : tmp14491;
  assign tmp14500 = s1 ? 1 : tmp14425;
  assign tmp14499 = s2 ? 1 : tmp14500;
  assign tmp14498 = s3 ? tmp14499 : 1;
  assign tmp14501 = s3 ? tmp14489 : 1;
  assign tmp14497 = s4 ? tmp14498 : tmp14501;
  assign tmp14486 = s5 ? tmp14487 : tmp14497;
  assign tmp14485 = s6 ? 1 : tmp14486;
  assign tmp14506 = s2 ? tmp14493 : 1;
  assign tmp14505 = s3 ? tmp14506 : tmp14495;
  assign tmp14504 = s4 ? tmp14488 : tmp14505;
  assign tmp14510 = s1 ? 1 : tmp14421;
  assign tmp14509 = s2 ? 1 : tmp14510;
  assign tmp14508 = s3 ? tmp14509 : 1;
  assign tmp14507 = s4 ? 1 : tmp14508;
  assign tmp14503 = s5 ? tmp14504 : tmp14507;
  assign tmp14502 = s6 ? 1 : tmp14503;
  assign tmp14484 = s7 ? tmp14485 : tmp14502;
  assign tmp14483 = s8 ? tmp14475 : tmp14484;
  assign tmp14414 = s9 ? tmp14415 : tmp14483;
  assign tmp14519 = s1 ? tmp14421 : 1;
  assign tmp14518 = s2 ? tmp14428 : tmp14519;
  assign tmp14517 = s3 ? tmp14518 : tmp14469;
  assign tmp14522 = s1 ? tmp14421 : tmp14440;
  assign tmp14521 = s2 ? 1 : tmp14522;
  assign tmp14520 = s3 ? tmp14521 : 1;
  assign tmp14516 = s4 ? tmp14517 : tmp14520;
  assign tmp14515 = s5 ? tmp14458 : tmp14516;
  assign tmp14514 = s6 ? tmp14418 : tmp14515;
  assign tmp14513 = s7 ? tmp14417 : tmp14514;
  assign tmp14512 = s8 ? tmp14513 : tmp14417;
  assign tmp14529 = s2 ? 1 : tmp14421;
  assign tmp14528 = s3 ? tmp14529 : 1;
  assign tmp14527 = s4 ? tmp14466 : tmp14528;
  assign tmp14526 = s5 ? tmp14458 : tmp14527;
  assign tmp14525 = s6 ? tmp14418 : tmp14526;
  assign tmp14531 = s5 ? tmp14504 : 1;
  assign tmp14530 = s6 ? 1 : tmp14531;
  assign tmp14524 = s7 ? tmp14525 : tmp14530;
  assign tmp14535 = s4 ? tmp14479 : 1;
  assign tmp14534 = s5 ? 1 : tmp14535;
  assign tmp14533 = s6 ? 1 : tmp14534;
  assign tmp14538 = s4 ? tmp14517 : tmp14528;
  assign tmp14537 = s5 ? tmp14458 : tmp14538;
  assign tmp14536 = s6 ? tmp14418 : tmp14537;
  assign tmp14532 = s7 ? tmp14533 : tmp14536;
  assign tmp14523 = s8 ? tmp14524 : tmp14532;
  assign tmp14511 = s9 ? tmp14512 : tmp14523;
  assign tmp14413 = s10 ? tmp14414 : tmp14511;
  assign tmp14542 = s7 ? tmp14456 : tmp14502;
  assign tmp14543 = s7 ? tmp14476 : tmp14514;
  assign tmp14541 = s8 ? tmp14542 : tmp14543;
  assign tmp14540 = s9 ? tmp14512 : tmp14541;
  assign tmp14539 = s10 ? tmp14414 : tmp14540;
  assign tmp14412 = s11 ? tmp14413 : tmp14539;
  assign tmp14553 = s2 ? 1 : tmp14440;
  assign tmp14552 = s3 ? tmp14553 : 1;
  assign tmp14551 = s4 ? tmp14479 : tmp14552;
  assign tmp14550 = s5 ? 1 : tmp14551;
  assign tmp14549 = s6 ? 1 : tmp14550;
  assign tmp14548 = s7 ? 1 : tmp14549;
  assign tmp14547 = s8 ? tmp14548 : tmp14475;
  assign tmp14554 = s8 ? tmp14475 : 1;
  assign tmp14546 = s9 ? tmp14547 : tmp14554;
  assign tmp14556 = s8 ? tmp14548 : 1;
  assign tmp14558 = s7 ? tmp14533 : 1;
  assign tmp14557 = s8 ? tmp14558 : tmp14533;
  assign tmp14555 = s9 ? tmp14556 : tmp14557;
  assign tmp14545 = s10 ? tmp14546 : tmp14555;
  assign tmp14562 = s7 ? tmp14549 : 1;
  assign tmp14563 = s7 ? tmp14476 : tmp14549;
  assign tmp14561 = s8 ? tmp14562 : tmp14563;
  assign tmp14560 = s9 ? tmp14556 : tmp14561;
  assign tmp14559 = s10 ? tmp14546 : tmp14560;
  assign tmp14544 = s11 ? tmp14545 : tmp14559;
  assign tmp14411 = s12 ? tmp14412 : tmp14544;
  assign tmp14410 = s13 ? 1 : tmp14411;
  assign tmp14409 = s14 ? 1 : tmp14410;
  assign tmp14578 = ~(l4 ? 1 : 0);
  assign tmp14577 = l2 ? 1 : tmp14578;
  assign tmp14576 = l1 ? 1 : tmp14577;
  assign tmp14575 = s0 ? 1 : tmp14576;
  assign tmp14580 = s1 ? tmp14425 : tmp14576;
  assign tmp14579 = s2 ? tmp14576 : tmp14580;
  assign tmp14574 = s3 ? tmp14575 : tmp14579;
  assign tmp14584 = s0 ? tmp14576 : 1;
  assign tmp14583 = s1 ? tmp14584 : tmp14576;
  assign tmp14585 = s1 ? tmp14584 : 1;
  assign tmp14582 = s2 ? tmp14583 : tmp14585;
  assign tmp14587 = s1 ? tmp14576 : tmp14575;
  assign tmp14586 = s2 ? 1 : tmp14587;
  assign tmp14581 = s3 ? tmp14582 : tmp14586;
  assign tmp14573 = s4 ? tmp14574 : tmp14581;
  assign tmp14593 = s0 ? tmp14576 : tmp14440;
  assign tmp14592 = s1 ? tmp14575 : tmp14593;
  assign tmp14591 = s2 ? tmp14585 : tmp14592;
  assign tmp14595 = s0 ? tmp14440 : tmp14576;
  assign tmp14596 = s1 ? 1 : tmp14576;
  assign tmp14594 = s2 ? tmp14595 : tmp14596;
  assign tmp14590 = s3 ? tmp14591 : tmp14594;
  assign tmp14599 = s1 ? tmp14575 : 1;
  assign tmp14600 = s1 ? 1 : tmp14584;
  assign tmp14598 = s2 ? tmp14599 : tmp14600;
  assign tmp14601 = s2 ? tmp14587 : 1;
  assign tmp14597 = s3 ? tmp14598 : tmp14601;
  assign tmp14589 = s4 ? tmp14590 : tmp14597;
  assign tmp14604 = s2 ? tmp14585 : 1;
  assign tmp14606 = s1 ? 1 : tmp14575;
  assign tmp14605 = s2 ? 1 : tmp14606;
  assign tmp14603 = s3 ? tmp14604 : tmp14605;
  assign tmp14608 = s2 ? tmp14585 : tmp14599;
  assign tmp14609 = s2 ? tmp14606 : tmp14599;
  assign tmp14607 = s3 ? tmp14608 : tmp14609;
  assign tmp14602 = s4 ? tmp14603 : tmp14607;
  assign tmp14588 = s5 ? tmp14589 : tmp14602;
  assign tmp14572 = s6 ? tmp14573 : tmp14588;
  assign tmp14615 = s1 ? tmp14576 : tmp14593;
  assign tmp14614 = s2 ? tmp14585 : tmp14615;
  assign tmp14616 = s2 ? tmp14576 : tmp14596;
  assign tmp14613 = s3 ? tmp14614 : tmp14616;
  assign tmp14618 = s2 ? tmp14599 : tmp14596;
  assign tmp14617 = s3 ? tmp14618 : tmp14601;
  assign tmp14612 = s4 ? tmp14613 : tmp14617;
  assign tmp14621 = s2 ? tmp14470 : tmp14596;
  assign tmp14620 = s3 ? tmp14604 : tmp14621;
  assign tmp14623 = s2 ? tmp14585 : tmp14576;
  assign tmp14624 = s2 ? tmp14596 : tmp14576;
  assign tmp14622 = s3 ? tmp14623 : tmp14624;
  assign tmp14619 = s4 ? tmp14620 : tmp14622;
  assign tmp14611 = s5 ? tmp14612 : tmp14619;
  assign tmp14610 = s6 ? tmp14573 : tmp14611;
  assign tmp14571 = s7 ? tmp14572 : tmp14610;
  assign tmp14628 = s3 ? tmp14575 : tmp14616;
  assign tmp14627 = s4 ? tmp14628 : tmp14581;
  assign tmp14633 = s1 ? tmp14575 : tmp14584;
  assign tmp14632 = s2 ? tmp14585 : tmp14633;
  assign tmp14634 = s2 ? tmp14575 : tmp14596;
  assign tmp14631 = s3 ? tmp14632 : tmp14634;
  assign tmp14630 = s4 ? tmp14631 : tmp14597;
  assign tmp14629 = s5 ? tmp14630 : tmp14602;
  assign tmp14626 = s6 ? tmp14627 : tmp14629;
  assign tmp14640 = s1 ? tmp14576 : tmp14584;
  assign tmp14639 = s2 ? tmp14585 : tmp14640;
  assign tmp14638 = s3 ? tmp14639 : tmp14616;
  assign tmp14642 = s2 ? tmp14599 : tmp14576;
  assign tmp14643 = s2 ? tmp14576 : 1;
  assign tmp14641 = s3 ? tmp14642 : tmp14643;
  assign tmp14637 = s4 ? tmp14638 : tmp14641;
  assign tmp14636 = s5 ? tmp14637 : tmp14619;
  assign tmp14635 = s6 ? tmp14627 : tmp14636;
  assign tmp14625 = s7 ? tmp14626 : tmp14635;
  assign tmp14570 = s8 ? tmp14571 : tmp14625;
  assign tmp14650 = s2 ? tmp14425 : 1;
  assign tmp14649 = s3 ? tmp14489 : tmp14650;
  assign tmp14648 = s4 ? tmp14649 : 1;
  assign tmp14647 = s5 ? tmp14648 : 1;
  assign tmp14646 = s6 ? 1 : tmp14647;
  assign tmp14653 = s4 ? tmp14501 : 1;
  assign tmp14652 = s5 ? tmp14653 : 1;
  assign tmp14651 = s6 ? 1 : tmp14652;
  assign tmp14645 = s7 ? tmp14646 : tmp14651;
  assign tmp14644 = s8 ? tmp14625 : tmp14645;
  assign tmp14569 = s9 ? tmp14570 : tmp14644;
  assign tmp14663 = s0 ? tmp14576 : tmp14421;
  assign tmp14662 = s1 ? tmp14575 : tmp14663;
  assign tmp14661 = s2 ? tmp14585 : tmp14662;
  assign tmp14665 = s0 ? tmp14421 : tmp14576;
  assign tmp14664 = s2 ? tmp14665 : tmp14596;
  assign tmp14660 = s3 ? tmp14661 : tmp14664;
  assign tmp14659 = s4 ? tmp14660 : tmp14597;
  assign tmp14658 = s5 ? tmp14659 : tmp14602;
  assign tmp14657 = s6 ? tmp14573 : tmp14658;
  assign tmp14671 = s1 ? tmp14576 : tmp14663;
  assign tmp14670 = s2 ? tmp14585 : tmp14671;
  assign tmp14669 = s3 ? tmp14670 : tmp14616;
  assign tmp14668 = s4 ? tmp14669 : tmp14641;
  assign tmp14667 = s5 ? tmp14668 : tmp14619;
  assign tmp14666 = s6 ? tmp14573 : tmp14667;
  assign tmp14656 = s7 ? tmp14657 : tmp14666;
  assign tmp14655 = s8 ? tmp14656 : tmp14657;
  assign tmp14677 = s3 ? tmp14618 : tmp14643;
  assign tmp14676 = s4 ? tmp14613 : tmp14677;
  assign tmp14679 = s3 ? tmp14623 : tmp14596;
  assign tmp14678 = s4 ? tmp14620 : tmp14679;
  assign tmp14675 = s5 ? tmp14676 : tmp14678;
  assign tmp14674 = s6 ? tmp14573 : tmp14675;
  assign tmp14673 = s7 ? tmp14674 : tmp14651;
  assign tmp14682 = s5 ? tmp14637 : tmp14678;
  assign tmp14681 = s6 ? tmp14627 : tmp14682;
  assign tmp14684 = s5 ? tmp14668 : tmp14678;
  assign tmp14683 = s6 ? tmp14573 : tmp14684;
  assign tmp14680 = s7 ? tmp14681 : tmp14683;
  assign tmp14672 = s8 ? tmp14673 : tmp14680;
  assign tmp14654 = s9 ? tmp14655 : tmp14672;
  assign tmp14568 = s10 ? tmp14569 : tmp14654;
  assign tmp14688 = s7 ? tmp14610 : tmp14651;
  assign tmp14689 = s7 ? tmp14635 : tmp14666;
  assign tmp14687 = s8 ? tmp14688 : tmp14689;
  assign tmp14686 = s9 ? tmp14655 : tmp14687;
  assign tmp14685 = s10 ? tmp14569 : tmp14686;
  assign tmp14567 = s11 ? tmp14568 : tmp14685;
  assign tmp14566 = s12 ? tmp14567 : 1;
  assign tmp14565 = s13 ? tmp14566 : 1;
  assign tmp14564 = s14 ? 1 : tmp14565;
  assign tmp14408 = s15 ? tmp14409 : tmp14564;
  assign tmp14407 = s16 ? tmp14408 : 1;
  assign tmp14706 = ~(l2 ? 1 : 0);
  assign tmp14705 = s0 ? 1 : tmp14706;
  assign tmp14704 = s1 ? tmp14705 : 1;
  assign tmp14703 = s2 ? tmp14704 : 1;
  assign tmp14702 = s3 ? tmp14703 : 1;
  assign tmp14710 = s0 ? tmp14422 : 0;
  assign tmp14709 = ~(s1 ? tmp14710 : 0);
  assign tmp14708 = s2 ? 1 : tmp14709;
  assign tmp14707 = s3 ? tmp14708 : 1;
  assign tmp14701 = s4 ? tmp14702 : tmp14707;
  assign tmp14700 = s5 ? 1 : tmp14701;
  assign tmp14699 = s6 ? 1 : tmp14700;
  assign tmp14713 = s4 ? tmp14702 : 1;
  assign tmp14712 = s5 ? 1 : tmp14713;
  assign tmp14711 = s6 ? 1 : tmp14712;
  assign tmp14698 = s7 ? tmp14699 : tmp14711;
  assign tmp14722 = ~(l1 ? 1 : 0);
  assign tmp14721 = s0 ? 1 : tmp14722;
  assign tmp14720 = s1 ? 1 : tmp14721;
  assign tmp14719 = s2 ? 1 : tmp14720;
  assign tmp14724 = s0 ? tmp14440 : 0;
  assign tmp14723 = ~(s2 ? tmp14724 : 0);
  assign tmp14718 = s3 ? tmp14719 : tmp14723;
  assign tmp14717 = s4 ? tmp14718 : 1;
  assign tmp14716 = s5 ? tmp14717 : tmp14701;
  assign tmp14715 = s6 ? 1 : tmp14716;
  assign tmp14728 = s3 ? tmp14719 : 1;
  assign tmp14732 = l1 ? tmp14422 : 0;
  assign tmp14734 = ~(l1 ? tmp14422 : 0);
  assign tmp14733 = ~(s0 ? 1 : tmp14734);
  assign tmp14731 = ~(s1 ? tmp14732 : tmp14733);
  assign tmp14730 = s2 ? 1 : tmp14731;
  assign tmp14729 = s3 ? tmp14730 : 1;
  assign tmp14727 = s4 ? tmp14728 : tmp14729;
  assign tmp14726 = s5 ? tmp14727 : tmp14713;
  assign tmp14725 = s6 ? 1 : tmp14726;
  assign tmp14714 = s7 ? tmp14715 : tmp14725;
  assign tmp14697 = s8 ? tmp14698 : tmp14714;
  assign tmp14741 = s2 ? tmp14494 : 1;
  assign tmp14740 = s3 ? tmp14741 : 1;
  assign tmp14743 = s2 ? 1 : tmp14470;
  assign tmp14742 = s3 ? tmp14743 : 1;
  assign tmp14739 = s4 ? tmp14740 : tmp14742;
  assign tmp14738 = s5 ? 1 : tmp14739;
  assign tmp14737 = s6 ? 1 : tmp14738;
  assign tmp14746 = s4 ? tmp14740 : 1;
  assign tmp14745 = s5 ? 1 : tmp14746;
  assign tmp14744 = s6 ? 1 : tmp14745;
  assign tmp14736 = s7 ? tmp14737 : tmp14744;
  assign tmp14735 = s8 ? tmp14714 : tmp14736;
  assign tmp14696 = s9 ? tmp14697 : tmp14735;
  assign tmp14748 = s8 ? tmp14698 : tmp14699;
  assign tmp14750 = s7 ? tmp14711 : tmp14744;
  assign tmp14757 = ~(s1 ? tmp14732 : 0);
  assign tmp14756 = s2 ? 1 : tmp14757;
  assign tmp14755 = s3 ? tmp14756 : 1;
  assign tmp14754 = s4 ? tmp14728 : tmp14755;
  assign tmp14753 = s5 ? tmp14754 : tmp14713;
  assign tmp14752 = s6 ? 1 : tmp14753;
  assign tmp14751 = s7 ? tmp14752 : tmp14711;
  assign tmp14749 = s8 ? tmp14750 : tmp14751;
  assign tmp14747 = s9 ? tmp14748 : tmp14749;
  assign tmp14695 = s10 ? tmp14696 : tmp14747;
  assign tmp14761 = s7 ? tmp14725 : tmp14711;
  assign tmp14760 = s8 ? tmp14750 : tmp14761;
  assign tmp14759 = s9 ? tmp14748 : tmp14760;
  assign tmp14758 = s10 ? tmp14696 : tmp14759;
  assign tmp14694 = s11 ? tmp14695 : tmp14758;
  assign tmp14773 = s0 ? 1 : 0;
  assign tmp14772 = s1 ? 1 : tmp14773;
  assign tmp14775 = ~(s0 ? 1 : 0);
  assign tmp14774 = s1 ? 1 : tmp14775;
  assign tmp14771 = s2 ? tmp14772 : tmp14774;
  assign tmp14770 = s3 ? 1 : tmp14771;
  assign tmp14769 = s4 ? 1 : tmp14770;
  assign tmp14780 = ~(s1 ? 1 : tmp14775);
  assign tmp14779 = s2 ? tmp14772 : tmp14780;
  assign tmp14778 = s3 ? 1 : tmp14779;
  assign tmp14783 = s1 ? tmp14773 : tmp14775;
  assign tmp14784 = ~(s1 ? tmp14773 : 1);
  assign tmp14782 = s2 ? tmp14783 : tmp14784;
  assign tmp14781 = ~(s3 ? tmp14782 : 1);
  assign tmp14777 = s4 ? tmp14778 : tmp14781;
  assign tmp14776 = s5 ? tmp14777 : 0;
  assign tmp14768 = s6 ? tmp14769 : tmp14776;
  assign tmp14790 = s1 ? 1 : 0;
  assign tmp14789 = s2 ? tmp14790 : tmp14780;
  assign tmp14788 = s3 ? 1 : tmp14789;
  assign tmp14792 = s2 ? tmp14783 : 0;
  assign tmp14791 = ~(s3 ? tmp14792 : 1);
  assign tmp14787 = s4 ? tmp14788 : tmp14791;
  assign tmp14786 = s5 ? tmp14787 : 0;
  assign tmp14785 = s6 ? tmp14769 : tmp14786;
  assign tmp14767 = s7 ? tmp14768 : tmp14785;
  assign tmp14799 = ~(s1 ? 1 : 0);
  assign tmp14798 = s2 ? tmp14772 : tmp14799;
  assign tmp14797 = s3 ? 1 : tmp14798;
  assign tmp14802 = s1 ? tmp14773 : 0;
  assign tmp14801 = s2 ? tmp14802 : 0;
  assign tmp14800 = ~(s3 ? tmp14801 : 1);
  assign tmp14796 = s4 ? tmp14797 : tmp14800;
  assign tmp14795 = s5 ? tmp14796 : 0;
  assign tmp14794 = s6 ? tmp14769 : tmp14795;
  assign tmp14808 = s0 ? 1 : tmp14734;
  assign tmp14807 = s1 ? 1 : tmp14808;
  assign tmp14806 = s2 ? 1 : tmp14807;
  assign tmp14811 = ~(s0 ? tmp14732 : 1);
  assign tmp14810 = s1 ? 1 : tmp14811;
  assign tmp14809 = s2 ? tmp14810 : tmp14774;
  assign tmp14805 = s3 ? tmp14806 : tmp14809;
  assign tmp14804 = s4 ? 1 : tmp14805;
  assign tmp14815 = s2 ? tmp14790 : tmp14799;
  assign tmp14814 = s3 ? 1 : tmp14815;
  assign tmp14813 = s4 ? tmp14814 : tmp14800;
  assign tmp14812 = s5 ? tmp14813 : 0;
  assign tmp14803 = s6 ? tmp14804 : tmp14812;
  assign tmp14793 = s7 ? tmp14794 : tmp14803;
  assign tmp14766 = s8 ? tmp14767 : tmp14793;
  assign tmp14821 = s2 ? tmp14790 : tmp14774;
  assign tmp14820 = s3 ? 1 : tmp14821;
  assign tmp14819 = s4 ? 1 : tmp14820;
  assign tmp14818 = s6 ? tmp14819 : tmp14786;
  assign tmp14817 = s7 ? tmp14768 : tmp14818;
  assign tmp14816 = s8 ? tmp14793 : tmp14817;
  assign tmp14765 = s9 ? tmp14766 : tmp14816;
  assign tmp14823 = s8 ? tmp14817 : tmp14768;
  assign tmp14828 = s3 ? tmp14806 : tmp14821;
  assign tmp14827 = s4 ? 1 : tmp14828;
  assign tmp14826 = s6 ? tmp14827 : tmp14812;
  assign tmp14825 = s7 ? tmp14826 : tmp14818;
  assign tmp14824 = s8 ? tmp14818 : tmp14825;
  assign tmp14822 = s9 ? tmp14823 : tmp14824;
  assign tmp14764 = s10 ? tmp14765 : tmp14822;
  assign tmp14832 = s7 ? tmp14803 : tmp14818;
  assign tmp14831 = s8 ? tmp14785 : tmp14832;
  assign tmp14830 = s9 ? tmp14823 : tmp14831;
  assign tmp14829 = s10 ? tmp14765 : tmp14830;
  assign tmp14763 = s11 ? tmp14764 : tmp14829;
  assign tmp14762 = s12 ? 1 : tmp14763;
  assign tmp14693 = s13 ? tmp14694 : tmp14762;
  assign tmp14846 = ~(s0 ? 1 : tmp14722);
  assign tmp14845 = s1 ? tmp14724 : tmp14846;
  assign tmp14847 = ~(s1 ? tmp14721 : tmp14722);
  assign tmp14844 = s2 ? tmp14845 : tmp14847;
  assign tmp14849 = s1 ? tmp14440 : tmp14724;
  assign tmp14848 = s2 ? tmp14849 : tmp14471;
  assign tmp14843 = s3 ? tmp14844 : tmp14848;
  assign tmp14852 = s1 ? tmp14440 : tmp14471;
  assign tmp14853 = s1 ? tmp14471 : tmp14440;
  assign tmp14851 = s2 ? tmp14852 : tmp14853;
  assign tmp14854 = ~(s1 ? tmp14773 : 0);
  assign tmp14850 = s3 ? tmp14851 : tmp14854;
  assign tmp14842 = s4 ? tmp14843 : tmp14850;
  assign tmp14841 = s5 ? tmp14842 : 0;
  assign tmp14840 = s6 ? tmp14440 : tmp14841;
  assign tmp14860 = s1 ? tmp14724 : tmp14440;
  assign tmp14859 = s2 ? tmp14860 : tmp14440;
  assign tmp14865 = l3 ? 1 : 0;
  assign tmp14864 = ~(l2 ? tmp14865 : 1);
  assign tmp14863 = l1 ? 1 : tmp14864;
  assign tmp14866 = s0 ? tmp14863 : 0;
  assign tmp14862 = s1 ? tmp14863 : tmp14866;
  assign tmp14861 = s2 ? tmp14862 : tmp14471;
  assign tmp14858 = s3 ? tmp14859 : tmp14861;
  assign tmp14868 = s2 ? tmp14852 : tmp14440;
  assign tmp14869 = ~(s2 ? tmp14773 : 1);
  assign tmp14867 = s3 ? tmp14868 : tmp14869;
  assign tmp14857 = s4 ? tmp14858 : tmp14867;
  assign tmp14856 = s5 ? tmp14857 : 0;
  assign tmp14855 = s6 ? tmp14440 : tmp14856;
  assign tmp14839 = ~(s7 ? tmp14840 : tmp14855);
  assign tmp14838 = s8 ? 1 : tmp14839;
  assign tmp14871 = s7 ? tmp14840 : tmp14855;
  assign tmp14870 = ~(s8 ? tmp14871 : 0);
  assign tmp14837 = s9 ? tmp14838 : tmp14870;
  assign tmp14880 = s1 ? tmp14863 : 0;
  assign tmp14879 = s2 ? tmp14880 : tmp14471;
  assign tmp14878 = s3 ? tmp14859 : tmp14879;
  assign tmp14877 = s4 ? tmp14878 : tmp14867;
  assign tmp14876 = s5 ? tmp14877 : 0;
  assign tmp14875 = s6 ? tmp14440 : tmp14876;
  assign tmp14874 = ~(s7 ? tmp14875 : 0);
  assign tmp14873 = s8 ? 1 : tmp14874;
  assign tmp14872 = s9 ? 1 : tmp14873;
  assign tmp14836 = s10 ? tmp14837 : tmp14872;
  assign tmp14884 = ~(s7 ? tmp14855 : 0);
  assign tmp14883 = s8 ? 1 : tmp14884;
  assign tmp14882 = s9 ? 1 : tmp14883;
  assign tmp14881 = s10 ? tmp14837 : tmp14882;
  assign tmp14835 = s11 ? tmp14836 : tmp14881;
  assign tmp14894 = s1 ? tmp14773 : 1;
  assign tmp14893 = s2 ? 1 : tmp14894;
  assign tmp14892 = s3 ? 1 : tmp14893;
  assign tmp14896 = s2 ? 1 : tmp14773;
  assign tmp14897 = s2 ? tmp14774 : 1;
  assign tmp14895 = s3 ? tmp14896 : tmp14897;
  assign tmp14891 = s4 ? tmp14892 : tmp14895;
  assign tmp14902 = ~(s1 ? tmp14773 : tmp14775);
  assign tmp14901 = s2 ? tmp14783 : tmp14902;
  assign tmp14903 = ~(s2 ? tmp14773 : 0);
  assign tmp14900 = s3 ? tmp14901 : tmp14903;
  assign tmp14899 = s4 ? tmp14900 : 1;
  assign tmp14898 = s5 ? tmp14899 : 1;
  assign tmp14890 = s6 ? tmp14891 : tmp14898;
  assign tmp14906 = s3 ? tmp14893 : 1;
  assign tmp14905 = s4 ? tmp14892 : tmp14906;
  assign tmp14910 = s2 ? tmp14894 : tmp14772;
  assign tmp14909 = s3 ? tmp14910 : 1;
  assign tmp14908 = s4 ? tmp14909 : 1;
  assign tmp14907 = s5 ? tmp14908 : 1;
  assign tmp14904 = s6 ? tmp14905 : tmp14907;
  assign tmp14889 = s7 ? tmp14890 : tmp14904;
  assign tmp14918 = l4 ? 1 : 0;
  assign tmp14917 = l2 ? tmp14918 : 0;
  assign tmp14916 = l1 ? tmp14422 : tmp14917;
  assign tmp14920 = l1 ? tmp14422 : tmp14918;
  assign tmp14919 = s0 ? tmp14920 : tmp14916;
  assign tmp14915 = s1 ? tmp14916 : tmp14919;
  assign tmp14923 = s0 ? tmp14916 : 1;
  assign tmp14922 = s1 ? tmp14923 : tmp14916;
  assign tmp14921 = s2 ? tmp14916 : tmp14922;
  assign tmp14914 = s3 ? tmp14915 : tmp14921;
  assign tmp14927 = s0 ? tmp14916 : tmp14422;
  assign tmp14926 = s1 ? tmp14927 : tmp14916;
  assign tmp14929 = s0 ? tmp14920 : 1;
  assign tmp14928 = s1 ? tmp14923 : tmp14929;
  assign tmp14925 = s2 ? tmp14926 : tmp14928;
  assign tmp14931 = s1 ? tmp14920 : tmp14773;
  assign tmp14933 = s0 ? tmp14918 : tmp14916;
  assign tmp14932 = s1 ? tmp14916 : tmp14933;
  assign tmp14930 = s2 ? tmp14931 : tmp14932;
  assign tmp14924 = s3 ? tmp14925 : tmp14930;
  assign tmp14913 = s4 ? tmp14914 : tmp14924;
  assign tmp14939 = s0 ? 1 : tmp14422;
  assign tmp14938 = s1 ? tmp14923 : tmp14939;
  assign tmp14941 = s0 ? 1 : tmp14916;
  assign tmp14940 = s1 ? tmp14941 : tmp14923;
  assign tmp14937 = s2 ? tmp14938 : tmp14940;
  assign tmp14944 = s0 ? tmp14918 : 0;
  assign tmp14943 = s1 ? tmp14944 : tmp14916;
  assign tmp14942 = s2 ? tmp14941 : tmp14943;
  assign tmp14936 = s3 ? tmp14937 : tmp14942;
  assign tmp14949 = ~(l1 ? tmp14422 : tmp14917);
  assign tmp14948 = s0 ? 1 : tmp14949;
  assign tmp14951 = l1 ? tmp14422 : 1;
  assign tmp14950 = ~(s0 ? tmp14951 : tmp14920);
  assign tmp14947 = s1 ? tmp14948 : tmp14950;
  assign tmp14953 = s0 ? tmp14951 : tmp14920;
  assign tmp14952 = ~(s1 ? tmp14953 : tmp14927);
  assign tmp14946 = s2 ? tmp14947 : tmp14952;
  assign tmp14956 = s0 ? tmp14920 : 0;
  assign tmp14955 = s1 ? tmp14916 : tmp14956;
  assign tmp14954 = ~(s2 ? tmp14955 : 0);
  assign tmp14945 = ~(s3 ? tmp14946 : tmp14954);
  assign tmp14935 = s4 ? tmp14936 : tmp14945;
  assign tmp14961 = s0 ? tmp14916 : 0;
  assign tmp14962 = ~(s0 ? 1 : tmp14578);
  assign tmp14960 = s1 ? tmp14961 : tmp14962;
  assign tmp14964 = s0 ? tmp14918 : tmp14422;
  assign tmp14963 = s1 ? tmp14964 : tmp14422;
  assign tmp14959 = s2 ? tmp14960 : tmp14963;
  assign tmp14958 = s3 ? tmp14959 : 0;
  assign tmp14968 = s0 ? 1 : tmp14578;
  assign tmp14967 = s1 ? 1 : tmp14968;
  assign tmp14969 = s1 ? tmp14948 : tmp14706;
  assign tmp14966 = s2 ? tmp14967 : tmp14969;
  assign tmp14971 = s1 ? tmp14944 : 0;
  assign tmp14970 = ~(s2 ? tmp14971 : 0);
  assign tmp14965 = ~(s3 ? tmp14966 : tmp14970);
  assign tmp14957 = s4 ? tmp14958 : tmp14965;
  assign tmp14934 = s5 ? tmp14935 : tmp14957;
  assign tmp14912 = s6 ? tmp14913 : tmp14934;
  assign tmp14976 = s1 ? tmp14923 : tmp14920;
  assign tmp14975 = s2 ? tmp14926 : tmp14976;
  assign tmp14978 = s1 ? tmp14920 : 0;
  assign tmp14977 = s2 ? tmp14978 : tmp14932;
  assign tmp14974 = s3 ? tmp14975 : tmp14977;
  assign tmp14973 = s4 ? tmp14914 : tmp14974;
  assign tmp14983 = s1 ? tmp14923 : tmp14422;
  assign tmp14984 = s1 ? tmp14916 : tmp14923;
  assign tmp14982 = s2 ? tmp14983 : tmp14984;
  assign tmp14985 = s2 ? tmp14916 : tmp14943;
  assign tmp14981 = s3 ? tmp14982 : tmp14985;
  assign tmp14988 = ~(s1 ? tmp14920 : tmp14916);
  assign tmp14987 = s2 ? tmp14947 : tmp14988;
  assign tmp14986 = ~(s3 ? tmp14987 : tmp14954);
  assign tmp14980 = s4 ? tmp14981 : tmp14986;
  assign tmp14992 = s1 ? tmp14961 : tmp14918;
  assign tmp14993 = s1 ? tmp14422 : 0;
  assign tmp14991 = s2 ? tmp14992 : tmp14993;
  assign tmp14990 = s3 ? tmp14991 : 0;
  assign tmp14996 = s1 ? 1 : tmp14578;
  assign tmp14995 = s2 ? tmp14996 : tmp14949;
  assign tmp14994 = ~(s3 ? tmp14995 : 1);
  assign tmp14989 = s4 ? tmp14990 : tmp14994;
  assign tmp14979 = s5 ? tmp14980 : tmp14989;
  assign tmp14972 = s6 ? tmp14973 : tmp14979;
  assign tmp14911 = ~(s7 ? tmp14912 : tmp14972);
  assign tmp14888 = s8 ? tmp14889 : tmp14911;
  assign tmp14998 = s7 ? tmp14912 : tmp14972;
  assign tmp14999 = ~(s7 ? tmp14890 : tmp14904);
  assign tmp14997 = ~(s8 ? tmp14998 : tmp14999);
  assign tmp14887 = s9 ? tmp14888 : tmp14997;
  assign tmp15001 = s8 ? tmp14889 : tmp14890;
  assign tmp15009 = s1 ? tmp14916 : 0;
  assign tmp15008 = ~(s2 ? tmp15009 : 0);
  assign tmp15007 = ~(s3 ? tmp14987 : tmp15008);
  assign tmp15006 = s4 ? tmp14981 : tmp15007;
  assign tmp15005 = s5 ? tmp15006 : tmp14989;
  assign tmp15004 = s6 ? tmp14973 : tmp15005;
  assign tmp15010 = ~(s6 ? tmp14905 : tmp14907);
  assign tmp15003 = ~(s7 ? tmp15004 : tmp15010);
  assign tmp15002 = s8 ? tmp14904 : tmp15003;
  assign tmp15000 = s9 ? tmp15001 : tmp15002;
  assign tmp14886 = s10 ? tmp14887 : tmp15000;
  assign tmp15014 = ~(s7 ? tmp14972 : tmp15010);
  assign tmp15013 = s8 ? tmp14904 : tmp15014;
  assign tmp15012 = s9 ? tmp15001 : tmp15013;
  assign tmp15011 = s10 ? tmp14887 : tmp15012;
  assign tmp14885 = s11 ? tmp14886 : tmp15011;
  assign tmp14834 = s12 ? tmp14835 : tmp14885;
  assign tmp15024 = l2 ? tmp14865 : 0;
  assign tmp15023 = l1 ? 1 : tmp15024;
  assign tmp15029 = ~(l2 ? tmp14865 : 0);
  assign tmp15028 = ~(l1 ? 1 : tmp15029);
  assign tmp15027 = s0 ? tmp15023 : tmp15028;
  assign tmp15026 = s1 ? tmp15027 : tmp15023;
  assign tmp15025 = s2 ? tmp15023 : tmp15026;
  assign tmp15022 = s3 ? tmp15023 : tmp15025;
  assign tmp15032 = s0 ? tmp15023 : 1;
  assign tmp15031 = s2 ? tmp15023 : tmp15032;
  assign tmp15035 = l1 ? 1 : tmp14865;
  assign tmp15034 = s1 ? tmp15035 : 1;
  assign tmp15037 = s0 ? 1 : tmp15023;
  assign tmp15036 = s1 ? tmp15023 : tmp15037;
  assign tmp15033 = s2 ? tmp15034 : tmp15036;
  assign tmp15030 = s3 ? tmp15031 : tmp15033;
  assign tmp15021 = s4 ? tmp15022 : tmp15030;
  assign tmp15044 = l1 ? 1 : tmp15029;
  assign tmp15045 = ~(l1 ? 1 : tmp15024);
  assign tmp15043 = ~(s0 ? tmp15044 : tmp15045);
  assign tmp15042 = s1 ? tmp15027 : tmp15043;
  assign tmp15047 = s0 ? tmp15044 : tmp15045;
  assign tmp15048 = ~(s0 ? tmp15023 : tmp15028);
  assign tmp15046 = ~(s1 ? tmp15047 : tmp15048);
  assign tmp15041 = s2 ? tmp15042 : tmp15046;
  assign tmp15051 = s0 ? tmp15023 : tmp14440;
  assign tmp15050 = ~(s1 ? 1 : tmp15051);
  assign tmp15049 = ~(s2 ? tmp15047 : tmp15050);
  assign tmp15040 = s3 ? tmp15041 : tmp15049;
  assign tmp15055 = s0 ? tmp14440 : tmp15023;
  assign tmp15054 = s1 ? tmp15055 : tmp14444;
  assign tmp15056 = s1 ? tmp14444 : tmp15023;
  assign tmp15053 = s2 ? tmp15054 : tmp15056;
  assign tmp15058 = s1 ? tmp15051 : 1;
  assign tmp15057 = s2 ? tmp15058 : 1;
  assign tmp15052 = s3 ? tmp15053 : tmp15057;
  assign tmp15039 = s4 ? tmp15040 : tmp15052;
  assign tmp15062 = s1 ? tmp15037 : tmp15055;
  assign tmp15061 = s2 ? tmp15058 : tmp15062;
  assign tmp15060 = s3 ? tmp15061 : 1;
  assign tmp15065 = s1 ? tmp15055 : tmp15051;
  assign tmp15064 = s2 ? 1 : tmp15065;
  assign tmp15063 = s3 ? tmp15064 : 1;
  assign tmp15059 = s4 ? tmp15060 : tmp15063;
  assign tmp15038 = s5 ? tmp15039 : tmp15059;
  assign tmp15020 = s6 ? tmp15021 : tmp15038;
  assign tmp15070 = s1 ? tmp15032 : tmp15035;
  assign tmp15069 = s2 ? tmp15023 : tmp15070;
  assign tmp15068 = s3 ? tmp15069 : tmp15033;
  assign tmp15067 = s4 ? tmp15022 : tmp15068;
  assign tmp15075 = s1 ? tmp15023 : tmp15027;
  assign tmp15074 = s2 ? tmp15026 : tmp15075;
  assign tmp15077 = s1 ? 1 : tmp15051;
  assign tmp15076 = s2 ? tmp15023 : tmp15077;
  assign tmp15073 = s3 ? tmp15074 : tmp15076;
  assign tmp15079 = s2 ? tmp15054 : tmp15023;
  assign tmp15078 = s3 ? tmp15079 : tmp15057;
  assign tmp15072 = s4 ? tmp15073 : tmp15078;
  assign tmp15083 = s1 ? tmp15023 : tmp15055;
  assign tmp15082 = s2 ? tmp15058 : tmp15083;
  assign tmp15081 = s3 ? tmp15082 : tmp14469;
  assign tmp15086 = s1 ? tmp15023 : tmp15051;
  assign tmp15085 = s2 ? 1 : tmp15086;
  assign tmp15084 = s3 ? tmp15085 : 1;
  assign tmp15080 = s4 ? tmp15081 : tmp15084;
  assign tmp15071 = s5 ? tmp15072 : tmp15080;
  assign tmp15066 = s6 ? tmp15067 : tmp15071;
  assign tmp15019 = s7 ? tmp15020 : tmp15066;
  assign tmp15093 = s1 ? tmp14721 : 1;
  assign tmp15092 = s2 ? 1 : tmp15093;
  assign tmp15091 = s3 ? 1 : tmp15092;
  assign tmp15090 = s4 ? tmp15091 : 1;
  assign tmp15099 = ~(s0 ? tmp14440 : 0);
  assign tmp15098 = s1 ? tmp14721 : tmp15099;
  assign tmp15100 = ~(s1 ? tmp14724 : tmp14846);
  assign tmp15097 = s2 ? tmp15098 : tmp15100;
  assign tmp15102 = ~(s1 ? 1 : tmp14444);
  assign tmp15101 = ~(s2 ? tmp14724 : tmp15102);
  assign tmp15096 = s3 ? tmp15097 : tmp15101;
  assign tmp15105 = s1 ? tmp14471 : tmp14444;
  assign tmp15104 = s2 ? tmp15105 : tmp14494;
  assign tmp15103 = s3 ? tmp15104 : tmp14741;
  assign tmp15095 = s4 ? tmp15096 : tmp15103;
  assign tmp15109 = s1 ? 1 : tmp14471;
  assign tmp15108 = s2 ? tmp14494 : tmp15109;
  assign tmp15107 = s3 ? tmp15108 : 1;
  assign tmp15111 = s2 ? 1 : tmp15105;
  assign tmp15110 = s3 ? tmp15111 : 1;
  assign tmp15106 = s4 ? tmp15107 : tmp15110;
  assign tmp15094 = s5 ? tmp15095 : tmp15106;
  assign tmp15089 = s6 ? tmp15090 : tmp15094;
  assign tmp15116 = s2 ? tmp15093 : tmp14720;
  assign tmp15117 = s2 ? 1 : tmp14493;
  assign tmp15115 = s3 ? tmp15116 : tmp15117;
  assign tmp15119 = s2 ? tmp15105 : 1;
  assign tmp15118 = s3 ? tmp15119 : tmp14741;
  assign tmp15114 = s4 ? tmp15115 : tmp15118;
  assign tmp15120 = s4 ? tmp14740 : tmp14480;
  assign tmp15113 = s5 ? tmp15114 : tmp15120;
  assign tmp15112 = s6 ? tmp15090 : tmp15113;
  assign tmp15088 = s7 ? tmp15089 : tmp15112;
  assign tmp15087 = s8 ? tmp15019 : tmp15088;
  assign tmp15018 = s9 ? tmp15019 : tmp15087;
  assign tmp15130 = ~(l1 ? 1 : tmp14706);
  assign tmp15129 = s0 ? tmp14421 : tmp15130;
  assign tmp15128 = s1 ? tmp15129 : tmp14421;
  assign tmp15127 = s2 ? tmp14421 : tmp15128;
  assign tmp15126 = s3 ? tmp14421 : tmp15127;
  assign tmp15132 = s2 ? tmp14421 : tmp14425;
  assign tmp15131 = s3 ? tmp15132 : tmp14429;
  assign tmp15125 = s4 ? tmp15126 : tmp15131;
  assign tmp15139 = l1 ? 1 : tmp14706;
  assign tmp15140 = ~(l1 ? 1 : tmp14422);
  assign tmp15138 = ~(s0 ? tmp15139 : tmp15140);
  assign tmp15137 = s1 ? tmp15129 : tmp15138;
  assign tmp15142 = s0 ? tmp15139 : tmp15140;
  assign tmp15143 = ~(s0 ? tmp14421 : tmp15130);
  assign tmp15141 = ~(s1 ? tmp15142 : tmp15143);
  assign tmp15136 = s2 ? tmp15137 : tmp15141;
  assign tmp15145 = ~(s1 ? 1 : tmp14439);
  assign tmp15144 = ~(s2 ? tmp15142 : tmp15145);
  assign tmp15135 = s3 ? tmp15136 : tmp15144;
  assign tmp15148 = s1 ? tmp14452 : tmp14444;
  assign tmp15149 = s1 ? tmp14444 : tmp14421;
  assign tmp15147 = s2 ? tmp15148 : tmp15149;
  assign tmp15146 = s3 ? tmp15147 : tmp14446;
  assign tmp15134 = s4 ? tmp15135 : tmp15146;
  assign tmp15152 = s2 ? tmp14447 : tmp14451;
  assign tmp15151 = s3 ? tmp15152 : 1;
  assign tmp15155 = s1 ? tmp14452 : tmp14439;
  assign tmp15154 = s2 ? 1 : tmp15155;
  assign tmp15153 = s3 ? tmp15154 : 1;
  assign tmp15150 = s4 ? tmp15151 : tmp15153;
  assign tmp15133 = s5 ? tmp15134 : tmp15150;
  assign tmp15124 = s6 ? tmp15125 : tmp15133;
  assign tmp15159 = s2 ? tmp14421 : tmp14428;
  assign tmp15158 = s3 ? tmp15159 : tmp14429;
  assign tmp15157 = s4 ? tmp15126 : tmp15158;
  assign tmp15164 = s1 ? tmp14421 : tmp15129;
  assign tmp15163 = s2 ? tmp15128 : tmp15164;
  assign tmp15162 = s3 ? tmp15163 : tmp14462;
  assign tmp15166 = s2 ? tmp15148 : tmp14421;
  assign tmp15165 = s3 ? tmp15166 : tmp14446;
  assign tmp15161 = s4 ? tmp15162 : tmp15165;
  assign tmp15169 = s2 ? tmp14447 : tmp14519;
  assign tmp15168 = s3 ? tmp15169 : tmp14469;
  assign tmp15167 = s4 ? tmp15168 : tmp14520;
  assign tmp15160 = s5 ? tmp15161 : tmp15167;
  assign tmp15156 = s6 ? tmp15157 : tmp15160;
  assign tmp15123 = s7 ? tmp15124 : tmp15156;
  assign tmp15122 = s8 ? tmp15123 : tmp15124;
  assign tmp15175 = s2 ? 1 : tmp15023;
  assign tmp15174 = s3 ? tmp15175 : 1;
  assign tmp15173 = s4 ? tmp15081 : tmp15174;
  assign tmp15172 = s5 ? tmp15072 : tmp15173;
  assign tmp15171 = s6 ? tmp15067 : tmp15172;
  assign tmp15178 = s4 ? tmp15168 : tmp14528;
  assign tmp15177 = s5 ? tmp15161 : tmp15178;
  assign tmp15176 = s6 ? tmp15157 : tmp15177;
  assign tmp15170 = s7 ? tmp15171 : tmp15176;
  assign tmp15121 = s9 ? tmp15122 : tmp15170;
  assign tmp15017 = s10 ? tmp15018 : tmp15121;
  assign tmp15181 = s7 ? tmp15066 : tmp15156;
  assign tmp15180 = s9 ? tmp15122 : tmp15181;
  assign tmp15179 = s10 ? tmp15018 : tmp15180;
  assign tmp15016 = s11 ? tmp15017 : tmp15179;
  assign tmp15015 = s12 ? tmp15016 : tmp14544;
  assign tmp14833 = s13 ? tmp14834 : tmp15015;
  assign tmp14692 = s14 ? tmp14693 : tmp14833;
  assign tmp15191 = s4 ? 1 : tmp14740;
  assign tmp15197 = s0 ? 1 : tmp15139;
  assign tmp15196 = s1 ? tmp15197 : 1;
  assign tmp15199 = s0 ? tmp15139 : 1;
  assign tmp15198 = s1 ? tmp15199 : 1;
  assign tmp15195 = s2 ? tmp15196 : tmp15198;
  assign tmp15194 = s3 ? tmp15195 : 1;
  assign tmp15201 = s2 ? tmp15109 : tmp15105;
  assign tmp15200 = s3 ? tmp15201 : 1;
  assign tmp15193 = s4 ? tmp15194 : tmp15200;
  assign tmp15192 = s5 ? tmp15193 : 1;
  assign tmp15190 = s6 ? tmp15191 : tmp15192;
  assign tmp15206 = s2 ? tmp15196 : 1;
  assign tmp15205 = s3 ? tmp15206 : 1;
  assign tmp15208 = s2 ? tmp15109 : 1;
  assign tmp15207 = s3 ? tmp15208 : 1;
  assign tmp15204 = s4 ? tmp15205 : tmp15207;
  assign tmp15203 = s5 ? tmp15204 : 1;
  assign tmp15202 = s6 ? tmp15191 : tmp15203;
  assign tmp15189 = s7 ? tmp15190 : tmp15202;
  assign tmp15214 = ~(l2 ? tmp14918 : 0);
  assign tmp15213 = l1 ? 1 : tmp15214;
  assign tmp15217 = s0 ? 1 : tmp15213;
  assign tmp15216 = s1 ? tmp15217 : tmp15213;
  assign tmp15215 = s2 ? tmp15216 : tmp15213;
  assign tmp15212 = s3 ? tmp15213 : tmp15215;
  assign tmp15221 = s0 ? tmp15213 : 0;
  assign tmp15220 = s1 ? tmp15221 : tmp15213;
  assign tmp15222 = s0 ? tmp15213 : 1;
  assign tmp15219 = s2 ? tmp15220 : tmp15222;
  assign tmp15224 = s1 ? tmp14918 : 0;
  assign tmp15225 = ~(l1 ? 1 : tmp15214);
  assign tmp15223 = ~(s2 ? tmp15224 : tmp15225);
  assign tmp15218 = s3 ? tmp15219 : tmp15223;
  assign tmp15211 = s4 ? tmp15212 : tmp15218;
  assign tmp15231 = s0 ? tmp15213 : tmp15139;
  assign tmp15230 = s1 ? tmp15231 : 1;
  assign tmp15233 = s0 ? tmp15139 : tmp15213;
  assign tmp15232 = s1 ? tmp15233 : tmp15213;
  assign tmp15229 = s2 ? tmp15230 : tmp15232;
  assign tmp15237 = l1 ? 1 : tmp14578;
  assign tmp15236 = s0 ? tmp15237 : 1;
  assign tmp15235 = s1 ? tmp15236 : tmp15213;
  assign tmp15234 = s2 ? tmp15213 : tmp15235;
  assign tmp15228 = s3 ? tmp15229 : tmp15234;
  assign tmp15241 = ~(s0 ? 1 : tmp14918);
  assign tmp15240 = s1 ? tmp15217 : tmp15241;
  assign tmp15243 = s0 ? 1 : tmp14918;
  assign tmp15244 = ~(s0 ? tmp15213 : 0);
  assign tmp15242 = ~(s1 ? tmp15243 : tmp15244);
  assign tmp15239 = s2 ? tmp15240 : tmp15242;
  assign tmp15247 = ~(s0 ? tmp14918 : 0);
  assign tmp15246 = s1 ? tmp15213 : tmp15247;
  assign tmp15245 = s2 ? tmp15246 : 1;
  assign tmp15238 = s3 ? tmp15239 : tmp15245;
  assign tmp15227 = s4 ? tmp15228 : tmp15238;
  assign tmp15252 = s0 ? 1 : tmp15237;
  assign tmp15251 = s1 ? tmp15222 : tmp15252;
  assign tmp15253 = s1 ? tmp15236 : 1;
  assign tmp15250 = s2 ? tmp15251 : tmp15253;
  assign tmp15249 = s3 ? tmp15250 : 1;
  assign tmp15256 = s1 ? 1 : tmp15252;
  assign tmp15257 = s1 ? tmp15217 : 1;
  assign tmp15255 = s2 ? tmp15256 : tmp15257;
  assign tmp15258 = s2 ? tmp15253 : 1;
  assign tmp15254 = s3 ? tmp15255 : tmp15258;
  assign tmp15248 = s4 ? tmp15249 : tmp15254;
  assign tmp15226 = s5 ? tmp15227 : tmp15248;
  assign tmp15210 = s6 ? tmp15211 : tmp15226;
  assign tmp15263 = s2 ? tmp15230 : tmp15213;
  assign tmp15262 = s3 ? tmp15263 : tmp15234;
  assign tmp15265 = s2 ? tmp15240 : tmp15213;
  assign tmp15267 = s1 ? tmp15213 : 1;
  assign tmp15266 = s2 ? tmp15267 : 1;
  assign tmp15264 = s3 ? tmp15265 : tmp15266;
  assign tmp15261 = s4 ? tmp15262 : tmp15264;
  assign tmp15271 = s1 ? tmp15222 : tmp15237;
  assign tmp15270 = s2 ? tmp15271 : tmp15253;
  assign tmp15269 = s3 ? tmp15270 : 1;
  assign tmp15274 = s1 ? 1 : tmp15237;
  assign tmp15273 = s2 ? tmp15274 : tmp15213;
  assign tmp15272 = s3 ? tmp15273 : tmp15253;
  assign tmp15268 = s4 ? tmp15269 : tmp15272;
  assign tmp15260 = s5 ? tmp15261 : tmp15268;
  assign tmp15259 = s6 ? tmp15211 : tmp15260;
  assign tmp15209 = s7 ? tmp15210 : tmp15259;
  assign tmp15188 = s8 ? tmp15189 : tmp15209;
  assign tmp15281 = s1 ? tmp15231 : tmp15213;
  assign tmp15280 = s2 ? tmp15281 : tmp15222;
  assign tmp15279 = s3 ? tmp15280 : tmp15223;
  assign tmp15278 = s4 ? tmp15212 : tmp15279;
  assign tmp15287 = ~(s0 ? tmp15213 : tmp15139);
  assign tmp15286 = ~(s1 ? tmp15243 : tmp15287);
  assign tmp15285 = s2 ? tmp15240 : tmp15286;
  assign tmp15284 = s3 ? tmp15285 : tmp15245;
  assign tmp15283 = s4 ? tmp15228 : tmp15284;
  assign tmp15282 = s5 ? tmp15283 : tmp15248;
  assign tmp15277 = s6 ? tmp15278 : tmp15282;
  assign tmp15288 = s6 ? tmp15278 : tmp15260;
  assign tmp15276 = s7 ? tmp15277 : tmp15288;
  assign tmp15294 = s2 ? tmp14494 : tmp14470;
  assign tmp15293 = s3 ? tmp15294 : 1;
  assign tmp15292 = s4 ? tmp15293 : tmp15200;
  assign tmp15291 = s5 ? tmp15292 : 1;
  assign tmp15290 = s6 ? tmp15191 : tmp15291;
  assign tmp15297 = s4 ? tmp14740 : tmp15207;
  assign tmp15296 = s5 ? tmp15297 : 1;
  assign tmp15295 = s6 ? tmp15191 : tmp15296;
  assign tmp15289 = s7 ? tmp15290 : tmp15295;
  assign tmp15275 = s8 ? tmp15276 : tmp15289;
  assign tmp15187 = s9 ? tmp15188 : tmp15275;
  assign tmp15302 = s4 ? 1 : tmp15205;
  assign tmp15307 = s1 ? tmp14471 : tmp15197;
  assign tmp15306 = s2 ? tmp15109 : tmp15307;
  assign tmp15305 = s3 ? tmp15306 : 1;
  assign tmp15304 = s4 ? tmp15194 : tmp15305;
  assign tmp15303 = s5 ? tmp15304 : 1;
  assign tmp15301 = s6 ? tmp15302 : tmp15303;
  assign tmp15308 = s6 ? tmp15302 : tmp15203;
  assign tmp15300 = s7 ? tmp15301 : tmp15308;
  assign tmp15299 = s8 ? tmp15300 : tmp15301;
  assign tmp15310 = s7 ? tmp15202 : tmp15295;
  assign tmp15315 = s3 ? tmp15273 : 1;
  assign tmp15314 = s4 ? tmp15269 : tmp15315;
  assign tmp15313 = s5 ? tmp15261 : tmp15314;
  assign tmp15312 = s6 ? tmp15278 : tmp15313;
  assign tmp15311 = s7 ? tmp15312 : tmp15308;
  assign tmp15309 = s8 ? tmp15310 : tmp15311;
  assign tmp15298 = s9 ? tmp15299 : tmp15309;
  assign tmp15186 = s10 ? tmp15187 : tmp15298;
  assign tmp15319 = s7 ? tmp15288 : tmp15308;
  assign tmp15318 = s8 ? tmp15310 : tmp15319;
  assign tmp15317 = s9 ? tmp15299 : tmp15318;
  assign tmp15316 = s10 ? tmp15187 : tmp15317;
  assign tmp15185 = s11 ? tmp15186 : tmp15316;
  assign tmp15184 = s12 ? tmp14567 : tmp15185;
  assign tmp15183 = s13 ? tmp15184 : 1;
  assign tmp15182 = s14 ? 1 : tmp15183;
  assign tmp14691 = s15 ? tmp14692 : tmp15182;
  assign tmp15333 = s2 ? tmp15148 : tmp14445;
  assign tmp15335 = s1 ? tmp14439 : tmp14471;
  assign tmp15334 = s2 ? tmp15335 : 1;
  assign tmp15332 = s3 ? tmp15333 : tmp15334;
  assign tmp15331 = s4 ? tmp14433 : tmp15332;
  assign tmp15338 = s2 ? tmp14428 : tmp14452;
  assign tmp15337 = s3 ? tmp15338 : 1;
  assign tmp15340 = s2 ? tmp14510 : tmp14455;
  assign tmp15339 = s3 ? tmp15340 : 1;
  assign tmp15336 = s4 ? tmp15337 : tmp15339;
  assign tmp15330 = s5 ? tmp15331 : tmp15336;
  assign tmp15329 = s6 ? tmp14418 : tmp15330;
  assign tmp15343 = s4 ? tmp14459 : tmp15165;
  assign tmp15342 = s5 ? tmp15343 : tmp14465;
  assign tmp15341 = s6 ? tmp14418 : tmp15342;
  assign tmp15328 = s7 ? tmp15329 : tmp15341;
  assign tmp15349 = s2 ? tmp14420 : tmp14510;
  assign tmp15348 = s3 ? tmp14434 : tmp15349;
  assign tmp15352 = s1 ? tmp14452 : 1;
  assign tmp15351 = s2 ? tmp15352 : tmp14500;
  assign tmp15353 = s2 ? tmp14519 : 1;
  assign tmp15350 = s3 ? tmp15351 : tmp15353;
  assign tmp15347 = s4 ? tmp15348 : tmp15350;
  assign tmp15346 = s5 ? tmp15347 : tmp14448;
  assign tmp15345 = s6 ? tmp14418 : tmp15346;
  assign tmp15358 = s2 ? tmp14421 : tmp14510;
  assign tmp15357 = s3 ? tmp14460 : tmp15358;
  assign tmp15360 = s2 ? tmp15352 : tmp14421;
  assign tmp15359 = s3 ? tmp15360 : tmp15353;
  assign tmp15356 = s4 ? tmp15357 : tmp15359;
  assign tmp15355 = s5 ? tmp15356 : tmp14465;
  assign tmp15354 = s6 ? tmp14418 : tmp15355;
  assign tmp15344 = s7 ? tmp15345 : tmp15354;
  assign tmp15327 = s8 ? tmp15328 : tmp15344;
  assign tmp15366 = s3 ? tmp14469 : 1;
  assign tmp15365 = s4 ? 1 : tmp15366;
  assign tmp15364 = s5 ? tmp15365 : tmp14497;
  assign tmp15363 = s6 ? 1 : tmp15364;
  assign tmp15371 = s2 ? tmp14428 : 1;
  assign tmp15370 = s3 ? tmp14499 : tmp15371;
  assign tmp15369 = s4 ? tmp15370 : tmp14501;
  assign tmp15368 = s5 ? tmp15365 : tmp15369;
  assign tmp15367 = s6 ? 1 : tmp15368;
  assign tmp15362 = s7 ? tmp15363 : tmp15367;
  assign tmp15361 = s8 ? tmp15344 : tmp15362;
  assign tmp15326 = s9 ? tmp15327 : tmp15361;
  assign tmp15373 = s8 ? tmp15344 : tmp15345;
  assign tmp15377 = s5 ? tmp15343 : tmp14527;
  assign tmp15376 = s6 ? tmp14418 : tmp15377;
  assign tmp15380 = s4 ? tmp15370 : 1;
  assign tmp15379 = s5 ? tmp15365 : tmp15380;
  assign tmp15378 = s6 ? 1 : tmp15379;
  assign tmp15375 = s7 ? tmp15376 : tmp15378;
  assign tmp15382 = s5 ? tmp15356 : tmp14527;
  assign tmp15381 = s6 ? tmp14418 : tmp15382;
  assign tmp15374 = s8 ? tmp15375 : tmp15381;
  assign tmp15372 = s9 ? tmp15373 : tmp15374;
  assign tmp15325 = s10 ? tmp15326 : tmp15372;
  assign tmp15386 = s7 ? tmp15341 : tmp15367;
  assign tmp15385 = s8 ? tmp15386 : tmp15354;
  assign tmp15384 = s9 ? tmp15373 : tmp15385;
  assign tmp15383 = s10 ? tmp15326 : tmp15384;
  assign tmp15324 = s11 ? tmp15325 : tmp15383;
  assign tmp15323 = s12 ? tmp15324 : tmp14544;
  assign tmp15322 = s13 ? 1 : tmp15323;
  assign tmp15321 = s14 ? 1 : tmp15322;
  assign tmp15320 = s15 ? tmp15321 : tmp14564;
  assign tmp14690 = s16 ? tmp14691 : tmp15320;
  assign tmp14406 = ~(s17 ? tmp14407 : tmp14690);
  assign s17n = tmp14406;

  assign tmp15404 = ~(l2 ? 1 : 0);
  assign tmp15403 = s0 ? 1 : tmp15404;
  assign tmp15402 = s1 ? tmp15403 : 1;
  assign tmp15401 = s2 ? tmp15402 : 1;
  assign tmp15400 = s3 ? tmp15401 : 1;
  assign tmp15409 = l2 ? 1 : 0;
  assign tmp15408 = s0 ? tmp15409 : 0;
  assign tmp15407 = ~(s1 ? tmp15408 : 0);
  assign tmp15406 = s2 ? 1 : tmp15407;
  assign tmp15405 = s3 ? tmp15406 : 1;
  assign tmp15399 = s4 ? tmp15400 : tmp15405;
  assign tmp15398 = s5 ? 1 : tmp15399;
  assign tmp15397 = s6 ? 1 : tmp15398;
  assign tmp15412 = s4 ? tmp15400 : 1;
  assign tmp15411 = s5 ? 1 : tmp15412;
  assign tmp15410 = s6 ? 1 : tmp15411;
  assign tmp15396 = s7 ? tmp15397 : tmp15410;
  assign tmp15421 = ~(l1 ? 1 : 0);
  assign tmp15420 = s0 ? 1 : tmp15421;
  assign tmp15419 = s1 ? 1 : tmp15420;
  assign tmp15418 = s2 ? 1 : tmp15419;
  assign tmp15424 = l1 ? 1 : 0;
  assign tmp15423 = s0 ? tmp15424 : 0;
  assign tmp15422 = ~(s2 ? tmp15423 : 0);
  assign tmp15417 = s3 ? tmp15418 : tmp15422;
  assign tmp15416 = s4 ? tmp15417 : 1;
  assign tmp15415 = s5 ? tmp15416 : tmp15399;
  assign tmp15414 = s6 ? 1 : tmp15415;
  assign tmp15428 = s3 ? tmp15418 : 1;
  assign tmp15432 = l1 ? tmp15409 : 0;
  assign tmp15434 = ~(l1 ? tmp15409 : 0);
  assign tmp15433 = ~(s0 ? 1 : tmp15434);
  assign tmp15431 = ~(s1 ? tmp15432 : tmp15433);
  assign tmp15430 = s2 ? 1 : tmp15431;
  assign tmp15429 = s3 ? tmp15430 : 1;
  assign tmp15427 = s4 ? tmp15428 : tmp15429;
  assign tmp15426 = s5 ? tmp15427 : tmp15412;
  assign tmp15425 = s6 ? 1 : tmp15426;
  assign tmp15413 = s7 ? tmp15414 : tmp15425;
  assign tmp15395 = s8 ? tmp15396 : tmp15413;
  assign tmp15441 = s0 ? tmp15432 : tmp15409;
  assign tmp15440 = s2 ? tmp15432 : tmp15441;
  assign tmp15443 = s1 ? tmp15432 : tmp15408;
  assign tmp15444 = s1 ? tmp15432 : tmp15433;
  assign tmp15442 = s2 ? tmp15443 : tmp15444;
  assign tmp15439 = s3 ? tmp15440 : tmp15442;
  assign tmp15438 = s4 ? tmp15432 : tmp15439;
  assign tmp15450 = s0 ? tmp15432 : 0;
  assign tmp15449 = s1 ? tmp15450 : tmp15433;
  assign tmp15452 = s0 ? 1 : tmp15434;
  assign tmp15451 = ~(s1 ? tmp15452 : tmp15434);
  assign tmp15448 = s2 ? tmp15449 : tmp15451;
  assign tmp15454 = s1 ? tmp15432 : tmp15423;
  assign tmp15456 = ~(s0 ? tmp15432 : tmp15409);
  assign tmp15455 = ~(s1 ? 1 : tmp15456);
  assign tmp15453 = s2 ? tmp15454 : tmp15455;
  assign tmp15447 = s3 ? tmp15448 : tmp15453;
  assign tmp15459 = s1 ? tmp15452 : tmp15456;
  assign tmp15460 = ~(s1 ? tmp15441 : tmp15432);
  assign tmp15458 = s2 ? tmp15459 : tmp15460;
  assign tmp15463 = ~(s0 ? tmp15409 : 0);
  assign tmp15462 = s1 ? tmp15403 : tmp15463;
  assign tmp15461 = s2 ? tmp15462 : 1;
  assign tmp15457 = ~(s3 ? tmp15458 : tmp15461);
  assign tmp15446 = s4 ? tmp15447 : tmp15457;
  assign tmp15468 = s0 ? 1 : tmp15424;
  assign tmp15467 = s1 ? tmp15468 : 1;
  assign tmp15466 = s2 ? tmp15467 : 1;
  assign tmp15465 = s3 ? tmp15466 : 1;
  assign tmp15472 = s0 ? tmp15424 : 1;
  assign tmp15471 = s1 ? tmp15472 : 1;
  assign tmp15470 = s2 ? 1 : tmp15471;
  assign tmp15469 = s3 ? tmp15470 : 1;
  assign tmp15464 = ~(s4 ? tmp15465 : tmp15469);
  assign tmp15445 = s5 ? tmp15446 : tmp15464;
  assign tmp15437 = s6 ? tmp15438 : tmp15445;
  assign tmp15477 = s1 ? tmp15441 : tmp15432;
  assign tmp15476 = s2 ? tmp15432 : tmp15477;
  assign tmp15479 = s1 ? tmp15432 : 0;
  assign tmp15478 = s2 ? tmp15479 : tmp15444;
  assign tmp15475 = s3 ? tmp15476 : tmp15478;
  assign tmp15474 = s4 ? tmp15432 : tmp15475;
  assign tmp15484 = s1 ? tmp15450 : tmp15432;
  assign tmp15483 = s2 ? tmp15484 : tmp15432;
  assign tmp15485 = s2 ? tmp15479 : tmp15455;
  assign tmp15482 = s3 ? tmp15483 : tmp15485;
  assign tmp15487 = s2 ? tmp15459 : tmp15434;
  assign tmp15486 = ~(s3 ? tmp15487 : tmp15401);
  assign tmp15481 = s4 ? tmp15482 : tmp15486;
  assign tmp15488 = ~(s4 ? tmp15465 : 1);
  assign tmp15480 = s5 ? tmp15481 : tmp15488;
  assign tmp15473 = s6 ? tmp15474 : tmp15480;
  assign tmp15436 = ~(s7 ? tmp15437 : tmp15473);
  assign tmp15435 = s8 ? tmp15413 : tmp15436;
  assign tmp15394 = s9 ? tmp15395 : tmp15435;
  assign tmp15498 = ~(s0 ? tmp15432 : tmp15424);
  assign tmp15497 = ~(s1 ? tmp15452 : tmp15498);
  assign tmp15496 = s2 ? tmp15449 : tmp15497;
  assign tmp15501 = s0 ? tmp15424 : tmp15432;
  assign tmp15500 = s1 ? tmp15501 : tmp15423;
  assign tmp15502 = ~(s1 ? 1 : tmp15434);
  assign tmp15499 = s2 ? tmp15500 : tmp15502;
  assign tmp15495 = s3 ? tmp15496 : tmp15499;
  assign tmp15505 = s1 ? tmp15452 : tmp15463;
  assign tmp15504 = s2 ? tmp15505 : 1;
  assign tmp15503 = ~(s3 ? tmp15458 : tmp15504);
  assign tmp15494 = s4 ? tmp15495 : tmp15503;
  assign tmp15506 = ~(s4 ? tmp15400 : tmp15405);
  assign tmp15493 = s5 ? tmp15494 : tmp15506;
  assign tmp15492 = s6 ? tmp15438 : tmp15493;
  assign tmp15513 = s0 ? tmp15432 : tmp15424;
  assign tmp15512 = s1 ? tmp15432 : tmp15513;
  assign tmp15511 = s2 ? tmp15484 : tmp15512;
  assign tmp15514 = s2 ? tmp15479 : tmp15502;
  assign tmp15510 = s3 ? tmp15511 : tmp15514;
  assign tmp15517 = s1 ? tmp15452 : 1;
  assign tmp15516 = s2 ? tmp15517 : 1;
  assign tmp15515 = ~(s3 ? tmp15487 : tmp15516);
  assign tmp15509 = s4 ? tmp15510 : tmp15515;
  assign tmp15518 = ~(s4 ? tmp15400 : 1);
  assign tmp15508 = s5 ? tmp15509 : tmp15518;
  assign tmp15507 = s6 ? tmp15474 : tmp15508;
  assign tmp15491 = s7 ? tmp15492 : tmp15507;
  assign tmp15490 = s8 ? tmp15491 : tmp15492;
  assign tmp15521 = ~(s6 ? tmp15474 : tmp15480);
  assign tmp15520 = s7 ? tmp15410 : tmp15521;
  assign tmp15528 = ~(s1 ? tmp15432 : 0);
  assign tmp15527 = s2 ? 1 : tmp15528;
  assign tmp15526 = s3 ? tmp15527 : 1;
  assign tmp15525 = s4 ? tmp15428 : tmp15526;
  assign tmp15524 = s5 ? tmp15525 : tmp15412;
  assign tmp15523 = s6 ? 1 : tmp15524;
  assign tmp15529 = ~(s6 ? tmp15474 : tmp15508);
  assign tmp15522 = s7 ? tmp15523 : tmp15529;
  assign tmp15519 = ~(s8 ? tmp15520 : tmp15522);
  assign tmp15489 = ~(s9 ? tmp15490 : tmp15519);
  assign tmp15393 = s10 ? tmp15394 : tmp15489;
  assign tmp15533 = s7 ? tmp15425 : tmp15529;
  assign tmp15532 = ~(s8 ? tmp15520 : tmp15533);
  assign tmp15531 = ~(s9 ? tmp15490 : tmp15532);
  assign tmp15530 = s10 ? tmp15394 : tmp15531;
  assign tmp15392 = s11 ? tmp15393 : tmp15530;
  assign tmp15545 = s0 ? 1 : 0;
  assign tmp15544 = s1 ? 1 : tmp15545;
  assign tmp15547 = ~(s0 ? 1 : 0);
  assign tmp15546 = s1 ? 1 : tmp15547;
  assign tmp15543 = s2 ? tmp15544 : tmp15546;
  assign tmp15542 = s3 ? 1 : tmp15543;
  assign tmp15541 = s4 ? 1 : tmp15542;
  assign tmp15552 = ~(s1 ? 1 : tmp15547);
  assign tmp15551 = s2 ? tmp15544 : tmp15552;
  assign tmp15550 = s3 ? 1 : tmp15551;
  assign tmp15555 = s1 ? tmp15545 : tmp15547;
  assign tmp15556 = ~(s1 ? tmp15545 : 1);
  assign tmp15554 = s2 ? tmp15555 : tmp15556;
  assign tmp15553 = ~(s3 ? tmp15554 : 1);
  assign tmp15549 = s4 ? tmp15550 : tmp15553;
  assign tmp15548 = s5 ? tmp15549 : 0;
  assign tmp15540 = s6 ? tmp15541 : tmp15548;
  assign tmp15562 = s1 ? 1 : 0;
  assign tmp15561 = s2 ? tmp15562 : tmp15552;
  assign tmp15560 = s3 ? 1 : tmp15561;
  assign tmp15564 = s2 ? tmp15555 : 0;
  assign tmp15563 = ~(s3 ? tmp15564 : 1);
  assign tmp15559 = s4 ? tmp15560 : tmp15563;
  assign tmp15558 = s5 ? tmp15559 : 0;
  assign tmp15557 = s6 ? tmp15541 : tmp15558;
  assign tmp15539 = s7 ? tmp15540 : tmp15557;
  assign tmp15571 = ~(s1 ? 1 : 0);
  assign tmp15570 = s2 ? tmp15544 : tmp15571;
  assign tmp15569 = s3 ? 1 : tmp15570;
  assign tmp15574 = s1 ? tmp15545 : 0;
  assign tmp15573 = s2 ? tmp15574 : 0;
  assign tmp15572 = ~(s3 ? tmp15573 : 1);
  assign tmp15568 = s4 ? tmp15569 : tmp15572;
  assign tmp15567 = s5 ? tmp15568 : 0;
  assign tmp15566 = s6 ? tmp15541 : tmp15567;
  assign tmp15579 = s1 ? 1 : tmp15452;
  assign tmp15578 = s2 ? 1 : tmp15579;
  assign tmp15582 = ~(s0 ? tmp15432 : 1);
  assign tmp15581 = s1 ? 1 : tmp15582;
  assign tmp15580 = s2 ? tmp15581 : tmp15546;
  assign tmp15577 = s3 ? tmp15578 : tmp15580;
  assign tmp15576 = s4 ? 1 : tmp15577;
  assign tmp15586 = s2 ? tmp15562 : tmp15571;
  assign tmp15585 = s3 ? 1 : tmp15586;
  assign tmp15584 = s4 ? tmp15585 : tmp15572;
  assign tmp15583 = s5 ? tmp15584 : 0;
  assign tmp15575 = s6 ? tmp15576 : tmp15583;
  assign tmp15565 = s7 ? tmp15566 : tmp15575;
  assign tmp15538 = s8 ? tmp15539 : tmp15565;
  assign tmp15594 = s0 ? tmp15432 : 1;
  assign tmp15593 = s1 ? tmp15432 : tmp15594;
  assign tmp15596 = s0 ? 1 : tmp15432;
  assign tmp15595 = s1 ? tmp15432 : tmp15596;
  assign tmp15592 = s2 ? tmp15593 : tmp15595;
  assign tmp15591 = s3 ? tmp15432 : tmp15592;
  assign tmp15590 = s4 ? tmp15432 : tmp15591;
  assign tmp15601 = ~(s1 ? tmp15403 : tmp15421);
  assign tmp15600 = s2 ? tmp15449 : tmp15601;
  assign tmp15603 = s1 ? tmp15424 : tmp15472;
  assign tmp15604 = s1 ? 1 : tmp15409;
  assign tmp15602 = s2 ? tmp15603 : tmp15604;
  assign tmp15599 = s3 ? tmp15600 : tmp15602;
  assign tmp15608 = s0 ? 1 : tmp15409;
  assign tmp15607 = s1 ? tmp15608 : tmp15409;
  assign tmp15606 = s2 ? tmp15607 : tmp15409;
  assign tmp15605 = s3 ? tmp15606 : 1;
  assign tmp15598 = s4 ? tmp15599 : tmp15605;
  assign tmp15597 = s5 ? tmp15598 : 1;
  assign tmp15589 = s6 ? tmp15590 : tmp15597;
  assign tmp15614 = s1 ? tmp15409 : tmp15424;
  assign tmp15613 = s2 ? tmp15484 : tmp15614;
  assign tmp15616 = s1 ? tmp15424 : 1;
  assign tmp15615 = s2 ? tmp15616 : tmp15604;
  assign tmp15612 = s3 ? tmp15613 : tmp15615;
  assign tmp15611 = s4 ? tmp15612 : tmp15605;
  assign tmp15610 = s5 ? tmp15611 : 1;
  assign tmp15609 = s6 ? tmp15590 : tmp15610;
  assign tmp15588 = ~(s7 ? tmp15589 : tmp15609);
  assign tmp15587 = s8 ? tmp15565 : tmp15588;
  assign tmp15537 = s9 ? tmp15538 : tmp15587;
  assign tmp15619 = s7 ? tmp15589 : tmp15609;
  assign tmp15618 = s8 ? tmp15619 : tmp15589;
  assign tmp15625 = s2 ? tmp15562 : tmp15546;
  assign tmp15624 = s3 ? 1 : tmp15625;
  assign tmp15623 = s4 ? 1 : tmp15624;
  assign tmp15622 = s6 ? tmp15623 : tmp15558;
  assign tmp15630 = s1 ? tmp15432 : 1;
  assign tmp15629 = s2 ? tmp15630 : tmp15595;
  assign tmp15628 = s3 ? tmp15432 : tmp15629;
  assign tmp15627 = s4 ? tmp15432 : tmp15628;
  assign tmp15626 = ~(s6 ? tmp15627 : tmp15610);
  assign tmp15621 = s7 ? tmp15622 : tmp15626;
  assign tmp15634 = s3 ? tmp15578 : tmp15625;
  assign tmp15633 = s4 ? 1 : tmp15634;
  assign tmp15632 = s6 ? tmp15633 : tmp15583;
  assign tmp15631 = s7 ? tmp15632 : tmp15626;
  assign tmp15620 = ~(s8 ? tmp15621 : tmp15631);
  assign tmp15617 = ~(s9 ? tmp15618 : tmp15620);
  assign tmp15536 = s10 ? tmp15537 : tmp15617;
  assign tmp15639 = ~(s6 ? tmp15590 : tmp15610);
  assign tmp15638 = s7 ? tmp15557 : tmp15639;
  assign tmp15640 = s7 ? tmp15575 : tmp15639;
  assign tmp15637 = ~(s8 ? tmp15638 : tmp15640);
  assign tmp15636 = ~(s9 ? tmp15618 : tmp15637);
  assign tmp15635 = s10 ? tmp15537 : tmp15636;
  assign tmp15535 = s11 ? tmp15536 : tmp15635;
  assign tmp15534 = s12 ? 1 : tmp15535;
  assign tmp15391 = s13 ? tmp15392 : tmp15534;
  assign tmp15654 = ~(s0 ? 1 : tmp15421);
  assign tmp15653 = s1 ? tmp15423 : tmp15654;
  assign tmp15655 = ~(s1 ? tmp15420 : tmp15421);
  assign tmp15652 = s2 ? tmp15653 : tmp15655;
  assign tmp15657 = s1 ? tmp15424 : tmp15423;
  assign tmp15656 = s2 ? tmp15657 : tmp15472;
  assign tmp15651 = s3 ? tmp15652 : tmp15656;
  assign tmp15660 = s1 ? tmp15472 : tmp15424;
  assign tmp15659 = s2 ? tmp15603 : tmp15660;
  assign tmp15661 = ~(s1 ? tmp15545 : 0);
  assign tmp15658 = s3 ? tmp15659 : tmp15661;
  assign tmp15650 = s4 ? tmp15651 : tmp15658;
  assign tmp15649 = s5 ? tmp15650 : 0;
  assign tmp15648 = s6 ? tmp15424 : tmp15649;
  assign tmp15667 = s1 ? tmp15423 : tmp15424;
  assign tmp15666 = s2 ? tmp15667 : tmp15424;
  assign tmp15672 = l3 ? 1 : 0;
  assign tmp15671 = ~(l2 ? tmp15672 : 1);
  assign tmp15670 = l1 ? 1 : tmp15671;
  assign tmp15673 = s0 ? tmp15670 : 0;
  assign tmp15669 = s1 ? tmp15670 : tmp15673;
  assign tmp15668 = s2 ? tmp15669 : tmp15472;
  assign tmp15665 = s3 ? tmp15666 : tmp15668;
  assign tmp15675 = s2 ? tmp15603 : tmp15424;
  assign tmp15676 = ~(s2 ? tmp15545 : 1);
  assign tmp15674 = s3 ? tmp15675 : tmp15676;
  assign tmp15664 = s4 ? tmp15665 : tmp15674;
  assign tmp15663 = s5 ? tmp15664 : 0;
  assign tmp15662 = s6 ? tmp15424 : tmp15663;
  assign tmp15647 = ~(s7 ? tmp15648 : tmp15662);
  assign tmp15646 = s8 ? 1 : tmp15647;
  assign tmp15645 = s9 ? tmp15646 : tmp15647;
  assign tmp15679 = s7 ? tmp15648 : tmp15662;
  assign tmp15678 = s8 ? tmp15679 : tmp15648;
  assign tmp15687 = s1 ? tmp15670 : 0;
  assign tmp15686 = s2 ? tmp15687 : tmp15472;
  assign tmp15685 = s3 ? tmp15666 : tmp15686;
  assign tmp15684 = s4 ? tmp15685 : tmp15674;
  assign tmp15683 = s5 ? tmp15684 : 0;
  assign tmp15682 = ~(s6 ? tmp15424 : tmp15683);
  assign tmp15681 = s7 ? 1 : tmp15682;
  assign tmp15680 = ~(s8 ? tmp15681 : tmp15682);
  assign tmp15677 = ~(s9 ? tmp15678 : tmp15680);
  assign tmp15644 = s10 ? tmp15645 : tmp15677;
  assign tmp15692 = ~(s6 ? tmp15424 : tmp15663);
  assign tmp15691 = s7 ? 1 : tmp15692;
  assign tmp15690 = ~(s8 ? tmp15691 : tmp15692);
  assign tmp15689 = ~(s9 ? tmp15678 : tmp15690);
  assign tmp15688 = s10 ? tmp15645 : tmp15689;
  assign tmp15643 = s11 ? tmp15644 : tmp15688;
  assign tmp15702 = s1 ? tmp15545 : 1;
  assign tmp15701 = s2 ? 1 : tmp15702;
  assign tmp15700 = s3 ? 1 : tmp15701;
  assign tmp15704 = s2 ? 1 : tmp15545;
  assign tmp15705 = s2 ? tmp15546 : 1;
  assign tmp15703 = s3 ? tmp15704 : tmp15705;
  assign tmp15699 = s4 ? tmp15700 : tmp15703;
  assign tmp15710 = ~(s1 ? tmp15545 : tmp15547);
  assign tmp15709 = s2 ? tmp15555 : tmp15710;
  assign tmp15711 = ~(s2 ? tmp15545 : 0);
  assign tmp15708 = s3 ? tmp15709 : tmp15711;
  assign tmp15707 = s4 ? tmp15708 : 1;
  assign tmp15706 = s5 ? tmp15707 : 1;
  assign tmp15698 = s6 ? tmp15699 : tmp15706;
  assign tmp15714 = s3 ? tmp15701 : 1;
  assign tmp15713 = s4 ? tmp15700 : tmp15714;
  assign tmp15718 = s2 ? tmp15702 : tmp15544;
  assign tmp15717 = s3 ? tmp15718 : 1;
  assign tmp15716 = s4 ? tmp15717 : 1;
  assign tmp15715 = s5 ? tmp15716 : 1;
  assign tmp15712 = s6 ? tmp15713 : tmp15715;
  assign tmp15697 = s7 ? tmp15698 : tmp15712;
  assign tmp15726 = l4 ? 1 : 0;
  assign tmp15725 = l2 ? tmp15726 : 0;
  assign tmp15724 = l1 ? tmp15409 : tmp15725;
  assign tmp15728 = l1 ? tmp15409 : tmp15726;
  assign tmp15727 = s0 ? tmp15728 : tmp15724;
  assign tmp15723 = s1 ? tmp15724 : tmp15727;
  assign tmp15731 = s0 ? tmp15724 : 1;
  assign tmp15730 = s1 ? tmp15731 : tmp15724;
  assign tmp15729 = s2 ? tmp15724 : tmp15730;
  assign tmp15722 = s3 ? tmp15723 : tmp15729;
  assign tmp15735 = s0 ? tmp15724 : tmp15409;
  assign tmp15734 = s1 ? tmp15735 : tmp15724;
  assign tmp15737 = s0 ? tmp15728 : 1;
  assign tmp15736 = s1 ? tmp15731 : tmp15737;
  assign tmp15733 = s2 ? tmp15734 : tmp15736;
  assign tmp15739 = s1 ? tmp15728 : tmp15545;
  assign tmp15741 = s0 ? tmp15726 : tmp15724;
  assign tmp15740 = s1 ? tmp15724 : tmp15741;
  assign tmp15738 = s2 ? tmp15739 : tmp15740;
  assign tmp15732 = s3 ? tmp15733 : tmp15738;
  assign tmp15721 = s4 ? tmp15722 : tmp15732;
  assign tmp15746 = s1 ? tmp15731 : tmp15608;
  assign tmp15748 = s0 ? 1 : tmp15724;
  assign tmp15747 = s1 ? tmp15748 : tmp15731;
  assign tmp15745 = s2 ? tmp15746 : tmp15747;
  assign tmp15751 = s0 ? tmp15726 : 0;
  assign tmp15750 = s1 ? tmp15751 : tmp15724;
  assign tmp15749 = s2 ? tmp15748 : tmp15750;
  assign tmp15744 = s3 ? tmp15745 : tmp15749;
  assign tmp15756 = ~(l1 ? tmp15409 : tmp15725);
  assign tmp15755 = s0 ? 1 : tmp15756;
  assign tmp15758 = l1 ? tmp15409 : 1;
  assign tmp15757 = ~(s0 ? tmp15758 : tmp15728);
  assign tmp15754 = s1 ? tmp15755 : tmp15757;
  assign tmp15760 = s0 ? tmp15758 : tmp15728;
  assign tmp15759 = ~(s1 ? tmp15760 : tmp15735);
  assign tmp15753 = s2 ? tmp15754 : tmp15759;
  assign tmp15763 = s0 ? tmp15728 : 0;
  assign tmp15762 = s1 ? tmp15724 : tmp15763;
  assign tmp15761 = ~(s2 ? tmp15762 : 0);
  assign tmp15752 = ~(s3 ? tmp15753 : tmp15761);
  assign tmp15743 = s4 ? tmp15744 : tmp15752;
  assign tmp15768 = s0 ? tmp15724 : 0;
  assign tmp15770 = ~(l4 ? 1 : 0);
  assign tmp15769 = ~(s0 ? 1 : tmp15770);
  assign tmp15767 = s1 ? tmp15768 : tmp15769;
  assign tmp15772 = s0 ? tmp15726 : tmp15409;
  assign tmp15771 = s1 ? tmp15772 : tmp15409;
  assign tmp15766 = s2 ? tmp15767 : tmp15771;
  assign tmp15765 = s3 ? tmp15766 : 0;
  assign tmp15776 = s0 ? 1 : tmp15770;
  assign tmp15775 = s1 ? 1 : tmp15776;
  assign tmp15777 = s1 ? tmp15755 : tmp15404;
  assign tmp15774 = s2 ? tmp15775 : tmp15777;
  assign tmp15779 = s1 ? tmp15751 : 0;
  assign tmp15778 = ~(s2 ? tmp15779 : 0);
  assign tmp15773 = ~(s3 ? tmp15774 : tmp15778);
  assign tmp15764 = s4 ? tmp15765 : tmp15773;
  assign tmp15742 = s5 ? tmp15743 : tmp15764;
  assign tmp15720 = s6 ? tmp15721 : tmp15742;
  assign tmp15784 = s1 ? tmp15731 : tmp15728;
  assign tmp15783 = s2 ? tmp15734 : tmp15784;
  assign tmp15786 = s1 ? tmp15728 : 0;
  assign tmp15785 = s2 ? tmp15786 : tmp15740;
  assign tmp15782 = s3 ? tmp15783 : tmp15785;
  assign tmp15781 = s4 ? tmp15722 : tmp15782;
  assign tmp15791 = s1 ? tmp15731 : tmp15409;
  assign tmp15792 = s1 ? tmp15724 : tmp15731;
  assign tmp15790 = s2 ? tmp15791 : tmp15792;
  assign tmp15793 = s2 ? tmp15724 : tmp15750;
  assign tmp15789 = s3 ? tmp15790 : tmp15793;
  assign tmp15796 = ~(s1 ? tmp15728 : tmp15724);
  assign tmp15795 = s2 ? tmp15754 : tmp15796;
  assign tmp15794 = ~(s3 ? tmp15795 : tmp15761);
  assign tmp15788 = s4 ? tmp15789 : tmp15794;
  assign tmp15800 = s1 ? tmp15768 : tmp15726;
  assign tmp15801 = s1 ? tmp15409 : 0;
  assign tmp15799 = s2 ? tmp15800 : tmp15801;
  assign tmp15798 = s3 ? tmp15799 : 0;
  assign tmp15804 = s1 ? 1 : tmp15770;
  assign tmp15803 = s2 ? tmp15804 : tmp15756;
  assign tmp15802 = ~(s3 ? tmp15803 : 1);
  assign tmp15797 = s4 ? tmp15798 : tmp15802;
  assign tmp15787 = s5 ? tmp15788 : tmp15797;
  assign tmp15780 = s6 ? tmp15781 : tmp15787;
  assign tmp15719 = ~(s7 ? tmp15720 : tmp15780);
  assign tmp15696 = s8 ? tmp15697 : tmp15719;
  assign tmp15806 = s7 ? tmp15720 : tmp15780;
  assign tmp15813 = s0 ? tmp15728 : tmp15758;
  assign tmp15812 = s1 ? tmp15813 : tmp15728;
  assign tmp15811 = s2 ? tmp15812 : tmp15737;
  assign tmp15816 = s0 ? tmp15726 : tmp15728;
  assign tmp15815 = s1 ? tmp15728 : tmp15816;
  assign tmp15814 = s2 ? tmp15739 : tmp15815;
  assign tmp15810 = s3 ? tmp15811 : tmp15814;
  assign tmp15809 = s4 ? tmp15728 : tmp15810;
  assign tmp15822 = s0 ? 1 : tmp15758;
  assign tmp15821 = s1 ? tmp15737 : tmp15822;
  assign tmp15824 = s0 ? 1 : tmp15728;
  assign tmp15823 = s1 ? tmp15824 : tmp15728;
  assign tmp15820 = s2 ? tmp15821 : tmp15823;
  assign tmp15828 = l1 ? 1 : tmp15726;
  assign tmp15829 = ~(l1 ? 1 : tmp15770);
  assign tmp15827 = s0 ? tmp15828 : tmp15829;
  assign tmp15826 = s1 ? tmp15728 : tmp15827;
  assign tmp15830 = s1 ? tmp15751 : tmp15728;
  assign tmp15825 = s2 ? tmp15826 : tmp15830;
  assign tmp15819 = s3 ? tmp15820 : tmp15825;
  assign tmp15835 = ~(l1 ? tmp15409 : tmp15726);
  assign tmp15834 = s0 ? 1 : tmp15835;
  assign tmp15833 = s1 ? tmp15834 : tmp15757;
  assign tmp15836 = ~(s1 ? tmp15760 : tmp15813);
  assign tmp15832 = s2 ? tmp15833 : tmp15836;
  assign tmp15840 = l1 ? 1 : tmp15770;
  assign tmp15839 = s0 ? tmp15840 : tmp15835;
  assign tmp15841 = ~(s0 ? tmp15728 : 0);
  assign tmp15838 = s1 ? tmp15839 : tmp15841;
  assign tmp15837 = s2 ? tmp15838 : 1;
  assign tmp15831 = ~(s3 ? tmp15832 : tmp15837);
  assign tmp15818 = s4 ? tmp15819 : tmp15831;
  assign tmp15846 = s0 ? tmp15840 : 1;
  assign tmp15845 = s1 ? tmp15846 : tmp15776;
  assign tmp15848 = s0 ? tmp15726 : tmp15421;
  assign tmp15847 = ~(s1 ? tmp15848 : tmp15421);
  assign tmp15844 = s2 ? tmp15845 : tmp15847;
  assign tmp15843 = s3 ? tmp15844 : 1;
  assign tmp15852 = s0 ? 1 : tmp15840;
  assign tmp15851 = s1 ? tmp15852 : tmp15424;
  assign tmp15850 = s2 ? tmp15775 : tmp15851;
  assign tmp15849 = s3 ? tmp15850 : tmp15778;
  assign tmp15842 = ~(s4 ? tmp15843 : tmp15849);
  assign tmp15817 = s5 ? tmp15818 : tmp15842;
  assign tmp15808 = s6 ? tmp15809 : tmp15817;
  assign tmp15857 = s1 ? tmp15737 : tmp15728;
  assign tmp15856 = s2 ? tmp15812 : tmp15857;
  assign tmp15858 = s2 ? tmp15786 : tmp15815;
  assign tmp15855 = s3 ? tmp15856 : tmp15858;
  assign tmp15854 = s4 ? tmp15728 : tmp15855;
  assign tmp15863 = s1 ? tmp15737 : tmp15758;
  assign tmp15862 = s2 ? tmp15863 : tmp15728;
  assign tmp15865 = s1 ? tmp15728 : tmp15829;
  assign tmp15864 = s2 ? tmp15865 : tmp15830;
  assign tmp15861 = s3 ? tmp15862 : tmp15864;
  assign tmp15867 = s2 ? tmp15833 : tmp15835;
  assign tmp15866 = ~(s3 ? tmp15867 : tmp15837);
  assign tmp15860 = s4 ? tmp15861 : tmp15866;
  assign tmp15871 = s1 ? tmp15846 : tmp15770;
  assign tmp15870 = s2 ? tmp15871 : tmp15616;
  assign tmp15869 = s3 ? tmp15870 : 1;
  assign tmp15873 = s2 ? tmp15804 : tmp15840;
  assign tmp15872 = s3 ? tmp15873 : 1;
  assign tmp15868 = ~(s4 ? tmp15869 : tmp15872);
  assign tmp15859 = s5 ? tmp15860 : tmp15868;
  assign tmp15853 = s6 ? tmp15854 : tmp15859;
  assign tmp15807 = s7 ? tmp15808 : tmp15853;
  assign tmp15805 = ~(s8 ? tmp15806 : tmp15807);
  assign tmp15695 = s9 ? tmp15696 : tmp15805;
  assign tmp15875 = s8 ? tmp15806 : tmp15720;
  assign tmp15883 = s1 ? tmp15839 : 1;
  assign tmp15882 = s2 ? tmp15883 : 1;
  assign tmp15881 = ~(s3 ? tmp15867 : tmp15882);
  assign tmp15880 = s4 ? tmp15861 : tmp15881;
  assign tmp15879 = s5 ? tmp15880 : tmp15868;
  assign tmp15878 = ~(s6 ? tmp15854 : tmp15879);
  assign tmp15877 = s7 ? tmp15712 : tmp15878;
  assign tmp15889 = s1 ? tmp15724 : 0;
  assign tmp15888 = ~(s2 ? tmp15889 : 0);
  assign tmp15887 = ~(s3 ? tmp15795 : tmp15888);
  assign tmp15886 = s4 ? tmp15789 : tmp15887;
  assign tmp15885 = s5 ? tmp15886 : tmp15797;
  assign tmp15884 = ~(s6 ? tmp15781 : tmp15885);
  assign tmp15876 = ~(s8 ? tmp15877 : tmp15884);
  assign tmp15874 = ~(s9 ? tmp15875 : tmp15876);
  assign tmp15694 = s10 ? tmp15695 : tmp15874;
  assign tmp15894 = ~(s6 ? tmp15854 : tmp15859);
  assign tmp15893 = s7 ? tmp15712 : tmp15894;
  assign tmp15895 = ~(s6 ? tmp15781 : tmp15787);
  assign tmp15892 = ~(s8 ? tmp15893 : tmp15895);
  assign tmp15891 = ~(s9 ? tmp15875 : tmp15892);
  assign tmp15890 = s10 ? tmp15695 : tmp15891;
  assign tmp15693 = s11 ? tmp15694 : tmp15890;
  assign tmp15642 = s12 ? tmp15643 : tmp15693;
  assign tmp15906 = l2 ? tmp15672 : 1;
  assign tmp15905 = l1 ? 1 : tmp15906;
  assign tmp15909 = l2 ? tmp15672 : 0;
  assign tmp15908 = l1 ? 1 : tmp15909;
  assign tmp15907 = s0 ? tmp15908 : tmp15905;
  assign tmp15904 = s1 ? tmp15905 : tmp15907;
  assign tmp15914 = ~(l2 ? tmp15672 : 0);
  assign tmp15913 = ~(l1 ? 1 : tmp15914);
  assign tmp15912 = s0 ? tmp15905 : tmp15913;
  assign tmp15911 = s1 ? tmp15912 : tmp15905;
  assign tmp15910 = s2 ? tmp15905 : tmp15911;
  assign tmp15903 = s3 ? tmp15904 : tmp15910;
  assign tmp15918 = s0 ? tmp15905 : tmp15908;
  assign tmp15917 = s1 ? tmp15918 : tmp15905;
  assign tmp15920 = s0 ? tmp15905 : 1;
  assign tmp15921 = s0 ? tmp15908 : 1;
  assign tmp15919 = s1 ? tmp15920 : tmp15921;
  assign tmp15916 = s2 ? tmp15917 : tmp15919;
  assign tmp15924 = l1 ? 1 : tmp15672;
  assign tmp15923 = s1 ? tmp15924 : 1;
  assign tmp15926 = s0 ? 1 : tmp15905;
  assign tmp15925 = s1 ? tmp15905 : tmp15926;
  assign tmp15922 = s2 ? tmp15923 : tmp15925;
  assign tmp15915 = s3 ? tmp15916 : tmp15922;
  assign tmp15902 = s4 ? tmp15903 : tmp15915;
  assign tmp15933 = l1 ? 1 : tmp15914;
  assign tmp15934 = ~(l1 ? 1 : tmp15906);
  assign tmp15932 = ~(s0 ? tmp15933 : tmp15934);
  assign tmp15931 = s1 ? tmp15912 : tmp15932;
  assign tmp15936 = s0 ? tmp15933 : tmp15934;
  assign tmp15937 = ~(s0 ? tmp15905 : tmp15913);
  assign tmp15935 = ~(s1 ? tmp15936 : tmp15937);
  assign tmp15930 = s2 ? tmp15931 : tmp15935;
  assign tmp15941 = l1 ? 1 : tmp15404;
  assign tmp15940 = s0 ? tmp15905 : tmp15941;
  assign tmp15939 = ~(s1 ? 1 : tmp15940);
  assign tmp15938 = ~(s2 ? tmp15936 : tmp15939);
  assign tmp15929 = s3 ? tmp15930 : tmp15938;
  assign tmp15944 = s1 ? tmp15926 : tmp15468;
  assign tmp15945 = s1 ? tmp15468 : tmp15918;
  assign tmp15943 = s2 ? tmp15944 : tmp15945;
  assign tmp15947 = s1 ? tmp15940 : 1;
  assign tmp15946 = s2 ? tmp15947 : 1;
  assign tmp15942 = s3 ? tmp15943 : tmp15946;
  assign tmp15928 = s4 ? tmp15929 : tmp15942;
  assign tmp15952 = s0 ? tmp15941 : tmp15905;
  assign tmp15951 = s1 ? tmp15926 : tmp15952;
  assign tmp15950 = s2 ? tmp15947 : tmp15951;
  assign tmp15949 = s3 ? tmp15950 : 1;
  assign tmp15955 = s1 ? tmp15952 : tmp15940;
  assign tmp15954 = s2 ? 1 : tmp15955;
  assign tmp15953 = s3 ? tmp15954 : 1;
  assign tmp15948 = s4 ? tmp15949 : tmp15953;
  assign tmp15927 = s5 ? tmp15928 : tmp15948;
  assign tmp15901 = s6 ? tmp15902 : tmp15927;
  assign tmp15960 = s1 ? tmp15920 : tmp15924;
  assign tmp15959 = s2 ? tmp15917 : tmp15960;
  assign tmp15958 = s3 ? tmp15959 : tmp15922;
  assign tmp15957 = s4 ? tmp15903 : tmp15958;
  assign tmp15965 = s1 ? tmp15905 : tmp15912;
  assign tmp15964 = s2 ? tmp15911 : tmp15965;
  assign tmp15967 = s1 ? 1 : tmp15940;
  assign tmp15966 = s2 ? tmp15905 : tmp15967;
  assign tmp15963 = s3 ? tmp15964 : tmp15966;
  assign tmp15969 = s2 ? tmp15944 : tmp15905;
  assign tmp15968 = s3 ? tmp15969 : tmp15946;
  assign tmp15962 = s4 ? tmp15963 : tmp15968;
  assign tmp15973 = s1 ? tmp15905 : 1;
  assign tmp15972 = s2 ? tmp15947 : tmp15973;
  assign tmp15971 = s3 ? tmp15972 : 1;
  assign tmp15975 = s2 ? 1 : tmp15905;
  assign tmp15974 = s3 ? tmp15975 : 1;
  assign tmp15970 = s4 ? tmp15971 : tmp15974;
  assign tmp15961 = s5 ? tmp15962 : tmp15970;
  assign tmp15956 = s6 ? tmp15957 : tmp15961;
  assign tmp15900 = s7 ? tmp15901 : tmp15956;
  assign tmp15985 = ~(l3 ? 1 : 0);
  assign tmp15984 = ~(l1 ? 1 : tmp15985);
  assign tmp15983 = s0 ? tmp15924 : tmp15984;
  assign tmp15982 = s1 ? tmp15983 : tmp15924;
  assign tmp15981 = s2 ? tmp15924 : tmp15982;
  assign tmp15980 = s3 ? tmp15924 : tmp15981;
  assign tmp15988 = s0 ? tmp15924 : 1;
  assign tmp15987 = s2 ? tmp15924 : tmp15988;
  assign tmp15991 = s0 ? tmp15424 : tmp15924;
  assign tmp15990 = s1 ? tmp15924 : tmp15991;
  assign tmp15989 = s2 ? tmp15923 : tmp15990;
  assign tmp15986 = s3 ? tmp15987 : tmp15989;
  assign tmp15979 = s4 ? tmp15980 : tmp15986;
  assign tmp15998 = l1 ? 1 : tmp15985;
  assign tmp15999 = ~(l1 ? 1 : tmp15672);
  assign tmp15997 = ~(s0 ? tmp15998 : tmp15999);
  assign tmp15996 = s1 ? tmp15983 : tmp15997;
  assign tmp16001 = s0 ? tmp15998 : tmp15999;
  assign tmp16002 = ~(s0 ? tmp15924 : tmp15984);
  assign tmp16000 = ~(s1 ? tmp16001 : tmp16002);
  assign tmp15995 = s2 ? tmp15996 : tmp16000;
  assign tmp16005 = s0 ? tmp15924 : tmp15424;
  assign tmp16004 = ~(s1 ? tmp15472 : tmp16005);
  assign tmp16003 = ~(s2 ? tmp16001 : tmp16004);
  assign tmp15994 = s3 ? tmp15995 : tmp16003;
  assign tmp16009 = s0 ? 1 : tmp15924;
  assign tmp16008 = s1 ? tmp16009 : tmp15468;
  assign tmp16010 = s1 ? tmp15468 : tmp15924;
  assign tmp16007 = s2 ? tmp16008 : tmp16010;
  assign tmp16012 = s1 ? tmp16005 : tmp15472;
  assign tmp16011 = s2 ? tmp16012 : 1;
  assign tmp16006 = s3 ? tmp16007 : tmp16011;
  assign tmp15993 = s4 ? tmp15994 : tmp16006;
  assign tmp16016 = s1 ? tmp16005 : tmp15424;
  assign tmp16015 = s2 ? tmp16016 : tmp15991;
  assign tmp16014 = s3 ? tmp16015 : 1;
  assign tmp16019 = s1 ? 1 : tmp15424;
  assign tmp16020 = s1 ? tmp15991 : tmp16005;
  assign tmp16018 = s2 ? tmp16019 : tmp16020;
  assign tmp16021 = s2 ? tmp15616 : 1;
  assign tmp16017 = s3 ? tmp16018 : tmp16021;
  assign tmp16013 = s4 ? tmp16014 : tmp16017;
  assign tmp15992 = s5 ? tmp15993 : tmp16013;
  assign tmp15978 = s6 ? tmp15979 : tmp15992;
  assign tmp16027 = s1 ? tmp15924 : tmp15983;
  assign tmp16026 = s2 ? tmp15982 : tmp16027;
  assign tmp16029 = s1 ? tmp15472 : tmp16005;
  assign tmp16028 = s2 ? tmp15924 : tmp16029;
  assign tmp16025 = s3 ? tmp16026 : tmp16028;
  assign tmp16031 = s2 ? tmp16008 : tmp15924;
  assign tmp16033 = s1 ? tmp16005 : 1;
  assign tmp16032 = s2 ? tmp16033 : 1;
  assign tmp16030 = s3 ? tmp16031 : tmp16032;
  assign tmp16024 = s4 ? tmp16025 : tmp16030;
  assign tmp16036 = s2 ? tmp16016 : tmp15990;
  assign tmp16035 = s3 ? tmp16036 : 1;
  assign tmp16039 = s1 ? tmp15924 : tmp16005;
  assign tmp16038 = s2 ? tmp15424 : tmp16039;
  assign tmp16037 = s3 ? tmp16038 : 1;
  assign tmp16034 = s4 ? tmp16035 : tmp16037;
  assign tmp16023 = s5 ? tmp16024 : tmp16034;
  assign tmp16022 = s6 ? tmp15979 : tmp16023;
  assign tmp15977 = s7 ? tmp15978 : tmp16022;
  assign tmp15976 = s8 ? tmp15900 : tmp15977;
  assign tmp15899 = s9 ? tmp15900 : tmp15976;
  assign tmp16048 = s0 ? tmp15424 : tmp15905;
  assign tmp16047 = s1 ? tmp15905 : tmp16048;
  assign tmp16046 = s2 ? tmp15923 : tmp16047;
  assign tmp16045 = s3 ? tmp15916 : tmp16046;
  assign tmp16044 = s4 ? tmp15903 : tmp16045;
  assign tmp16053 = ~(s1 ? tmp15472 : tmp15940);
  assign tmp16052 = ~(s2 ? tmp15936 : tmp16053);
  assign tmp16051 = s3 ? tmp15930 : tmp16052;
  assign tmp16056 = s1 ? tmp15940 : tmp15472;
  assign tmp16055 = s2 ? tmp16056 : 1;
  assign tmp16054 = s3 ? tmp15943 : tmp16055;
  assign tmp16050 = s4 ? tmp16051 : tmp16054;
  assign tmp16060 = s1 ? tmp15940 : tmp15424;
  assign tmp16061 = s1 ? tmp16048 : tmp15952;
  assign tmp16059 = s2 ? tmp16060 : tmp16061;
  assign tmp16058 = s3 ? tmp16059 : 1;
  assign tmp16063 = s2 ? tmp16019 : tmp15955;
  assign tmp16062 = s3 ? tmp16063 : tmp16021;
  assign tmp16057 = s4 ? tmp16058 : tmp16062;
  assign tmp16049 = s5 ? tmp16050 : tmp16057;
  assign tmp16043 = s6 ? tmp16044 : tmp16049;
  assign tmp16066 = s3 ? tmp15959 : tmp16046;
  assign tmp16065 = s4 ? tmp15903 : tmp16066;
  assign tmp16071 = s1 ? tmp15472 : tmp15940;
  assign tmp16070 = s2 ? tmp15905 : tmp16071;
  assign tmp16069 = s3 ? tmp15964 : tmp16070;
  assign tmp16068 = s4 ? tmp16069 : tmp15968;
  assign tmp16074 = s2 ? tmp16060 : tmp15973;
  assign tmp16073 = s3 ? tmp16074 : 1;
  assign tmp16076 = s2 ? tmp15424 : tmp15905;
  assign tmp16075 = s3 ? tmp16076 : 1;
  assign tmp16072 = s4 ? tmp16073 : tmp16075;
  assign tmp16067 = s5 ? tmp16068 : tmp16072;
  assign tmp16064 = s6 ? tmp16065 : tmp16067;
  assign tmp16042 = s7 ? tmp16043 : tmp16064;
  assign tmp16041 = s8 ? tmp16042 : tmp16043;
  assign tmp16084 = l1 ? 1 : tmp15409;
  assign tmp16083 = s0 ? tmp16084 : 1;
  assign tmp16082 = s1 ? 1 : tmp16083;
  assign tmp16088 = ~(l1 ? 1 : tmp15404);
  assign tmp16087 = s0 ? 1 : tmp16088;
  assign tmp16086 = s1 ? tmp16087 : 1;
  assign tmp16085 = s2 ? 1 : tmp16086;
  assign tmp16081 = s3 ? tmp16082 : tmp16085;
  assign tmp16092 = s0 ? 1 : tmp16084;
  assign tmp16091 = s1 ? tmp16092 : 1;
  assign tmp16090 = s2 ? tmp16091 : 1;
  assign tmp16089 = s3 ? tmp16090 : 1;
  assign tmp16080 = s4 ? tmp16081 : tmp16089;
  assign tmp16097 = s1 ? 1 : tmp16087;
  assign tmp16096 = s2 ? tmp16086 : tmp16097;
  assign tmp16100 = s0 ? 1 : tmp15941;
  assign tmp16099 = s1 ? 1 : tmp16100;
  assign tmp16098 = s2 ? 1 : tmp16099;
  assign tmp16095 = s3 ? tmp16096 : tmp16098;
  assign tmp16103 = s1 ? 1 : tmp15468;
  assign tmp16102 = s2 ? tmp16103 : 1;
  assign tmp16105 = s1 ? tmp16100 : 1;
  assign tmp16104 = s2 ? tmp16105 : 1;
  assign tmp16101 = s3 ? tmp16102 : tmp16104;
  assign tmp16094 = s4 ? tmp16095 : tmp16101;
  assign tmp16107 = s3 ? tmp16104 : 1;
  assign tmp16106 = s4 ? tmp16107 : 1;
  assign tmp16093 = s5 ? tmp16094 : tmp16106;
  assign tmp16079 = s6 ? tmp16080 : tmp16093;
  assign tmp16112 = s2 ? tmp15424 : tmp15924;
  assign tmp16111 = s3 ? tmp16112 : 1;
  assign tmp16110 = s4 ? tmp16035 : tmp16111;
  assign tmp16109 = s5 ? tmp16024 : tmp16110;
  assign tmp16108 = s6 ? tmp15979 : tmp16109;
  assign tmp16078 = s7 ? tmp16079 : tmp16108;
  assign tmp16077 = s8 ? tmp16078 : tmp16064;
  assign tmp16040 = s9 ? tmp16041 : tmp16077;
  assign tmp15898 = s10 ? tmp15899 : tmp16040;
  assign tmp16116 = s7 ? tmp16079 : tmp16022;
  assign tmp16115 = s8 ? tmp16116 : tmp16064;
  assign tmp16114 = s9 ? tmp16041 : tmp16115;
  assign tmp16113 = s10 ? tmp15899 : tmp16114;
  assign tmp15897 = s11 ? tmp15898 : tmp16113;
  assign tmp15896 = s12 ? tmp15897 : 1;
  assign tmp15641 = s13 ? tmp15642 : tmp15896;
  assign tmp15390 = s14 ? tmp15391 : tmp15641;
  assign tmp16126 = s4 ? 1 : tmp15465;
  assign tmp16132 = s0 ? tmp15941 : 1;
  assign tmp16131 = s1 ? tmp16132 : 1;
  assign tmp16130 = s2 ? tmp16105 : tmp16131;
  assign tmp16129 = s3 ? tmp16130 : 1;
  assign tmp16135 = s1 ? 1 : tmp15472;
  assign tmp16136 = s1 ? tmp15472 : tmp15468;
  assign tmp16134 = s2 ? tmp16135 : tmp16136;
  assign tmp16133 = s3 ? tmp16134 : 1;
  assign tmp16128 = s4 ? tmp16129 : tmp16133;
  assign tmp16127 = s5 ? tmp16128 : 1;
  assign tmp16125 = s6 ? tmp16126 : tmp16127;
  assign tmp16141 = s2 ? tmp16135 : 1;
  assign tmp16140 = s3 ? tmp16141 : 1;
  assign tmp16139 = s4 ? tmp16107 : tmp16140;
  assign tmp16138 = s5 ? tmp16139 : 1;
  assign tmp16137 = s6 ? tmp16126 : tmp16138;
  assign tmp16124 = s7 ? tmp16125 : tmp16137;
  assign tmp16147 = ~(l2 ? tmp15726 : 0);
  assign tmp16146 = l1 ? 1 : tmp16147;
  assign tmp16150 = s0 ? 1 : tmp16146;
  assign tmp16149 = s1 ? tmp16150 : tmp16146;
  assign tmp16148 = s2 ? tmp16149 : tmp16146;
  assign tmp16145 = s3 ? tmp16146 : tmp16148;
  assign tmp16154 = s0 ? tmp16146 : 0;
  assign tmp16153 = s1 ? tmp16154 : tmp16146;
  assign tmp16155 = s0 ? tmp16146 : 1;
  assign tmp16152 = s2 ? tmp16153 : tmp16155;
  assign tmp16157 = s1 ? tmp15726 : 0;
  assign tmp16158 = ~(l1 ? 1 : tmp16147);
  assign tmp16156 = ~(s2 ? tmp16157 : tmp16158);
  assign tmp16151 = s3 ? tmp16152 : tmp16156;
  assign tmp16144 = s4 ? tmp16145 : tmp16151;
  assign tmp16164 = s0 ? tmp16146 : tmp15941;
  assign tmp16163 = s1 ? tmp16164 : 1;
  assign tmp16166 = s0 ? tmp15941 : tmp16146;
  assign tmp16165 = s1 ? tmp16166 : tmp16146;
  assign tmp16162 = s2 ? tmp16163 : tmp16165;
  assign tmp16168 = s1 ? tmp15846 : tmp16146;
  assign tmp16167 = s2 ? tmp16146 : tmp16168;
  assign tmp16161 = s3 ? tmp16162 : tmp16167;
  assign tmp16172 = ~(s0 ? 1 : tmp15726);
  assign tmp16171 = s1 ? tmp16150 : tmp16172;
  assign tmp16174 = s0 ? 1 : tmp15726;
  assign tmp16175 = ~(s0 ? tmp16146 : 0);
  assign tmp16173 = ~(s1 ? tmp16174 : tmp16175);
  assign tmp16170 = s2 ? tmp16171 : tmp16173;
  assign tmp16178 = ~(s0 ? tmp15726 : 0);
  assign tmp16177 = s1 ? tmp16146 : tmp16178;
  assign tmp16176 = s2 ? tmp16177 : 1;
  assign tmp16169 = s3 ? tmp16170 : tmp16176;
  assign tmp16160 = s4 ? tmp16161 : tmp16169;
  assign tmp16182 = s1 ? tmp16155 : tmp15852;
  assign tmp16183 = s1 ? tmp15846 : 1;
  assign tmp16181 = s2 ? tmp16182 : tmp16183;
  assign tmp16180 = s3 ? tmp16181 : 1;
  assign tmp16186 = s1 ? 1 : tmp15852;
  assign tmp16187 = s1 ? tmp16150 : 1;
  assign tmp16185 = s2 ? tmp16186 : tmp16187;
  assign tmp16188 = s2 ? tmp16183 : 1;
  assign tmp16184 = s3 ? tmp16185 : tmp16188;
  assign tmp16179 = s4 ? tmp16180 : tmp16184;
  assign tmp16159 = s5 ? tmp16160 : tmp16179;
  assign tmp16143 = s6 ? tmp16144 : tmp16159;
  assign tmp16193 = s2 ? tmp16163 : tmp16146;
  assign tmp16192 = s3 ? tmp16193 : tmp16167;
  assign tmp16195 = s2 ? tmp16171 : tmp16146;
  assign tmp16197 = s1 ? tmp16146 : 1;
  assign tmp16196 = s2 ? tmp16197 : 1;
  assign tmp16194 = s3 ? tmp16195 : tmp16196;
  assign tmp16191 = s4 ? tmp16192 : tmp16194;
  assign tmp16201 = s1 ? tmp16155 : tmp15840;
  assign tmp16200 = s2 ? tmp16201 : tmp16183;
  assign tmp16199 = s3 ? tmp16200 : 1;
  assign tmp16204 = s1 ? 1 : tmp15840;
  assign tmp16203 = s2 ? tmp16204 : tmp16146;
  assign tmp16202 = s3 ? tmp16203 : tmp16183;
  assign tmp16198 = s4 ? tmp16199 : tmp16202;
  assign tmp16190 = s5 ? tmp16191 : tmp16198;
  assign tmp16189 = s6 ? tmp16144 : tmp16190;
  assign tmp16142 = s7 ? tmp16143 : tmp16189;
  assign tmp16123 = s8 ? tmp16124 : tmp16142;
  assign tmp16211 = s1 ? tmp16164 : tmp16146;
  assign tmp16210 = s2 ? tmp16211 : tmp16155;
  assign tmp16209 = s3 ? tmp16210 : tmp16156;
  assign tmp16208 = s4 ? tmp16145 : tmp16209;
  assign tmp16217 = ~(s0 ? tmp16146 : tmp15941);
  assign tmp16216 = ~(s1 ? tmp16174 : tmp16217);
  assign tmp16215 = s2 ? tmp16171 : tmp16216;
  assign tmp16214 = s3 ? tmp16215 : tmp16176;
  assign tmp16213 = s4 ? tmp16161 : tmp16214;
  assign tmp16212 = s5 ? tmp16213 : tmp16179;
  assign tmp16207 = s6 ? tmp16208 : tmp16212;
  assign tmp16218 = s6 ? tmp16208 : tmp16190;
  assign tmp16206 = s7 ? tmp16207 : tmp16218;
  assign tmp16225 = s0 ? tmp15840 : tmp15424;
  assign tmp16224 = s1 ? tmp16225 : tmp15840;
  assign tmp16223 = s2 ? tmp16224 : tmp15846;
  assign tmp16226 = ~(s2 ? tmp16157 : tmp15829);
  assign tmp16222 = s3 ? tmp16223 : tmp16226;
  assign tmp16221 = s4 ? tmp15840 : tmp16222;
  assign tmp16231 = s1 ? tmp16225 : tmp15424;
  assign tmp16233 = s0 ? tmp15424 : tmp15840;
  assign tmp16232 = s1 ? tmp16233 : tmp15840;
  assign tmp16230 = s2 ? tmp16231 : tmp16232;
  assign tmp16235 = s1 ? tmp15846 : tmp15840;
  assign tmp16234 = s2 ? tmp15840 : tmp16235;
  assign tmp16229 = s3 ? tmp16230 : tmp16234;
  assign tmp16238 = s1 ? tmp15852 : tmp16172;
  assign tmp16240 = ~(s0 ? tmp15840 : tmp15424);
  assign tmp16239 = ~(s1 ? tmp16174 : tmp16240);
  assign tmp16237 = s2 ? tmp16238 : tmp16239;
  assign tmp16242 = s1 ? tmp15840 : tmp16178;
  assign tmp16241 = s2 ? tmp16242 : 1;
  assign tmp16236 = s3 ? tmp16237 : tmp16241;
  assign tmp16228 = s4 ? tmp16229 : tmp16236;
  assign tmp16246 = s1 ? tmp15846 : tmp15852;
  assign tmp16247 = s1 ? tmp15840 : tmp15468;
  assign tmp16245 = s2 ? tmp16246 : tmp16247;
  assign tmp16244 = s3 ? tmp16245 : 1;
  assign tmp16250 = s1 ? tmp15852 : tmp15472;
  assign tmp16249 = s2 ? tmp16186 : tmp16250;
  assign tmp16248 = s3 ? tmp16249 : tmp16188;
  assign tmp16243 = s4 ? tmp16244 : tmp16248;
  assign tmp16227 = s5 ? tmp16228 : tmp16243;
  assign tmp16220 = s6 ? tmp16221 : tmp16227;
  assign tmp16255 = s2 ? tmp16231 : tmp15840;
  assign tmp16254 = s3 ? tmp16255 : tmp16234;
  assign tmp16257 = s2 ? tmp16238 : tmp15840;
  assign tmp16259 = s1 ? tmp15840 : 1;
  assign tmp16258 = s2 ? tmp16259 : 1;
  assign tmp16256 = s3 ? tmp16257 : tmp16258;
  assign tmp16253 = s4 ? tmp16254 : tmp16256;
  assign tmp16262 = s2 ? tmp16235 : tmp16259;
  assign tmp16261 = s3 ? tmp16262 : 1;
  assign tmp16264 = s2 ? tmp16204 : tmp15840;
  assign tmp16263 = s3 ? tmp16264 : tmp16183;
  assign tmp16260 = s4 ? tmp16261 : tmp16263;
  assign tmp16252 = s5 ? tmp16253 : tmp16260;
  assign tmp16251 = s6 ? tmp16221 : tmp16252;
  assign tmp16219 = s7 ? tmp16220 : tmp16251;
  assign tmp16205 = s8 ? tmp16206 : tmp16219;
  assign tmp16122 = s9 ? tmp16123 : tmp16205;
  assign tmp16269 = s4 ? tmp16146 : tmp16209;
  assign tmp16274 = s1 ? tmp16164 : tmp15941;
  assign tmp16273 = s2 ? tmp16274 : tmp16165;
  assign tmp16272 = s3 ? tmp16273 : tmp16167;
  assign tmp16271 = s4 ? tmp16272 : tmp16214;
  assign tmp16278 = s1 ? tmp16146 : tmp16100;
  assign tmp16277 = s2 ? tmp16182 : tmp16278;
  assign tmp16276 = s3 ? tmp16277 : 1;
  assign tmp16281 = s1 ? tmp16150 : tmp16132;
  assign tmp16280 = s2 ? tmp16186 : tmp16281;
  assign tmp16279 = s3 ? tmp16280 : tmp16188;
  assign tmp16275 = s4 ? tmp16276 : tmp16279;
  assign tmp16270 = s5 ? tmp16271 : tmp16275;
  assign tmp16268 = s6 ? tmp16269 : tmp16270;
  assign tmp16286 = s2 ? tmp16274 : tmp16146;
  assign tmp16285 = s3 ? tmp16286 : tmp16167;
  assign tmp16284 = s4 ? tmp16285 : tmp16194;
  assign tmp16289 = s2 ? tmp16201 : tmp16197;
  assign tmp16288 = s3 ? tmp16289 : 1;
  assign tmp16287 = s4 ? tmp16288 : tmp16202;
  assign tmp16283 = s5 ? tmp16284 : tmp16287;
  assign tmp16282 = s6 ? tmp16269 : tmp16283;
  assign tmp16267 = s7 ? tmp16268 : tmp16282;
  assign tmp16266 = s8 ? tmp16267 : tmp16268;
  assign tmp16295 = s3 ? tmp16264 : 1;
  assign tmp16294 = s4 ? tmp16261 : tmp16295;
  assign tmp16293 = s5 ? tmp16253 : tmp16294;
  assign tmp16292 = s6 ? tmp16221 : tmp16293;
  assign tmp16291 = s7 ? tmp16137 : tmp16292;
  assign tmp16299 = s3 ? tmp16203 : 1;
  assign tmp16298 = s4 ? tmp16288 : tmp16299;
  assign tmp16297 = s5 ? tmp16284 : tmp16298;
  assign tmp16296 = s6 ? tmp16269 : tmp16297;
  assign tmp16290 = s8 ? tmp16291 : tmp16296;
  assign tmp16265 = s9 ? tmp16266 : tmp16290;
  assign tmp16121 = s10 ? tmp16122 : tmp16265;
  assign tmp16303 = s7 ? tmp16137 : tmp16251;
  assign tmp16302 = s8 ? tmp16303 : tmp16282;
  assign tmp16301 = s9 ? tmp16266 : tmp16302;
  assign tmp16300 = s10 ? tmp16122 : tmp16301;
  assign tmp16120 = s11 ? tmp16121 : tmp16300;
  assign tmp16119 = s12 ? 1 : tmp16120;
  assign tmp16118 = s13 ? tmp16119 : 1;
  assign tmp16117 = s14 ? 1 : tmp16118;
  assign tmp15389 = s15 ? tmp15390 : tmp16117;
  assign tmp15388 = s16 ? 1 : tmp15389;
  assign tmp16315 = s4 ? tmp15465 : tmp15469;
  assign tmp16314 = s5 ? 1 : tmp16315;
  assign tmp16313 = s6 ? 1 : tmp16314;
  assign tmp16318 = s4 ? tmp15465 : 1;
  assign tmp16317 = s5 ? 1 : tmp16318;
  assign tmp16316 = s6 ? 1 : tmp16317;
  assign tmp16312 = s7 ? tmp16313 : tmp16316;
  assign tmp16311 = s8 ? tmp15413 : tmp16312;
  assign tmp16310 = s9 ? tmp15395 : tmp16311;
  assign tmp16320 = s8 ? tmp15396 : tmp15397;
  assign tmp16322 = s7 ? tmp15410 : tmp16316;
  assign tmp16323 = s7 ? tmp15523 : tmp15410;
  assign tmp16321 = s8 ? tmp16322 : tmp16323;
  assign tmp16319 = s9 ? tmp16320 : tmp16321;
  assign tmp16309 = s10 ? tmp16310 : tmp16319;
  assign tmp16327 = s7 ? tmp15425 : tmp15410;
  assign tmp16326 = s8 ? tmp16322 : tmp16327;
  assign tmp16325 = s9 ? tmp16320 : tmp16326;
  assign tmp16324 = s10 ? tmp16310 : tmp16325;
  assign tmp16308 = s11 ? tmp16309 : tmp16324;
  assign tmp16333 = s7 ? tmp15540 : tmp15622;
  assign tmp16332 = s8 ? tmp15565 : tmp16333;
  assign tmp16331 = s9 ? tmp15538 : tmp16332;
  assign tmp16335 = s8 ? tmp16333 : tmp15540;
  assign tmp16337 = s7 ? tmp15632 : tmp15622;
  assign tmp16336 = s8 ? tmp15622 : tmp16337;
  assign tmp16334 = s9 ? tmp16335 : tmp16336;
  assign tmp16330 = s10 ? tmp16331 : tmp16334;
  assign tmp16341 = s7 ? tmp15575 : tmp15622;
  assign tmp16340 = s8 ? tmp15557 : tmp16341;
  assign tmp16339 = s9 ? tmp16335 : tmp16340;
  assign tmp16338 = s10 ? tmp16331 : tmp16339;
  assign tmp16329 = s11 ? tmp16330 : tmp16338;
  assign tmp16328 = s12 ? 1 : tmp16329;
  assign tmp16307 = s13 ? tmp16308 : tmp16328;
  assign tmp16347 = ~(s8 ? tmp15679 : 0);
  assign tmp16346 = s9 ? tmp15646 : tmp16347;
  assign tmp16351 = s6 ? tmp15424 : tmp15683;
  assign tmp16350 = ~(s7 ? tmp16351 : 0);
  assign tmp16349 = s8 ? 1 : tmp16350;
  assign tmp16348 = s9 ? 1 : tmp16349;
  assign tmp16345 = s10 ? tmp16346 : tmp16348;
  assign tmp16355 = ~(s7 ? tmp15662 : 0);
  assign tmp16354 = s8 ? 1 : tmp16355;
  assign tmp16353 = s9 ? 1 : tmp16354;
  assign tmp16352 = s10 ? tmp16346 : tmp16353;
  assign tmp16344 = s11 ? tmp16345 : tmp16352;
  assign tmp16360 = ~(s7 ? tmp15698 : tmp15712);
  assign tmp16359 = ~(s8 ? tmp15806 : tmp16360);
  assign tmp16358 = s9 ? tmp15696 : tmp16359;
  assign tmp16362 = s8 ? tmp15697 : tmp15698;
  assign tmp16365 = s6 ? tmp15781 : tmp15885;
  assign tmp16366 = ~(s6 ? tmp15713 : tmp15715);
  assign tmp16364 = ~(s7 ? tmp16365 : tmp16366);
  assign tmp16363 = s8 ? tmp15712 : tmp16364;
  assign tmp16361 = s9 ? tmp16362 : tmp16363;
  assign tmp16357 = s10 ? tmp16358 : tmp16361;
  assign tmp16370 = ~(s7 ? tmp15780 : tmp16366);
  assign tmp16369 = s8 ? tmp15712 : tmp16370;
  assign tmp16368 = s9 ? tmp16362 : tmp16369;
  assign tmp16367 = s10 ? tmp16358 : tmp16368;
  assign tmp16356 = s11 ? tmp16357 : tmp16367;
  assign tmp16343 = s12 ? tmp16344 : tmp16356;
  assign tmp16382 = ~(s1 ? 1 : tmp15920);
  assign tmp16381 = ~(s2 ? tmp15936 : tmp16382);
  assign tmp16380 = s3 ? tmp15930 : tmp16381;
  assign tmp16385 = s1 ? tmp15926 : 1;
  assign tmp16386 = s1 ? 1 : tmp15918;
  assign tmp16384 = s2 ? tmp16385 : tmp16386;
  assign tmp16388 = s1 ? tmp15920 : 1;
  assign tmp16387 = s2 ? tmp16388 : 1;
  assign tmp16383 = s3 ? tmp16384 : tmp16387;
  assign tmp16379 = s4 ? tmp16380 : tmp16383;
  assign tmp16393 = s0 ? tmp15905 : tmp15424;
  assign tmp16392 = s1 ? tmp16393 : 1;
  assign tmp16391 = s2 ? tmp16392 : tmp15926;
  assign tmp16390 = s3 ? tmp16391 : 1;
  assign tmp16396 = s1 ? tmp16048 : tmp15920;
  assign tmp16395 = s2 ? 1 : tmp16396;
  assign tmp16394 = s3 ? tmp16395 : 1;
  assign tmp16389 = s4 ? tmp16390 : tmp16394;
  assign tmp16378 = s5 ? tmp16379 : tmp16389;
  assign tmp16377 = s6 ? tmp15902 : tmp16378;
  assign tmp16402 = s1 ? 1 : tmp15920;
  assign tmp16401 = s2 ? tmp15905 : tmp16402;
  assign tmp16400 = s3 ? tmp15964 : tmp16401;
  assign tmp16404 = s2 ? tmp16385 : tmp15905;
  assign tmp16403 = s3 ? tmp16404 : tmp16387;
  assign tmp16399 = s4 ? tmp16400 : tmp16403;
  assign tmp16408 = s1 ? tmp15905 : tmp15920;
  assign tmp16407 = s2 ? 1 : tmp16408;
  assign tmp16406 = s3 ? tmp16407 : 1;
  assign tmp16405 = s4 ? tmp16390 : tmp16406;
  assign tmp16398 = s5 ? tmp16399 : tmp16405;
  assign tmp16397 = s6 ? tmp15957 : tmp16398;
  assign tmp16376 = s7 ? tmp16377 : tmp16397;
  assign tmp16411 = s5 ? tmp15928 : tmp16389;
  assign tmp16410 = s6 ? tmp15902 : tmp16411;
  assign tmp16413 = s5 ? tmp15962 : tmp16405;
  assign tmp16412 = s6 ? tmp15957 : tmp16413;
  assign tmp16409 = s7 ? tmp16410 : tmp16412;
  assign tmp16375 = s8 ? tmp16376 : tmp16409;
  assign tmp16420 = s1 ? tmp15420 : 1;
  assign tmp16419 = s2 ? 1 : tmp16420;
  assign tmp16418 = s3 ? 1 : tmp16419;
  assign tmp16417 = s4 ? tmp16418 : 1;
  assign tmp16426 = ~(s0 ? tmp15424 : 0);
  assign tmp16425 = s1 ? tmp15420 : tmp16426;
  assign tmp16427 = ~(s1 ? tmp15423 : tmp15654);
  assign tmp16424 = s2 ? tmp16425 : tmp16427;
  assign tmp16429 = ~(s1 ? 1 : tmp16100);
  assign tmp16428 = ~(s2 ? tmp15423 : tmp16429);
  assign tmp16423 = s3 ? tmp16424 : tmp16428;
  assign tmp16430 = s3 ? 1 : tmp16104;
  assign tmp16422 = s4 ? tmp16423 : tmp16430;
  assign tmp16434 = s1 ? 1 : tmp16132;
  assign tmp16433 = s2 ? tmp15467 : tmp16434;
  assign tmp16432 = s3 ? tmp16433 : 1;
  assign tmp16437 = s1 ? tmp15472 : tmp16100;
  assign tmp16436 = s2 ? 1 : tmp16437;
  assign tmp16435 = s3 ? tmp16436 : 1;
  assign tmp16431 = s4 ? tmp16432 : tmp16435;
  assign tmp16421 = s5 ? tmp16422 : tmp16431;
  assign tmp16416 = s6 ? tmp16417 : tmp16421;
  assign tmp16442 = s2 ? tmp16420 : tmp15419;
  assign tmp16441 = s3 ? tmp16442 : tmp16098;
  assign tmp16440 = s4 ? tmp16441 : tmp16430;
  assign tmp16446 = s1 ? 1 : tmp15941;
  assign tmp16445 = s2 ? 1 : tmp16446;
  assign tmp16444 = s3 ? tmp16445 : 1;
  assign tmp16443 = s4 ? tmp15465 : tmp16444;
  assign tmp16439 = s5 ? tmp16440 : tmp16443;
  assign tmp16438 = s6 ? tmp16417 : tmp16439;
  assign tmp16415 = s7 ? tmp16416 : tmp16438;
  assign tmp16414 = s8 ? tmp16409 : tmp16415;
  assign tmp16374 = s9 ? tmp16375 : tmp16414;
  assign tmp16453 = s2 ? tmp16091 : tmp16082;
  assign tmp16452 = s3 ? tmp16453 : 1;
  assign tmp16451 = s4 ? tmp16081 : tmp16452;
  assign tmp16459 = ~(s0 ? tmp15941 : 0);
  assign tmp16458 = s1 ? tmp16087 : tmp16459;
  assign tmp16461 = s0 ? tmp15941 : 0;
  assign tmp16462 = ~(s0 ? 1 : tmp16088);
  assign tmp16460 = ~(s1 ? tmp16461 : tmp16462);
  assign tmp16457 = s2 ? tmp16458 : tmp16460;
  assign tmp16463 = ~(s2 ? tmp16461 : 0);
  assign tmp16456 = s3 ? tmp16457 : tmp16463;
  assign tmp16466 = s1 ? 1 : tmp16092;
  assign tmp16465 = s2 ? 1 : tmp16466;
  assign tmp16464 = s3 ? tmp16465 : 1;
  assign tmp16455 = s4 ? tmp16456 : tmp16464;
  assign tmp16454 = s5 ? tmp16455 : tmp16315;
  assign tmp16450 = s6 ? tmp16451 : tmp16454;
  assign tmp16470 = s3 ? tmp16096 : 1;
  assign tmp16469 = s4 ? tmp16470 : 1;
  assign tmp16468 = s5 ? tmp16469 : tmp16318;
  assign tmp16467 = s6 ? tmp16080 : tmp16468;
  assign tmp16449 = s7 ? tmp16450 : tmp16467;
  assign tmp16448 = s8 ? tmp16449 : tmp16450;
  assign tmp16475 = s4 ? tmp16390 : tmp15974;
  assign tmp16474 = s5 ? tmp16399 : tmp16475;
  assign tmp16473 = s6 ? tmp15957 : tmp16474;
  assign tmp16481 = s0 ? tmp16084 : tmp16088;
  assign tmp16480 = s1 ? tmp16481 : tmp16084;
  assign tmp16479 = s2 ? tmp16084 : tmp16480;
  assign tmp16478 = s3 ? tmp16084 : tmp16479;
  assign tmp16484 = s1 ? tmp16083 : 1;
  assign tmp16483 = s2 ? tmp16084 : tmp16484;
  assign tmp16486 = s1 ? tmp16084 : tmp16092;
  assign tmp16485 = s2 ? 1 : tmp16486;
  assign tmp16482 = s3 ? tmp16483 : tmp16485;
  assign tmp16477 = s4 ? tmp16478 : tmp16482;
  assign tmp16491 = s1 ? tmp16084 : tmp16481;
  assign tmp16490 = s2 ? tmp16480 : tmp16491;
  assign tmp16494 = s0 ? tmp16084 : tmp15941;
  assign tmp16493 = s1 ? 1 : tmp16494;
  assign tmp16492 = s2 ? tmp16084 : tmp16493;
  assign tmp16489 = s3 ? tmp16490 : tmp16492;
  assign tmp16496 = s2 ? tmp16091 : tmp16084;
  assign tmp16498 = s1 ? tmp16494 : 1;
  assign tmp16497 = s2 ? tmp16498 : 1;
  assign tmp16495 = s3 ? tmp16496 : tmp16497;
  assign tmp16488 = s4 ? tmp16489 : tmp16495;
  assign tmp16503 = s0 ? tmp16084 : tmp15424;
  assign tmp16502 = s1 ? tmp16503 : 1;
  assign tmp16504 = s1 ? tmp16084 : 1;
  assign tmp16501 = s2 ? tmp16502 : tmp16504;
  assign tmp16505 = s2 ? tmp16131 : 1;
  assign tmp16500 = s3 ? tmp16501 : tmp16505;
  assign tmp16507 = s2 ? 1 : tmp16084;
  assign tmp16506 = s3 ? tmp16507 : 1;
  assign tmp16499 = s4 ? tmp16500 : tmp16506;
  assign tmp16487 = s5 ? tmp16488 : tmp16499;
  assign tmp16476 = s6 ? tmp16477 : tmp16487;
  assign tmp16472 = s7 ? tmp16473 : tmp16476;
  assign tmp16510 = s5 ? tmp15962 : tmp16475;
  assign tmp16509 = s6 ? tmp15957 : tmp16510;
  assign tmp16508 = s7 ? tmp16509 : tmp16467;
  assign tmp16471 = s8 ? tmp16472 : tmp16508;
  assign tmp16447 = s9 ? tmp16448 : tmp16471;
  assign tmp16373 = s10 ? tmp16374 : tmp16447;
  assign tmp16520 = s1 ? tmp16084 : tmp15941;
  assign tmp16519 = s2 ? 1 : tmp16520;
  assign tmp16518 = s3 ? tmp16519 : 1;
  assign tmp16517 = s4 ? tmp16500 : tmp16518;
  assign tmp16516 = s5 ? tmp16488 : tmp16517;
  assign tmp16515 = s6 ? tmp16477 : tmp16516;
  assign tmp16514 = s7 ? tmp16397 : tmp16515;
  assign tmp16521 = s7 ? tmp16412 : tmp16467;
  assign tmp16513 = s8 ? tmp16514 : tmp16521;
  assign tmp16512 = s9 ? tmp16448 : tmp16513;
  assign tmp16511 = s10 ? tmp16374 : tmp16512;
  assign tmp16372 = s11 ? tmp16373 : tmp16511;
  assign tmp16371 = s12 ? tmp16372 : 1;
  assign tmp16342 = s13 ? tmp16343 : tmp16371;
  assign tmp16306 = s14 ? tmp16307 : tmp16342;
  assign tmp16534 = s2 ? tmp15467 : tmp15471;
  assign tmp16533 = s3 ? tmp16534 : 1;
  assign tmp16532 = s4 ? tmp16533 : tmp16133;
  assign tmp16531 = s5 ? tmp16532 : 1;
  assign tmp16530 = s6 ? tmp16126 : tmp16531;
  assign tmp16537 = s4 ? tmp15465 : tmp16140;
  assign tmp16536 = s5 ? tmp16537 : 1;
  assign tmp16535 = s6 ? tmp16126 : tmp16536;
  assign tmp16529 = s7 ? tmp16530 : tmp16535;
  assign tmp16528 = s8 ? tmp16206 : tmp16529;
  assign tmp16527 = s9 ? tmp16123 : tmp16528;
  assign tmp16542 = s4 ? 1 : tmp16107;
  assign tmp16546 = s2 ? tmp16135 : tmp16437;
  assign tmp16545 = s3 ? tmp16546 : 1;
  assign tmp16544 = s4 ? tmp16129 : tmp16545;
  assign tmp16543 = s5 ? tmp16544 : 1;
  assign tmp16541 = s6 ? tmp16542 : tmp16543;
  assign tmp16547 = s6 ? tmp16542 : tmp16138;
  assign tmp16540 = s7 ? tmp16541 : tmp16547;
  assign tmp16539 = s8 ? tmp16540 : tmp16541;
  assign tmp16549 = s7 ? tmp16137 : tmp16535;
  assign tmp16553 = s4 ? tmp16199 : tmp16299;
  assign tmp16552 = s5 ? tmp16191 : tmp16553;
  assign tmp16551 = s6 ? tmp16208 : tmp16552;
  assign tmp16550 = s7 ? tmp16551 : tmp16547;
  assign tmp16548 = s8 ? tmp16549 : tmp16550;
  assign tmp16538 = s9 ? tmp16539 : tmp16548;
  assign tmp16526 = s10 ? tmp16527 : tmp16538;
  assign tmp16557 = s7 ? tmp16218 : tmp16547;
  assign tmp16556 = s8 ? tmp16549 : tmp16557;
  assign tmp16555 = s9 ? tmp16539 : tmp16556;
  assign tmp16554 = s10 ? tmp16527 : tmp16555;
  assign tmp16525 = s11 ? tmp16526 : tmp16554;
  assign tmp16524 = s12 ? 1 : tmp16525;
  assign tmp16523 = s13 ? tmp16524 : 1;
  assign tmp16522 = s14 ? 1 : tmp16523;
  assign tmp16305 = s15 ? tmp16306 : tmp16522;
  assign tmp16572 = ~(s1 ? tmp15472 : tmp15920);
  assign tmp16571 = ~(s2 ? tmp15936 : tmp16572);
  assign tmp16570 = s3 ? tmp15930 : tmp16571;
  assign tmp16569 = s4 ? tmp16570 : tmp16383;
  assign tmp16576 = s1 ? tmp16393 : tmp15424;
  assign tmp16575 = s2 ? tmp16576 : tmp15926;
  assign tmp16574 = s3 ? tmp16575 : 1;
  assign tmp16578 = s2 ? tmp16446 : tmp16396;
  assign tmp16577 = s3 ? tmp16578 : tmp16021;
  assign tmp16573 = s4 ? tmp16574 : tmp16577;
  assign tmp16568 = s5 ? tmp16569 : tmp16573;
  assign tmp16567 = s6 ? tmp16044 : tmp16568;
  assign tmp16584 = s1 ? tmp15472 : tmp15920;
  assign tmp16583 = s2 ? tmp15905 : tmp16584;
  assign tmp16582 = s3 ? tmp15964 : tmp16583;
  assign tmp16581 = s4 ? tmp16582 : tmp16403;
  assign tmp16587 = s2 ? tmp15424 : tmp16408;
  assign tmp16586 = s3 ? tmp16587 : 1;
  assign tmp16585 = s4 ? tmp16574 : tmp16586;
  assign tmp16580 = s5 ? tmp16581 : tmp16585;
  assign tmp16579 = s6 ? tmp16065 : tmp16580;
  assign tmp16566 = s7 ? tmp16567 : tmp16579;
  assign tmp16594 = s1 ? tmp16048 : tmp15926;
  assign tmp16593 = s2 ? tmp16576 : tmp16594;
  assign tmp16592 = s3 ? tmp16593 : 1;
  assign tmp16596 = s2 ? tmp16019 : tmp16396;
  assign tmp16595 = s3 ? tmp16596 : tmp16021;
  assign tmp16591 = s4 ? tmp16592 : tmp16595;
  assign tmp16590 = s5 ? tmp16050 : tmp16591;
  assign tmp16589 = s6 ? tmp16044 : tmp16590;
  assign tmp16598 = s5 ? tmp16068 : tmp16585;
  assign tmp16597 = s6 ? tmp16065 : tmp16598;
  assign tmp16588 = s7 ? tmp16589 : tmp16597;
  assign tmp16565 = s8 ? tmp16566 : tmp16588;
  assign tmp16607 = s0 ? tmp15941 : tmp15924;
  assign tmp16606 = s1 ? tmp15991 : tmp16607;
  assign tmp16605 = s2 ? tmp16016 : tmp16606;
  assign tmp16604 = s3 ? tmp16605 : 1;
  assign tmp16611 = s0 ? tmp15924 : tmp15941;
  assign tmp16610 = s1 ? tmp15991 : tmp16611;
  assign tmp16609 = s2 ? tmp16019 : tmp16610;
  assign tmp16608 = s3 ? tmp16609 : tmp16021;
  assign tmp16603 = s4 ? tmp16604 : tmp16608;
  assign tmp16602 = s5 ? tmp15993 : tmp16603;
  assign tmp16601 = s6 ? tmp15979 : tmp16602;
  assign tmp16617 = s1 ? tmp15924 : tmp16607;
  assign tmp16616 = s2 ? tmp16016 : tmp16617;
  assign tmp16615 = s3 ? tmp16616 : tmp16505;
  assign tmp16620 = s1 ? tmp15924 : tmp16611;
  assign tmp16619 = s2 ? tmp15424 : tmp16620;
  assign tmp16618 = s3 ? tmp16619 : 1;
  assign tmp16614 = s4 ? tmp16615 : tmp16618;
  assign tmp16613 = s5 ? tmp16024 : tmp16614;
  assign tmp16612 = s6 ? tmp15979 : tmp16613;
  assign tmp16600 = s7 ? tmp16601 : tmp16612;
  assign tmp16599 = s8 ? tmp16588 : tmp16600;
  assign tmp16564 = s9 ? tmp16565 : tmp16599;
  assign tmp16622 = s8 ? tmp16588 : tmp16589;
  assign tmp16627 = s4 ? tmp16574 : tmp16075;
  assign tmp16626 = s5 ? tmp16581 : tmp16627;
  assign tmp16625 = s6 ? tmp16065 : tmp16626;
  assign tmp16633 = s0 ? tmp15908 : tmp15913;
  assign tmp16632 = s1 ? tmp16633 : tmp15908;
  assign tmp16631 = s2 ? tmp15908 : tmp16632;
  assign tmp16630 = s3 ? tmp15908 : tmp16631;
  assign tmp16636 = s1 ? tmp15921 : tmp15924;
  assign tmp16635 = s2 ? tmp15908 : tmp16636;
  assign tmp16639 = s0 ? tmp15424 : tmp15908;
  assign tmp16638 = s1 ? tmp15908 : tmp16639;
  assign tmp16637 = s2 ? tmp15923 : tmp16638;
  assign tmp16634 = s3 ? tmp16635 : tmp16637;
  assign tmp16629 = s4 ? tmp16630 : tmp16634;
  assign tmp16644 = s1 ? tmp15908 : tmp16633;
  assign tmp16643 = s2 ? tmp16632 : tmp16644;
  assign tmp16647 = s0 ? tmp15908 : tmp15424;
  assign tmp16646 = s1 ? tmp15472 : tmp16647;
  assign tmp16645 = s2 ? tmp15908 : tmp16646;
  assign tmp16642 = s3 ? tmp16643 : tmp16645;
  assign tmp16651 = s0 ? 1 : tmp15908;
  assign tmp16650 = s1 ? tmp16651 : tmp15468;
  assign tmp16649 = s2 ? tmp16650 : tmp15908;
  assign tmp16653 = s1 ? tmp16647 : 1;
  assign tmp16652 = s2 ? tmp16653 : 1;
  assign tmp16648 = s3 ? tmp16649 : tmp16652;
  assign tmp16641 = s4 ? tmp16642 : tmp16648;
  assign tmp16657 = s1 ? tmp16647 : tmp15424;
  assign tmp16659 = s0 ? tmp15941 : tmp15908;
  assign tmp16658 = s1 ? tmp15908 : tmp16659;
  assign tmp16656 = s2 ? tmp16657 : tmp16658;
  assign tmp16655 = s3 ? tmp16656 : tmp16505;
  assign tmp16661 = s2 ? tmp15424 : tmp15908;
  assign tmp16660 = s3 ? tmp16661 : 1;
  assign tmp16654 = s4 ? tmp16655 : tmp16660;
  assign tmp16640 = s5 ? tmp16641 : tmp16654;
  assign tmp16628 = s6 ? tmp16629 : tmp16640;
  assign tmp16624 = s7 ? tmp16625 : tmp16628;
  assign tmp16663 = s5 ? tmp16068 : tmp16627;
  assign tmp16662 = s6 ? tmp16065 : tmp16663;
  assign tmp16623 = s8 ? tmp16624 : tmp16662;
  assign tmp16621 = s9 ? tmp16622 : tmp16623;
  assign tmp16563 = s10 ? tmp16564 : tmp16621;
  assign tmp16674 = s0 ? tmp15908 : tmp15941;
  assign tmp16673 = s1 ? tmp15908 : tmp16674;
  assign tmp16672 = s2 ? tmp15424 : tmp16673;
  assign tmp16671 = s3 ? tmp16672 : 1;
  assign tmp16670 = s4 ? tmp16655 : tmp16671;
  assign tmp16669 = s5 ? tmp16641 : tmp16670;
  assign tmp16668 = s6 ? tmp16629 : tmp16669;
  assign tmp16667 = s7 ? tmp16579 : tmp16668;
  assign tmp16666 = s8 ? tmp16667 : tmp16597;
  assign tmp16665 = s9 ? tmp16622 : tmp16666;
  assign tmp16664 = s10 ? tmp16564 : tmp16665;
  assign tmp16562 = s11 ? tmp16563 : tmp16664;
  assign tmp16561 = s12 ? tmp16562 : 1;
  assign tmp16560 = s13 ? tmp15642 : tmp16561;
  assign tmp16559 = s14 ? tmp15391 : tmp16560;
  assign tmp16558 = s15 ? tmp16559 : tmp16117;
  assign tmp16304 = s16 ? tmp16305 : tmp16558;
  assign tmp15387 = ~(s17 ? tmp15388 : tmp16304);
  assign s16n = tmp15387;

  assign tmp16690 = l2 ? 1 : 0;
  assign tmp16692 = l1 ? 1 : 0;
  assign tmp16693 = ~(l2 ? 1 : 0);
  assign tmp16691 = ~(s0 ? tmp16692 : tmp16693);
  assign tmp16689 = s1 ? tmp16690 : tmp16691;
  assign tmp16696 = s0 ? tmp16690 : 0;
  assign tmp16695 = s1 ? tmp16696 : tmp16690;
  assign tmp16694 = s2 ? tmp16690 : tmp16695;
  assign tmp16688 = s3 ? tmp16689 : tmp16694;
  assign tmp16700 = ~(s0 ? tmp16692 : 1);
  assign tmp16699 = s1 ? tmp16696 : tmp16700;
  assign tmp16698 = s2 ? tmp16695 : tmp16699;
  assign tmp16703 = s0 ? 1 : 0;
  assign tmp16702 = s1 ? tmp16692 : tmp16703;
  assign tmp16705 = s0 ? 1 : tmp16690;
  assign tmp16704 = ~(s1 ? tmp16690 : tmp16705);
  assign tmp16701 = ~(s2 ? tmp16702 : tmp16704);
  assign tmp16697 = s3 ? tmp16698 : tmp16701;
  assign tmp16687 = s4 ? tmp16688 : tmp16697;
  assign tmp16710 = s1 ? tmp16696 : 0;
  assign tmp16712 = s0 ? 1 : tmp16693;
  assign tmp16711 = ~(s1 ? tmp16712 : tmp16693);
  assign tmp16709 = s2 ? tmp16710 : tmp16711;
  assign tmp16714 = s1 ? 1 : tmp16690;
  assign tmp16713 = s2 ? tmp16690 : tmp16714;
  assign tmp16708 = s3 ? tmp16709 : tmp16713;
  assign tmp16718 = ~(l1 ? 1 : 0);
  assign tmp16717 = s1 ? tmp16705 : tmp16718;
  assign tmp16720 = ~(s0 ? tmp16690 : 0);
  assign tmp16719 = ~(s1 ? tmp16692 : tmp16720);
  assign tmp16716 = s2 ? tmp16717 : tmp16719;
  assign tmp16721 = s2 ? tmp16689 : 1;
  assign tmp16715 = s3 ? tmp16716 : tmp16721;
  assign tmp16707 = s4 ? tmp16708 : tmp16715;
  assign tmp16726 = s0 ? tmp16690 : 1;
  assign tmp16725 = s1 ? tmp16726 : 1;
  assign tmp16727 = s1 ? tmp16703 : 0;
  assign tmp16724 = s2 ? tmp16725 : tmp16727;
  assign tmp16729 = ~(s1 ? 1 : tmp16705);
  assign tmp16728 = ~(s2 ? tmp16727 : tmp16729);
  assign tmp16723 = s3 ? tmp16724 : tmp16728;
  assign tmp16732 = s1 ? tmp16705 : 0;
  assign tmp16731 = s2 ? tmp16725 : tmp16732;
  assign tmp16734 = s1 ? 1 : tmp16705;
  assign tmp16735 = s1 ? tmp16705 : 1;
  assign tmp16733 = s2 ? tmp16734 : tmp16735;
  assign tmp16730 = s3 ? tmp16731 : tmp16733;
  assign tmp16722 = s4 ? tmp16723 : tmp16730;
  assign tmp16706 = s5 ? tmp16707 : tmp16722;
  assign tmp16686 = s6 ? tmp16687 : tmp16706;
  assign tmp16740 = s1 ? tmp16696 : tmp16718;
  assign tmp16739 = s2 ? tmp16695 : tmp16740;
  assign tmp16742 = s1 ? tmp16692 : 0;
  assign tmp16741 = ~(s2 ? tmp16742 : tmp16704);
  assign tmp16738 = s3 ? tmp16739 : tmp16741;
  assign tmp16737 = s4 ? tmp16688 : tmp16738;
  assign tmp16746 = s2 ? tmp16710 : tmp16690;
  assign tmp16745 = s3 ? tmp16746 : tmp16713;
  assign tmp16749 = ~(s1 ? tmp16692 : tmp16693);
  assign tmp16748 = s2 ? tmp16717 : tmp16749;
  assign tmp16747 = s3 ? tmp16748 : tmp16721;
  assign tmp16744 = s4 ? tmp16745 : tmp16747;
  assign tmp16752 = s2 ? tmp16725 : 0;
  assign tmp16753 = s2 ? 1 : tmp16714;
  assign tmp16751 = s3 ? tmp16752 : tmp16753;
  assign tmp16755 = s2 ? 1 : tmp16690;
  assign tmp16754 = s3 ? tmp16755 : tmp16714;
  assign tmp16750 = s4 ? tmp16751 : tmp16754;
  assign tmp16743 = s5 ? tmp16744 : tmp16750;
  assign tmp16736 = s6 ? tmp16737 : tmp16743;
  assign tmp16685 = s7 ? tmp16686 : tmp16736;
  assign tmp16762 = ~(s1 ? tmp16712 : tmp16720);
  assign tmp16761 = s2 ? tmp16710 : tmp16762;
  assign tmp16764 = ~(s1 ? 1 : tmp16690);
  assign tmp16763 = ~(s2 ? tmp16712 : tmp16764);
  assign tmp16760 = s3 ? tmp16761 : tmp16763;
  assign tmp16759 = s4 ? tmp16760 : tmp16715;
  assign tmp16758 = s5 ? tmp16759 : tmp16722;
  assign tmp16757 = s6 ? tmp16687 : tmp16758;
  assign tmp16770 = s1 ? tmp16690 : tmp16696;
  assign tmp16769 = s2 ? tmp16710 : tmp16770;
  assign tmp16768 = s3 ? tmp16769 : tmp16713;
  assign tmp16772 = s2 ? tmp16717 : tmp16690;
  assign tmp16773 = s2 ? tmp16690 : 1;
  assign tmp16771 = s3 ? tmp16772 : tmp16773;
  assign tmp16767 = s4 ? tmp16768 : tmp16771;
  assign tmp16766 = s5 ? tmp16767 : tmp16750;
  assign tmp16765 = s6 ? tmp16737 : tmp16766;
  assign tmp16756 = s7 ? tmp16757 : tmp16765;
  assign tmp16684 = s8 ? tmp16685 : tmp16756;
  assign tmp16781 = s0 ? tmp16692 : 1;
  assign tmp16780 = s1 ? tmp16781 : tmp16692;
  assign tmp16779 = s2 ? tmp16692 : tmp16780;
  assign tmp16778 = s3 ? tmp16692 : tmp16779;
  assign tmp16783 = s2 ? tmp16692 : tmp16781;
  assign tmp16786 = ~(s0 ? 1 : tmp16718);
  assign tmp16785 = s1 ? tmp16692 : tmp16786;
  assign tmp16784 = s2 ? tmp16702 : tmp16785;
  assign tmp16782 = s3 ? tmp16783 : tmp16784;
  assign tmp16777 = s4 ? tmp16778 : tmp16782;
  assign tmp16791 = s1 ? tmp16781 : 1;
  assign tmp16793 = s0 ? 1 : tmp16692;
  assign tmp16792 = s1 ? tmp16793 : tmp16692;
  assign tmp16790 = s2 ? tmp16791 : tmp16792;
  assign tmp16795 = ~(s1 ? 1 : tmp16718);
  assign tmp16794 = s2 ? tmp16692 : tmp16795;
  assign tmp16789 = s3 ? tmp16790 : tmp16794;
  assign tmp16799 = s0 ? 1 : tmp16718;
  assign tmp16798 = s1 ? tmp16799 : tmp16718;
  assign tmp16797 = s2 ? tmp16798 : tmp16718;
  assign tmp16800 = ~(s2 ? tmp16692 : 0);
  assign tmp16796 = ~(s3 ? tmp16797 : tmp16800);
  assign tmp16788 = s4 ? tmp16789 : tmp16796;
  assign tmp16805 = s0 ? tmp16692 : 0;
  assign tmp16804 = s1 ? tmp16805 : 0;
  assign tmp16806 = ~(s1 ? tmp16703 : 0);
  assign tmp16803 = s2 ? tmp16804 : tmp16806;
  assign tmp16808 = ~(s1 ? 1 : tmp16799);
  assign tmp16807 = s2 ? tmp16727 : tmp16808;
  assign tmp16802 = s3 ? tmp16803 : tmp16807;
  assign tmp16811 = ~(s1 ? tmp16799 : 0);
  assign tmp16810 = s2 ? tmp16804 : tmp16811;
  assign tmp16813 = s1 ? 1 : tmp16799;
  assign tmp16814 = s1 ? tmp16799 : 1;
  assign tmp16812 = ~(s2 ? tmp16813 : tmp16814);
  assign tmp16809 = s3 ? tmp16810 : tmp16812;
  assign tmp16801 = s4 ? tmp16802 : tmp16809;
  assign tmp16787 = s5 ? tmp16788 : tmp16801;
  assign tmp16776 = s6 ? tmp16777 : tmp16787;
  assign tmp16818 = s2 ? tmp16742 : tmp16785;
  assign tmp16817 = s3 ? tmp16779 : tmp16818;
  assign tmp16816 = s4 ? tmp16778 : tmp16817;
  assign tmp16822 = s2 ? tmp16791 : tmp16692;
  assign tmp16821 = s3 ? tmp16822 : tmp16794;
  assign tmp16820 = s4 ? tmp16821 : tmp16796;
  assign tmp16825 = s2 ? tmp16804 : 1;
  assign tmp16827 = s1 ? 1 : tmp16718;
  assign tmp16826 = ~(s2 ? 1 : tmp16827);
  assign tmp16824 = s3 ? tmp16825 : tmp16826;
  assign tmp16829 = s2 ? 1 : tmp16718;
  assign tmp16828 = ~(s3 ? tmp16829 : tmp16827);
  assign tmp16823 = s4 ? tmp16824 : tmp16828;
  assign tmp16819 = s5 ? tmp16820 : tmp16823;
  assign tmp16815 = s6 ? tmp16816 : tmp16819;
  assign tmp16775 = ~(s7 ? tmp16776 : tmp16815);
  assign tmp16774 = s8 ? tmp16756 : tmp16775;
  assign tmp16683 = s9 ? tmp16684 : tmp16774;
  assign tmp16835 = s4 ? tmp16745 : tmp16771;
  assign tmp16834 = s5 ? tmp16835 : tmp16750;
  assign tmp16833 = s6 ? tmp16737 : tmp16834;
  assign tmp16832 = s7 ? tmp16686 : tmp16833;
  assign tmp16831 = s8 ? tmp16832 : tmp16686;
  assign tmp16841 = s3 ? tmp16748 : tmp16773;
  assign tmp16840 = s4 ? tmp16745 : tmp16841;
  assign tmp16839 = s5 ? tmp16840 : tmp16750;
  assign tmp16838 = s6 ? tmp16737 : tmp16839;
  assign tmp16842 = ~(s6 ? tmp16816 : tmp16819);
  assign tmp16837 = s7 ? tmp16838 : tmp16842;
  assign tmp16843 = s7 ? tmp16765 : tmp16833;
  assign tmp16836 = s8 ? tmp16837 : tmp16843;
  assign tmp16830 = s9 ? tmp16831 : tmp16836;
  assign tmp16682 = s10 ? tmp16683 : tmp16830;
  assign tmp16847 = s7 ? tmp16736 : tmp16842;
  assign tmp16846 = s8 ? tmp16847 : tmp16843;
  assign tmp16845 = s9 ? tmp16831 : tmp16846;
  assign tmp16844 = s10 ? tmp16683 : tmp16845;
  assign tmp16681 = ~(s11 ? tmp16682 : tmp16844);
  assign tmp16680 = s12 ? 1 : tmp16681;
  assign tmp16858 = l1 ? tmp16690 : 0;
  assign tmp16860 = ~(l1 ? tmp16690 : 0);
  assign tmp16859 = ~(s0 ? 1 : tmp16860);
  assign tmp16857 = s1 ? tmp16858 : tmp16859;
  assign tmp16863 = s0 ? tmp16858 : 0;
  assign tmp16862 = s1 ? tmp16863 : tmp16858;
  assign tmp16861 = s2 ? tmp16858 : tmp16862;
  assign tmp16856 = s3 ? tmp16857 : tmp16861;
  assign tmp16866 = s1 ? tmp16863 : 0;
  assign tmp16865 = s2 ? tmp16862 : tmp16866;
  assign tmp16868 = s1 ? 1 : tmp16703;
  assign tmp16870 = s0 ? 1 : tmp16858;
  assign tmp16869 = ~(s1 ? tmp16858 : tmp16870);
  assign tmp16867 = ~(s2 ? tmp16868 : tmp16869);
  assign tmp16864 = s3 ? tmp16865 : tmp16867;
  assign tmp16855 = s4 ? tmp16856 : tmp16864;
  assign tmp16875 = s1 ? tmp16863 : tmp16859;
  assign tmp16877 = s0 ? 1 : tmp16860;
  assign tmp16878 = ~(s0 ? tmp16858 : 0);
  assign tmp16876 = ~(s1 ? tmp16877 : tmp16878);
  assign tmp16874 = s2 ? tmp16875 : tmp16876;
  assign tmp16880 = ~(s1 ? 1 : tmp16858);
  assign tmp16879 = ~(s2 ? tmp16877 : tmp16880);
  assign tmp16873 = s3 ? tmp16874 : tmp16879;
  assign tmp16883 = s1 ? tmp16870 : 0;
  assign tmp16884 = ~(s1 ? 1 : tmp16878);
  assign tmp16882 = s2 ? tmp16883 : tmp16884;
  assign tmp16887 = ~(s0 ? 1 : tmp16693);
  assign tmp16886 = s1 ? tmp16858 : tmp16887;
  assign tmp16885 = s2 ? tmp16886 : 1;
  assign tmp16881 = s3 ? tmp16882 : tmp16885;
  assign tmp16872 = s4 ? tmp16873 : tmp16881;
  assign tmp16892 = s0 ? tmp16858 : 1;
  assign tmp16891 = s1 ? tmp16892 : 1;
  assign tmp16890 = s2 ? tmp16891 : tmp16858;
  assign tmp16893 = s2 ? tmp16725 : tmp16734;
  assign tmp16889 = s3 ? tmp16890 : tmp16893;
  assign tmp16896 = s1 ? tmp16870 : tmp16858;
  assign tmp16895 = s2 ? tmp16690 : tmp16896;
  assign tmp16894 = s3 ? tmp16895 : tmp16733;
  assign tmp16888 = s4 ? tmp16889 : tmp16894;
  assign tmp16871 = s5 ? tmp16872 : tmp16888;
  assign tmp16854 = s6 ? tmp16855 : tmp16871;
  assign tmp16901 = s1 ? 1 : 0;
  assign tmp16900 = ~(s2 ? tmp16901 : tmp16869);
  assign tmp16899 = s3 ? tmp16865 : tmp16900;
  assign tmp16898 = s4 ? tmp16856 : tmp16899;
  assign tmp16906 = s1 ? tmp16858 : tmp16863;
  assign tmp16905 = s2 ? tmp16862 : tmp16906;
  assign tmp16908 = s1 ? 1 : tmp16858;
  assign tmp16907 = s2 ? tmp16858 : tmp16908;
  assign tmp16904 = s3 ? tmp16905 : tmp16907;
  assign tmp16910 = s2 ? tmp16883 : tmp16858;
  assign tmp16912 = s1 ? tmp16858 : tmp16690;
  assign tmp16911 = s2 ? tmp16912 : 1;
  assign tmp16909 = s3 ? tmp16910 : tmp16911;
  assign tmp16903 = s4 ? tmp16904 : tmp16909;
  assign tmp16915 = s2 ? tmp16891 : tmp16714;
  assign tmp16914 = s3 ? tmp16890 : tmp16915;
  assign tmp16917 = s2 ? 1 : tmp16858;
  assign tmp16916 = s3 ? tmp16917 : tmp16690;
  assign tmp16913 = s4 ? tmp16914 : tmp16916;
  assign tmp16902 = s5 ? tmp16903 : tmp16913;
  assign tmp16897 = s6 ? tmp16898 : tmp16902;
  assign tmp16853 = s7 ? tmp16854 : tmp16897;
  assign tmp16924 = ~(l3 ? 1 : 0);
  assign tmp16923 = l1 ? tmp16690 : tmp16924;
  assign tmp16927 = l3 ? 1 : 0;
  assign tmp16926 = l1 ? 1 : tmp16927;
  assign tmp16928 = ~(l1 ? tmp16690 : tmp16924);
  assign tmp16925 = ~(s0 ? tmp16926 : tmp16928);
  assign tmp16922 = s1 ? tmp16923 : tmp16925;
  assign tmp16931 = s0 ? tmp16923 : tmp16924;
  assign tmp16930 = s1 ? tmp16931 : tmp16923;
  assign tmp16929 = s2 ? tmp16923 : tmp16930;
  assign tmp16921 = s3 ? tmp16922 : tmp16929;
  assign tmp16935 = s0 ? tmp16923 : 0;
  assign tmp16934 = s1 ? tmp16935 : tmp16923;
  assign tmp16937 = ~(s0 ? tmp16926 : 1);
  assign tmp16936 = s1 ? tmp16935 : tmp16937;
  assign tmp16933 = s2 ? tmp16934 : tmp16936;
  assign tmp16939 = s1 ? tmp16926 : tmp16703;
  assign tmp16941 = s0 ? 1 : tmp16923;
  assign tmp16940 = ~(s1 ? tmp16923 : tmp16941);
  assign tmp16938 = ~(s2 ? tmp16939 : tmp16940);
  assign tmp16932 = s3 ? tmp16933 : tmp16938;
  assign tmp16920 = s4 ? tmp16921 : tmp16932;
  assign tmp16947 = ~(s0 ? 1 : tmp16928);
  assign tmp16946 = s1 ? tmp16935 : tmp16947;
  assign tmp16949 = s0 ? 1 : tmp16928;
  assign tmp16950 = ~(s0 ? tmp16923 : tmp16924);
  assign tmp16948 = ~(s1 ? tmp16949 : tmp16950);
  assign tmp16945 = s2 ? tmp16946 : tmp16948;
  assign tmp16952 = s0 ? tmp16927 : tmp16928;
  assign tmp16953 = ~(s1 ? 1 : tmp16923);
  assign tmp16951 = ~(s2 ? tmp16952 : tmp16953);
  assign tmp16944 = s3 ? tmp16945 : tmp16951;
  assign tmp16957 = ~(s0 ? 1 : tmp16692);
  assign tmp16956 = s1 ? tmp16941 : tmp16957;
  assign tmp16959 = ~(s0 ? tmp16923 : 0);
  assign tmp16958 = ~(s1 ? tmp16793 : tmp16959);
  assign tmp16955 = s2 ? tmp16956 : tmp16958;
  assign tmp16961 = s1 ? tmp16923 : tmp16691;
  assign tmp16960 = s2 ? tmp16961 : 1;
  assign tmp16954 = s3 ? tmp16955 : tmp16960;
  assign tmp16943 = s4 ? tmp16944 : tmp16954;
  assign tmp16966 = s0 ? tmp16923 : 1;
  assign tmp16965 = s1 ? tmp16966 : 1;
  assign tmp16968 = s0 ? tmp16690 : tmp16923;
  assign tmp16967 = s1 ? tmp16941 : tmp16968;
  assign tmp16964 = s2 ? tmp16965 : tmp16967;
  assign tmp16963 = s3 ? tmp16964 : tmp16893;
  assign tmp16971 = s1 ? tmp16690 : 1;
  assign tmp16973 = s0 ? tmp16923 : tmp16690;
  assign tmp16972 = s1 ? tmp16941 : tmp16973;
  assign tmp16970 = s2 ? tmp16971 : tmp16972;
  assign tmp16969 = s3 ? tmp16970 : tmp16733;
  assign tmp16962 = s4 ? tmp16963 : tmp16969;
  assign tmp16942 = s5 ? tmp16943 : tmp16962;
  assign tmp16919 = s6 ? tmp16920 : tmp16942;
  assign tmp16979 = ~(l1 ? 1 : tmp16927);
  assign tmp16978 = s1 ? tmp16935 : tmp16979;
  assign tmp16977 = s2 ? tmp16934 : tmp16978;
  assign tmp16981 = s1 ? tmp16926 : 0;
  assign tmp16980 = ~(s2 ? tmp16981 : tmp16940);
  assign tmp16976 = s3 ? tmp16977 : tmp16980;
  assign tmp16975 = s4 ? tmp16921 : tmp16976;
  assign tmp16986 = s1 ? tmp16923 : tmp16931;
  assign tmp16985 = s2 ? tmp16934 : tmp16986;
  assign tmp16988 = s1 ? 1 : tmp16923;
  assign tmp16987 = s2 ? tmp16923 : tmp16988;
  assign tmp16984 = s3 ? tmp16985 : tmp16987;
  assign tmp16990 = s2 ? tmp16956 : tmp16923;
  assign tmp16992 = s1 ? tmp16923 : tmp16690;
  assign tmp16991 = s2 ? tmp16992 : 1;
  assign tmp16989 = s3 ? tmp16990 : tmp16991;
  assign tmp16983 = s4 ? tmp16984 : tmp16989;
  assign tmp16995 = s2 ? tmp16965 : tmp16992;
  assign tmp16994 = s3 ? tmp16995 : tmp16915;
  assign tmp16998 = s1 ? tmp16923 : tmp16858;
  assign tmp16997 = s2 ? 1 : tmp16998;
  assign tmp16996 = s3 ? tmp16997 : tmp16690;
  assign tmp16993 = s4 ? tmp16994 : tmp16996;
  assign tmp16982 = s5 ? tmp16983 : tmp16993;
  assign tmp16974 = s6 ? tmp16975 : tmp16982;
  assign tmp16918 = s7 ? tmp16919 : tmp16974;
  assign tmp16852 = s8 ? tmp16853 : tmp16918;
  assign tmp17007 = s0 ? tmp16690 : tmp16858;
  assign tmp17006 = s1 ? tmp17007 : tmp16858;
  assign tmp17005 = s2 ? tmp16891 : tmp17006;
  assign tmp17004 = s3 ? tmp17005 : tmp16893;
  assign tmp17003 = s4 ? tmp17004 : tmp16894;
  assign tmp17002 = s5 ? tmp16872 : tmp17003;
  assign tmp17001 = s6 ? tmp16855 : tmp17002;
  assign tmp17012 = s2 ? tmp16891 : tmp16912;
  assign tmp17013 = s2 ? tmp16725 : tmp16714;
  assign tmp17011 = s3 ? tmp17012 : tmp17013;
  assign tmp17010 = s4 ? tmp17011 : tmp16916;
  assign tmp17009 = s5 ? tmp16903 : tmp17010;
  assign tmp17008 = s6 ? tmp16898 : tmp17009;
  assign tmp17000 = s7 ? tmp17001 : tmp17008;
  assign tmp16999 = s8 ? tmp16918 : tmp17000;
  assign tmp16851 = s9 ? tmp16852 : tmp16999;
  assign tmp17020 = s3 ? tmp17012 : tmp16915;
  assign tmp17019 = s4 ? tmp17020 : tmp16916;
  assign tmp17018 = s5 ? tmp16903 : tmp17019;
  assign tmp17017 = s6 ? tmp16898 : tmp17018;
  assign tmp17016 = s7 ? tmp16854 : tmp17017;
  assign tmp17015 = s8 ? tmp17016 : tmp16854;
  assign tmp17022 = s7 ? tmp16897 : tmp17008;
  assign tmp17028 = s2 ? 1 : tmp16923;
  assign tmp17027 = s3 ? tmp17028 : tmp16690;
  assign tmp17026 = s4 ? tmp16994 : tmp17027;
  assign tmp17025 = s5 ? tmp16983 : tmp17026;
  assign tmp17024 = s6 ? tmp16975 : tmp17025;
  assign tmp17023 = s7 ? tmp17024 : tmp17017;
  assign tmp17021 = s8 ? tmp17022 : tmp17023;
  assign tmp17014 = s9 ? tmp17015 : tmp17021;
  assign tmp16850 = s10 ? tmp16851 : tmp17014;
  assign tmp17032 = s7 ? tmp16974 : tmp17017;
  assign tmp17031 = s8 ? tmp17022 : tmp17032;
  assign tmp17030 = s9 ? tmp17015 : tmp17031;
  assign tmp17029 = s10 ? tmp16851 : tmp17030;
  assign tmp16849 = s11 ? tmp16850 : tmp17029;
  assign tmp17041 = s1 ? tmp16690 : tmp16887;
  assign tmp17040 = s3 ? tmp17041 : tmp16694;
  assign tmp17043 = s2 ? tmp16695 : tmp16710;
  assign tmp17044 = ~(s2 ? tmp16868 : tmp16693);
  assign tmp17042 = s3 ? tmp17043 : tmp17044;
  assign tmp17039 = s4 ? tmp17040 : tmp17042;
  assign tmp17049 = s1 ? tmp16696 : tmp16887;
  assign tmp17048 = s2 ? tmp17049 : tmp16762;
  assign tmp17047 = s3 ? tmp17048 : tmp16763;
  assign tmp17052 = ~(s1 ? 1 : tmp16720);
  assign tmp17051 = s2 ? tmp16732 : tmp17052;
  assign tmp17053 = s2 ? tmp17041 : 1;
  assign tmp17050 = s3 ? tmp17051 : tmp17053;
  assign tmp17046 = s4 ? tmp17047 : tmp17050;
  assign tmp17056 = s2 ? tmp16725 : tmp16690;
  assign tmp17055 = s3 ? tmp17056 : tmp16893;
  assign tmp17059 = s1 ? tmp16705 : tmp16690;
  assign tmp17058 = s2 ? tmp16690 : tmp17059;
  assign tmp17057 = s3 ? tmp17058 : tmp16733;
  assign tmp17054 = s4 ? tmp17055 : tmp17057;
  assign tmp17045 = s5 ? tmp17046 : tmp17054;
  assign tmp17038 = s6 ? tmp17039 : tmp17045;
  assign tmp17063 = ~(s2 ? tmp16901 : tmp16693);
  assign tmp17062 = s3 ? tmp17043 : tmp17063;
  assign tmp17061 = s4 ? tmp17040 : tmp17062;
  assign tmp17067 = s2 ? tmp16695 : tmp16770;
  assign tmp17066 = s3 ? tmp17067 : tmp16713;
  assign tmp17069 = s2 ? tmp16732 : tmp16690;
  assign tmp17068 = s3 ? tmp17069 : tmp16773;
  assign tmp17065 = s4 ? tmp17066 : tmp17068;
  assign tmp17071 = s3 ? tmp17056 : tmp16915;
  assign tmp17072 = s3 ? tmp16858 : tmp16690;
  assign tmp17070 = s4 ? tmp17071 : tmp17072;
  assign tmp17064 = s5 ? tmp17065 : tmp17070;
  assign tmp17060 = s6 ? tmp17061 : tmp17064;
  assign tmp17037 = s7 ? tmp17038 : tmp17060;
  assign tmp17078 = l1 ? tmp16690 : 1;
  assign tmp17080 = ~(l1 ? tmp16690 : 1);
  assign tmp17079 = ~(s0 ? tmp16692 : tmp17080);
  assign tmp17077 = s1 ? tmp17078 : tmp17079;
  assign tmp17083 = s0 ? tmp17078 : 1;
  assign tmp17082 = s1 ? tmp17083 : tmp17078;
  assign tmp17081 = s2 ? tmp17078 : tmp17082;
  assign tmp17076 = s3 ? tmp17077 : tmp17081;
  assign tmp17087 = s0 ? tmp17078 : 0;
  assign tmp17086 = s1 ? tmp17087 : tmp17078;
  assign tmp17088 = s1 ? tmp17087 : tmp16700;
  assign tmp17085 = s2 ? tmp17086 : tmp17088;
  assign tmp17089 = ~(s2 ? tmp16702 : tmp17080);
  assign tmp17084 = s3 ? tmp17085 : tmp17089;
  assign tmp17075 = s4 ? tmp17076 : tmp17084;
  assign tmp17095 = ~(s0 ? 1 : tmp17080);
  assign tmp17094 = s1 ? tmp17087 : tmp17095;
  assign tmp17097 = s0 ? 1 : tmp17080;
  assign tmp17098 = ~(s0 ? tmp17078 : 1);
  assign tmp17096 = ~(s1 ? tmp17097 : tmp17098);
  assign tmp17093 = s2 ? tmp17094 : tmp17096;
  assign tmp17100 = s0 ? 1 : tmp17078;
  assign tmp17101 = s1 ? 1 : tmp17078;
  assign tmp17099 = s2 ? tmp17100 : tmp17101;
  assign tmp17092 = s3 ? tmp17093 : tmp17099;
  assign tmp17104 = s1 ? tmp17100 : tmp16957;
  assign tmp17106 = ~(s0 ? tmp17078 : 0);
  assign tmp17105 = ~(s1 ? tmp16793 : tmp17106);
  assign tmp17103 = s2 ? tmp17104 : tmp17105;
  assign tmp17108 = s1 ? tmp17078 : tmp16691;
  assign tmp17107 = s2 ? tmp17108 : 1;
  assign tmp17102 = s3 ? tmp17103 : tmp17107;
  assign tmp17091 = s4 ? tmp17092 : tmp17102;
  assign tmp17112 = s1 ? tmp17083 : 1;
  assign tmp17114 = s0 ? tmp16690 : tmp17078;
  assign tmp17113 = s1 ? tmp17078 : tmp17114;
  assign tmp17111 = s2 ? tmp17112 : tmp17113;
  assign tmp17110 = s3 ? tmp17111 : tmp16893;
  assign tmp17118 = s0 ? tmp17078 : tmp16690;
  assign tmp17117 = s1 ? tmp17100 : tmp17118;
  assign tmp17116 = s2 ? tmp16971 : tmp17117;
  assign tmp17115 = s3 ? tmp17116 : tmp16733;
  assign tmp17109 = s4 ? tmp17110 : tmp17115;
  assign tmp17090 = s5 ? tmp17091 : tmp17109;
  assign tmp17074 = s6 ? tmp17075 : tmp17090;
  assign tmp17123 = s1 ? tmp17087 : tmp16718;
  assign tmp17122 = s2 ? tmp17086 : tmp17123;
  assign tmp17124 = ~(s2 ? tmp16742 : tmp17080);
  assign tmp17121 = s3 ? tmp17122 : tmp17124;
  assign tmp17120 = s4 ? tmp17076 : tmp17121;
  assign tmp17129 = s1 ? tmp17078 : tmp17083;
  assign tmp17128 = s2 ? tmp17086 : tmp17129;
  assign tmp17130 = s2 ? tmp17078 : tmp17101;
  assign tmp17127 = s3 ? tmp17128 : tmp17130;
  assign tmp17132 = s2 ? tmp17104 : tmp17078;
  assign tmp17134 = s1 ? tmp17078 : tmp16690;
  assign tmp17133 = s2 ? tmp17134 : 1;
  assign tmp17131 = s3 ? tmp17132 : tmp17133;
  assign tmp17126 = s4 ? tmp17127 : tmp17131;
  assign tmp17137 = s2 ? tmp17112 : tmp17134;
  assign tmp17136 = s3 ? tmp17137 : tmp16915;
  assign tmp17140 = s1 ? tmp17078 : tmp16858;
  assign tmp17139 = s2 ? 1 : tmp17140;
  assign tmp17138 = s3 ? tmp17139 : tmp16690;
  assign tmp17135 = s4 ? tmp17136 : tmp17138;
  assign tmp17125 = s5 ? tmp17126 : tmp17135;
  assign tmp17119 = s6 ? tmp17120 : tmp17125;
  assign tmp17073 = s7 ? tmp17074 : tmp17119;
  assign tmp17036 = s8 ? tmp17037 : tmp17073;
  assign tmp17147 = s2 ? tmp17049 : tmp16711;
  assign tmp17146 = s3 ? tmp17147 : tmp16713;
  assign tmp17145 = s4 ? tmp17146 : tmp17050;
  assign tmp17144 = s5 ? tmp17145 : tmp17054;
  assign tmp17143 = s6 ? tmp17039 : tmp17144;
  assign tmp17152 = s2 ? tmp16695 : tmp16690;
  assign tmp17151 = s3 ? tmp17152 : tmp16713;
  assign tmp17150 = s4 ? tmp17151 : tmp17068;
  assign tmp17154 = s3 ? tmp17056 : tmp17013;
  assign tmp17153 = s4 ? tmp17154 : tmp16690;
  assign tmp17149 = s5 ? tmp17150 : tmp17153;
  assign tmp17148 = s6 ? tmp17061 : tmp17149;
  assign tmp17142 = s7 ? tmp17143 : tmp17148;
  assign tmp17141 = s8 ? tmp17073 : tmp17142;
  assign tmp17035 = s9 ? tmp17036 : tmp17141;
  assign tmp17159 = s5 ? tmp17150 : tmp17070;
  assign tmp17158 = s6 ? tmp17061 : tmp17159;
  assign tmp17157 = s7 ? tmp17143 : tmp17158;
  assign tmp17156 = s8 ? tmp17157 : tmp17143;
  assign tmp17164 = s3 ? tmp16755 : tmp16690;
  assign tmp17163 = s4 ? tmp17071 : tmp17164;
  assign tmp17162 = s5 ? tmp17065 : tmp17163;
  assign tmp17161 = s6 ? tmp17061 : tmp17162;
  assign tmp17170 = s2 ? 1 : tmp17078;
  assign tmp17169 = s3 ? tmp17170 : tmp16690;
  assign tmp17168 = s4 ? tmp17136 : tmp17169;
  assign tmp17167 = s5 ? tmp17126 : tmp17168;
  assign tmp17166 = s6 ? tmp17120 : tmp17167;
  assign tmp17172 = s5 ? tmp17150 : tmp17163;
  assign tmp17171 = s6 ? tmp17061 : tmp17172;
  assign tmp17165 = s7 ? tmp17166 : tmp17171;
  assign tmp17160 = s8 ? tmp17161 : tmp17165;
  assign tmp17155 = s9 ? tmp17156 : tmp17160;
  assign tmp17034 = s10 ? tmp17035 : tmp17155;
  assign tmp17176 = s7 ? tmp17119 : tmp17158;
  assign tmp17175 = s8 ? tmp17060 : tmp17176;
  assign tmp17174 = s9 ? tmp17156 : tmp17175;
  assign tmp17173 = s10 ? tmp17035 : tmp17174;
  assign tmp17033 = s11 ? tmp17034 : tmp17173;
  assign tmp16848 = ~(s12 ? tmp16849 : tmp17033);
  assign tmp16679 = s13 ? tmp16680 : tmp16848;
  assign tmp16678 = s14 ? 1 : tmp16679;
  assign tmp17191 = ~(l4 ? 1 : 0);
  assign tmp17190 = l2 ? 1 : tmp17191;
  assign tmp17189 = l1 ? tmp16690 : tmp17190;
  assign tmp17193 = ~(l1 ? tmp16690 : tmp17190);
  assign tmp17192 = ~(s0 ? tmp16692 : tmp17193);
  assign tmp17188 = s1 ? tmp17189 : tmp17192;
  assign tmp17195 = s1 ? tmp16696 : tmp17189;
  assign tmp17194 = s2 ? tmp17189 : tmp17195;
  assign tmp17187 = s3 ? tmp17188 : tmp17194;
  assign tmp17199 = s0 ? tmp17189 : 0;
  assign tmp17198 = s1 ? tmp17199 : tmp17189;
  assign tmp17200 = s1 ? tmp17199 : tmp16700;
  assign tmp17197 = s2 ? tmp17198 : tmp17200;
  assign tmp17203 = s0 ? tmp17078 : tmp17189;
  assign tmp17202 = ~(s1 ? tmp17189 : tmp17203);
  assign tmp17201 = ~(s2 ? tmp16702 : tmp17202);
  assign tmp17196 = s3 ? tmp17197 : tmp17201;
  assign tmp17186 = s4 ? tmp17187 : tmp17196;
  assign tmp17208 = s1 ? tmp17199 : tmp16887;
  assign tmp17210 = s0 ? 1 : tmp17193;
  assign tmp17211 = ~(s0 ? tmp17189 : 0);
  assign tmp17209 = ~(s1 ? tmp17210 : tmp17211);
  assign tmp17207 = s2 ? tmp17208 : tmp17209;
  assign tmp17213 = ~(s1 ? tmp17083 : tmp17189);
  assign tmp17212 = ~(s2 ? tmp17210 : tmp17213);
  assign tmp17206 = s3 ? tmp17207 : tmp17212;
  assign tmp17217 = s0 ? 1 : tmp17189;
  assign tmp17216 = s1 ? tmp17217 : tmp16718;
  assign tmp17218 = ~(s1 ? tmp16692 : tmp17211);
  assign tmp17215 = s2 ? tmp17216 : tmp17218;
  assign tmp17219 = s2 ? tmp17188 : 1;
  assign tmp17214 = s3 ? tmp17215 : tmp17219;
  assign tmp17205 = s4 ? tmp17206 : tmp17214;
  assign tmp17224 = s0 ? tmp17189 : 1;
  assign tmp17223 = s1 ? tmp17224 : 1;
  assign tmp17222 = s2 ? tmp17223 : tmp17059;
  assign tmp17226 = s1 ? 1 : tmp17217;
  assign tmp17225 = s2 ? tmp16725 : tmp17226;
  assign tmp17221 = s3 ? tmp17222 : tmp17225;
  assign tmp17229 = s1 ? tmp17224 : tmp17100;
  assign tmp17230 = s1 ? tmp17217 : tmp16690;
  assign tmp17228 = s2 ? tmp17229 : tmp17230;
  assign tmp17232 = s1 ? tmp17217 : 1;
  assign tmp17231 = s2 ? tmp17226 : tmp17232;
  assign tmp17227 = s3 ? tmp17228 : tmp17231;
  assign tmp17220 = s4 ? tmp17221 : tmp17227;
  assign tmp17204 = s5 ? tmp17205 : tmp17220;
  assign tmp17185 = s6 ? tmp17186 : tmp17204;
  assign tmp17237 = s1 ? tmp17199 : tmp16718;
  assign tmp17236 = s2 ? tmp17198 : tmp17237;
  assign tmp17238 = ~(s2 ? tmp16742 : tmp17202);
  assign tmp17235 = s3 ? tmp17236 : tmp17238;
  assign tmp17234 = s4 ? tmp17187 : tmp17235;
  assign tmp17243 = s1 ? tmp17199 : tmp16690;
  assign tmp17244 = s1 ? tmp17189 : tmp17199;
  assign tmp17242 = s2 ? tmp17243 : tmp17244;
  assign tmp17246 = s1 ? tmp17083 : tmp17189;
  assign tmp17245 = s2 ? tmp17189 : tmp17246;
  assign tmp17241 = s3 ? tmp17242 : tmp17245;
  assign tmp17249 = ~(s1 ? tmp16692 : tmp17193);
  assign tmp17248 = s2 ? tmp17216 : tmp17249;
  assign tmp17247 = s3 ? tmp17248 : tmp17219;
  assign tmp17240 = s4 ? tmp17241 : tmp17247;
  assign tmp17252 = s2 ? tmp17223 : tmp16690;
  assign tmp17254 = s1 ? 1 : tmp17189;
  assign tmp17253 = s2 ? tmp16891 : tmp17254;
  assign tmp17251 = s3 ? tmp17252 : tmp17253;
  assign tmp17257 = s1 ? tmp17224 : tmp17078;
  assign tmp17256 = s2 ? tmp17257 : tmp17189;
  assign tmp17258 = s2 ? tmp17254 : tmp17189;
  assign tmp17255 = s3 ? tmp17256 : tmp17258;
  assign tmp17250 = s4 ? tmp17251 : tmp17255;
  assign tmp17239 = s5 ? tmp17240 : tmp17250;
  assign tmp17233 = s6 ? tmp17234 : tmp17239;
  assign tmp17184 = s7 ? tmp17185 : tmp17233;
  assign tmp17262 = s3 ? tmp17188 : tmp17245;
  assign tmp17261 = s4 ? tmp17262 : tmp17196;
  assign tmp17267 = s1 ? tmp17199 : tmp17095;
  assign tmp17269 = ~(s0 ? tmp17189 : 1);
  assign tmp17268 = ~(s1 ? tmp17210 : tmp17269);
  assign tmp17266 = s2 ? tmp17267 : tmp17268;
  assign tmp17270 = s2 ? tmp17217 : tmp17254;
  assign tmp17265 = s3 ? tmp17266 : tmp17270;
  assign tmp17273 = s1 ? tmp17217 : tmp16957;
  assign tmp17274 = ~(s1 ? tmp16793 : tmp17211);
  assign tmp17272 = s2 ? tmp17273 : tmp17274;
  assign tmp17271 = s3 ? tmp17272 : tmp17219;
  assign tmp17264 = s4 ? tmp17265 : tmp17271;
  assign tmp17278 = s1 ? tmp17100 : tmp17114;
  assign tmp17277 = s2 ? tmp17223 : tmp17278;
  assign tmp17276 = s3 ? tmp17277 : tmp17225;
  assign tmp17281 = s1 ? tmp17217 : tmp17118;
  assign tmp17280 = s2 ? tmp17223 : tmp17281;
  assign tmp17279 = s3 ? tmp17280 : tmp17231;
  assign tmp17275 = s4 ? tmp17276 : tmp17279;
  assign tmp17263 = s5 ? tmp17264 : tmp17275;
  assign tmp17260 = s6 ? tmp17261 : tmp17263;
  assign tmp17283 = s4 ? tmp17262 : tmp17235;
  assign tmp17288 = s1 ? tmp17199 : tmp17078;
  assign tmp17289 = s1 ? tmp17189 : tmp17224;
  assign tmp17287 = s2 ? tmp17288 : tmp17289;
  assign tmp17290 = s2 ? tmp17189 : tmp17254;
  assign tmp17286 = s3 ? tmp17287 : tmp17290;
  assign tmp17292 = s2 ? tmp17273 : tmp17189;
  assign tmp17293 = s2 ? tmp17189 : 1;
  assign tmp17291 = s3 ? tmp17292 : tmp17293;
  assign tmp17285 = s4 ? tmp17286 : tmp17291;
  assign tmp17296 = s2 ? tmp17223 : tmp17134;
  assign tmp17295 = s3 ? tmp17296 : tmp17253;
  assign tmp17298 = s2 ? tmp17223 : tmp17189;
  assign tmp17297 = s3 ? tmp17298 : tmp17258;
  assign tmp17294 = s4 ? tmp17295 : tmp17297;
  assign tmp17284 = s5 ? tmp17285 : tmp17294;
  assign tmp17282 = s6 ? tmp17283 : tmp17284;
  assign tmp17259 = s7 ? tmp17260 : tmp17282;
  assign tmp17183 = s8 ? tmp17184 : tmp17259;
  assign tmp17304 = s2 ? tmp17078 : tmp17086;
  assign tmp17303 = s3 ? tmp17077 : tmp17304;
  assign tmp17302 = s4 ? tmp17303 : tmp17084;
  assign tmp17309 = s1 ? tmp17087 : tmp16887;
  assign tmp17311 = ~(s0 ? tmp17078 : tmp16690);
  assign tmp17310 = ~(s1 ? tmp17097 : tmp17311);
  assign tmp17308 = s2 ? tmp17309 : tmp17310;
  assign tmp17312 = s2 ? tmp17114 : tmp17082;
  assign tmp17307 = s3 ? tmp17308 : tmp17312;
  assign tmp17315 = s1 ? tmp17100 : tmp16718;
  assign tmp17316 = ~(s1 ? tmp16692 : tmp17106);
  assign tmp17314 = s2 ? tmp17315 : tmp17316;
  assign tmp17317 = s2 ? tmp17077 : 1;
  assign tmp17313 = s3 ? tmp17314 : tmp17317;
  assign tmp17306 = s4 ? tmp17307 : tmp17313;
  assign tmp17320 = s2 ? tmp17112 : tmp17059;
  assign tmp17322 = s1 ? 1 : tmp17100;
  assign tmp17321 = s2 ? tmp16725 : tmp17322;
  assign tmp17319 = s3 ? tmp17320 : tmp17321;
  assign tmp17325 = s1 ? tmp17083 : tmp17100;
  assign tmp17326 = s1 ? tmp17100 : tmp16690;
  assign tmp17324 = s2 ? tmp17325 : tmp17326;
  assign tmp17328 = s1 ? tmp17100 : 1;
  assign tmp17327 = s2 ? tmp17322 : tmp17328;
  assign tmp17323 = s3 ? tmp17324 : tmp17327;
  assign tmp17318 = s4 ? tmp17319 : tmp17323;
  assign tmp17305 = s5 ? tmp17306 : tmp17318;
  assign tmp17301 = s6 ? tmp17302 : tmp17305;
  assign tmp17330 = s4 ? tmp17303 : tmp17121;
  assign tmp17335 = s1 ? tmp17087 : tmp16690;
  assign tmp17336 = s1 ? tmp17078 : tmp17118;
  assign tmp17334 = s2 ? tmp17335 : tmp17336;
  assign tmp17333 = s3 ? tmp17334 : tmp17081;
  assign tmp17338 = s2 ? tmp17315 : tmp17078;
  assign tmp17339 = s2 ? tmp17078 : 1;
  assign tmp17337 = s3 ? tmp17338 : tmp17339;
  assign tmp17332 = s4 ? tmp17333 : tmp17337;
  assign tmp17342 = s2 ? tmp17112 : tmp16690;
  assign tmp17343 = s2 ? tmp16725 : tmp17101;
  assign tmp17341 = s3 ? tmp17342 : tmp17343;
  assign tmp17345 = s2 ? tmp17082 : tmp17078;
  assign tmp17346 = s2 ? tmp17101 : tmp17078;
  assign tmp17344 = s3 ? tmp17345 : tmp17346;
  assign tmp17340 = s4 ? tmp17341 : tmp17344;
  assign tmp17331 = s5 ? tmp17332 : tmp17340;
  assign tmp17329 = s6 ? tmp17330 : tmp17331;
  assign tmp17300 = s7 ? tmp17301 : tmp17329;
  assign tmp17299 = s8 ? tmp17259 : tmp17300;
  assign tmp17182 = s9 ? tmp17183 : tmp17299;
  assign tmp17356 = ~(s0 ? tmp17189 : tmp16690);
  assign tmp17355 = ~(s1 ? tmp17210 : tmp17356);
  assign tmp17354 = s2 ? tmp17208 : tmp17355;
  assign tmp17358 = s0 ? tmp16690 : tmp17189;
  assign tmp17357 = s2 ? tmp17358 : tmp17246;
  assign tmp17353 = s3 ? tmp17354 : tmp17357;
  assign tmp17352 = s4 ? tmp17353 : tmp17214;
  assign tmp17351 = s5 ? tmp17352 : tmp17220;
  assign tmp17350 = s6 ? tmp17186 : tmp17351;
  assign tmp17365 = s0 ? tmp17189 : tmp16690;
  assign tmp17364 = s1 ? tmp17189 : tmp17365;
  assign tmp17363 = s2 ? tmp17243 : tmp17364;
  assign tmp17362 = s3 ? tmp17363 : tmp17245;
  assign tmp17367 = s2 ? tmp17216 : tmp17189;
  assign tmp17366 = s3 ? tmp17367 : tmp17293;
  assign tmp17361 = s4 ? tmp17362 : tmp17366;
  assign tmp17360 = s5 ? tmp17361 : tmp17250;
  assign tmp17359 = s6 ? tmp17234 : tmp17360;
  assign tmp17349 = s7 ? tmp17350 : tmp17359;
  assign tmp17348 = s8 ? tmp17349 : tmp17350;
  assign tmp17373 = s3 ? tmp17248 : tmp17293;
  assign tmp17372 = s4 ? tmp17241 : tmp17373;
  assign tmp17375 = s3 ? tmp17256 : tmp17254;
  assign tmp17374 = s4 ? tmp17251 : tmp17375;
  assign tmp17371 = s5 ? tmp17372 : tmp17374;
  assign tmp17370 = s6 ? tmp17234 : tmp17371;
  assign tmp17379 = s3 ? tmp17345 : tmp17101;
  assign tmp17378 = s4 ? tmp17341 : tmp17379;
  assign tmp17377 = s5 ? tmp17332 : tmp17378;
  assign tmp17376 = s6 ? tmp17330 : tmp17377;
  assign tmp17369 = s7 ? tmp17370 : tmp17376;
  assign tmp17384 = s3 ? tmp17298 : tmp17254;
  assign tmp17383 = s4 ? tmp17295 : tmp17384;
  assign tmp17382 = s5 ? tmp17285 : tmp17383;
  assign tmp17381 = s6 ? tmp17283 : tmp17382;
  assign tmp17386 = s5 ? tmp17361 : tmp17374;
  assign tmp17385 = s6 ? tmp17234 : tmp17386;
  assign tmp17380 = s7 ? tmp17381 : tmp17385;
  assign tmp17368 = s8 ? tmp17369 : tmp17380;
  assign tmp17347 = s9 ? tmp17348 : tmp17368;
  assign tmp17181 = s10 ? tmp17182 : tmp17347;
  assign tmp17390 = s7 ? tmp17233 : tmp17329;
  assign tmp17391 = s7 ? tmp17282 : tmp17359;
  assign tmp17389 = s8 ? tmp17390 : tmp17391;
  assign tmp17388 = s9 ? tmp17348 : tmp17389;
  assign tmp17387 = s10 ? tmp17182 : tmp17388;
  assign tmp17180 = s11 ? tmp17181 : tmp17387;
  assign tmp17179 = s12 ? tmp17180 : 1;
  assign tmp17178 = s13 ? tmp17179 : 1;
  assign tmp17177 = ~(s14 ? 1 : tmp17178);
  assign tmp16677 = s15 ? tmp16678 : tmp17177;
  assign tmp17403 = s4 ? tmp16768 : tmp16747;
  assign tmp17402 = s5 ? tmp17403 : tmp16750;
  assign tmp17401 = s6 ? tmp16737 : tmp17402;
  assign tmp17400 = s7 ? tmp16757 : tmp17401;
  assign tmp17411 = l4 ? 1 : 0;
  assign tmp17410 = l2 ? tmp17411 : 1;
  assign tmp17409 = l1 ? 1 : tmp17410;
  assign tmp17413 = l1 ? 1 : tmp17411;
  assign tmp17412 = s0 ? tmp17413 : tmp17409;
  assign tmp17408 = s1 ? tmp17409 : tmp17412;
  assign tmp17416 = s0 ? tmp17409 : 1;
  assign tmp17415 = s1 ? tmp17416 : tmp17409;
  assign tmp17414 = s2 ? tmp17409 : tmp17415;
  assign tmp17407 = s3 ? tmp17408 : tmp17414;
  assign tmp17420 = s0 ? tmp17413 : 1;
  assign tmp17419 = s1 ? tmp17416 : tmp17420;
  assign tmp17418 = s2 ? tmp17415 : tmp17419;
  assign tmp17422 = s1 ? tmp17413 : tmp16703;
  assign tmp17424 = s0 ? tmp17411 : tmp17409;
  assign tmp17423 = s1 ? tmp17409 : tmp17424;
  assign tmp17421 = s2 ? tmp17422 : tmp17423;
  assign tmp17417 = s3 ? tmp17418 : tmp17421;
  assign tmp17406 = s4 ? tmp17407 : tmp17417;
  assign tmp17429 = s1 ? tmp17416 : 1;
  assign tmp17431 = s0 ? 1 : tmp17409;
  assign tmp17430 = s1 ? tmp17431 : tmp17416;
  assign tmp17428 = s2 ? tmp17429 : tmp17430;
  assign tmp17434 = s0 ? tmp17411 : 0;
  assign tmp17433 = s1 ? tmp17434 : tmp17409;
  assign tmp17432 = s2 ? tmp17431 : tmp17433;
  assign tmp17427 = s3 ? tmp17428 : tmp17432;
  assign tmp17439 = ~(l1 ? 1 : tmp17410);
  assign tmp17438 = s0 ? 1 : tmp17439;
  assign tmp17440 = ~(s0 ? 1 : tmp17413);
  assign tmp17437 = s1 ? tmp17438 : tmp17440;
  assign tmp17442 = s0 ? 1 : tmp17413;
  assign tmp17441 = ~(s1 ? tmp17442 : tmp17416);
  assign tmp17436 = s2 ? tmp17437 : tmp17441;
  assign tmp17445 = s0 ? tmp17413 : tmp16693;
  assign tmp17444 = s1 ? tmp17409 : tmp17445;
  assign tmp17443 = ~(s2 ? tmp17444 : 0);
  assign tmp17435 = ~(s3 ? tmp17436 : tmp17443);
  assign tmp17426 = s4 ? tmp17427 : tmp17435;
  assign tmp17450 = s0 ? tmp17409 : 0;
  assign tmp17451 = ~(s0 ? 1 : tmp17191);
  assign tmp17449 = s1 ? tmp17450 : tmp17451;
  assign tmp17453 = s0 ? tmp17411 : 1;
  assign tmp17452 = s1 ? tmp17453 : 1;
  assign tmp17448 = s2 ? tmp17449 : tmp17452;
  assign tmp17454 = s2 ? tmp16727 : tmp16729;
  assign tmp17447 = s3 ? tmp17448 : tmp17454;
  assign tmp17458 = s0 ? 1 : tmp17191;
  assign tmp17457 = s1 ? tmp16726 : tmp17458;
  assign tmp17459 = s1 ? tmp17438 : 0;
  assign tmp17456 = s2 ? tmp17457 : tmp17459;
  assign tmp17462 = ~(s0 ? 1 : tmp16690);
  assign tmp17461 = s1 ? tmp17434 : tmp17462;
  assign tmp17463 = ~(s1 ? tmp16705 : 1);
  assign tmp17460 = ~(s2 ? tmp17461 : tmp17463);
  assign tmp17455 = ~(s3 ? tmp17456 : tmp17460);
  assign tmp17446 = s4 ? tmp17447 : tmp17455;
  assign tmp17425 = s5 ? tmp17426 : tmp17446;
  assign tmp17405 = s6 ? tmp17406 : tmp17425;
  assign tmp17468 = s1 ? tmp17416 : tmp17413;
  assign tmp17467 = s2 ? tmp17415 : tmp17468;
  assign tmp17470 = s1 ? tmp17413 : 0;
  assign tmp17469 = s2 ? tmp17470 : tmp17423;
  assign tmp17466 = s3 ? tmp17467 : tmp17469;
  assign tmp17465 = s4 ? tmp17407 : tmp17466;
  assign tmp17475 = s1 ? tmp17409 : tmp17416;
  assign tmp17474 = s2 ? tmp17429 : tmp17475;
  assign tmp17476 = s2 ? tmp17409 : tmp17433;
  assign tmp17473 = s3 ? tmp17474 : tmp17476;
  assign tmp17479 = ~(s1 ? tmp17413 : tmp17409);
  assign tmp17478 = s2 ? tmp17437 : tmp17479;
  assign tmp17477 = ~(s3 ? tmp17478 : tmp17443);
  assign tmp17472 = s4 ? tmp17473 : tmp17477;
  assign tmp17483 = s1 ? tmp17450 : tmp17411;
  assign tmp17482 = s2 ? tmp17483 : 1;
  assign tmp17484 = ~(s2 ? 1 : tmp16714);
  assign tmp17481 = s3 ? tmp17482 : tmp17484;
  assign tmp17487 = s1 ? 1 : tmp17191;
  assign tmp17486 = s2 ? tmp17487 : tmp17439;
  assign tmp17485 = ~(s3 ? tmp17486 : tmp16714);
  assign tmp17480 = s4 ? tmp17481 : tmp17485;
  assign tmp17471 = s5 ? tmp17472 : tmp17480;
  assign tmp17464 = s6 ? tmp17465 : tmp17471;
  assign tmp17404 = ~(s7 ? tmp17405 : tmp17464);
  assign tmp17399 = s8 ? tmp17400 : tmp17404;
  assign tmp17489 = s7 ? tmp17405 : tmp17464;
  assign tmp17495 = s1 ? tmp17420 : tmp17413;
  assign tmp17494 = s2 ? tmp17495 : tmp17420;
  assign tmp17498 = s0 ? tmp17411 : tmp17413;
  assign tmp17497 = s1 ? tmp17413 : tmp17498;
  assign tmp17496 = s2 ? tmp17422 : tmp17497;
  assign tmp17493 = s3 ? tmp17494 : tmp17496;
  assign tmp17492 = s4 ? tmp17413 : tmp17493;
  assign tmp17503 = s1 ? tmp17420 : 1;
  assign tmp17504 = s1 ? tmp17442 : tmp17413;
  assign tmp17502 = s2 ? tmp17503 : tmp17504;
  assign tmp17506 = s1 ? tmp17434 : tmp17413;
  assign tmp17505 = s2 ? tmp17413 : tmp17506;
  assign tmp17501 = s3 ? tmp17502 : tmp17505;
  assign tmp17511 = ~(l1 ? 1 : tmp17411);
  assign tmp17510 = s0 ? 1 : tmp17511;
  assign tmp17509 = s1 ? tmp17510 : tmp17440;
  assign tmp17512 = ~(s1 ? tmp17442 : tmp17420);
  assign tmp17508 = s2 ? tmp17509 : tmp17512;
  assign tmp17515 = s0 ? tmp17413 : tmp16692;
  assign tmp17514 = s1 ? tmp17413 : tmp17515;
  assign tmp17513 = ~(s2 ? tmp17514 : 0);
  assign tmp17507 = ~(s3 ? tmp17508 : tmp17513);
  assign tmp17500 = s4 ? tmp17501 : tmp17507;
  assign tmp17520 = s0 ? tmp17413 : 0;
  assign tmp17519 = s1 ? tmp17520 : tmp17451;
  assign tmp17518 = s2 ? tmp17519 : tmp17452;
  assign tmp17517 = s3 ? tmp17518 : tmp16807;
  assign tmp17523 = s1 ? tmp16805 : tmp17451;
  assign tmp17524 = ~(s1 ? tmp17510 : 0);
  assign tmp17522 = s2 ? tmp17523 : tmp17524;
  assign tmp17526 = s1 ? tmp17434 : tmp16786;
  assign tmp17527 = ~(s1 ? tmp16799 : 1);
  assign tmp17525 = s2 ? tmp17526 : tmp17527;
  assign tmp17521 = s3 ? tmp17522 : tmp17525;
  assign tmp17516 = s4 ? tmp17517 : tmp17521;
  assign tmp17499 = s5 ? tmp17500 : tmp17516;
  assign tmp17491 = s6 ? tmp17492 : tmp17499;
  assign tmp17531 = s2 ? tmp17470 : tmp17497;
  assign tmp17530 = s3 ? tmp17495 : tmp17531;
  assign tmp17529 = s4 ? tmp17413 : tmp17530;
  assign tmp17535 = s2 ? tmp17503 : tmp17413;
  assign tmp17534 = s3 ? tmp17535 : tmp17505;
  assign tmp17537 = s2 ? tmp17509 : tmp17511;
  assign tmp17536 = ~(s3 ? tmp17537 : tmp17513);
  assign tmp17533 = s4 ? tmp17534 : tmp17536;
  assign tmp17541 = s1 ? tmp17520 : tmp17411;
  assign tmp17540 = s2 ? tmp17541 : 1;
  assign tmp17539 = s3 ? tmp17540 : tmp16826;
  assign tmp17543 = s2 ? tmp17487 : tmp17511;
  assign tmp17542 = ~(s3 ? tmp17543 : tmp16827);
  assign tmp17538 = s4 ? tmp17539 : tmp17542;
  assign tmp17532 = s5 ? tmp17533 : tmp17538;
  assign tmp17528 = s6 ? tmp17529 : tmp17532;
  assign tmp17490 = s7 ? tmp17491 : tmp17528;
  assign tmp17488 = ~(s8 ? tmp17489 : tmp17490);
  assign tmp17398 = s9 ? tmp17399 : tmp17488;
  assign tmp17545 = s8 ? tmp17489 : tmp17405;
  assign tmp17550 = s4 ? tmp16768 : tmp16841;
  assign tmp17549 = s5 ? tmp17550 : tmp16750;
  assign tmp17548 = s6 ? tmp16737 : tmp17549;
  assign tmp17556 = s1 ? tmp17413 : tmp16692;
  assign tmp17555 = ~(s2 ? tmp17556 : 0);
  assign tmp17554 = ~(s3 ? tmp17537 : tmp17555);
  assign tmp17553 = s4 ? tmp17534 : tmp17554;
  assign tmp17552 = s5 ? tmp17553 : tmp17538;
  assign tmp17551 = ~(s6 ? tmp17529 : tmp17552);
  assign tmp17547 = s7 ? tmp17548 : tmp17551;
  assign tmp17562 = s1 ? tmp17409 : tmp16693;
  assign tmp17561 = ~(s2 ? tmp17562 : 0);
  assign tmp17560 = ~(s3 ? tmp17478 : tmp17561);
  assign tmp17559 = s4 ? tmp17473 : tmp17560;
  assign tmp17558 = s5 ? tmp17559 : tmp17480;
  assign tmp17557 = ~(s6 ? tmp17465 : tmp17558);
  assign tmp17546 = ~(s8 ? tmp17547 : tmp17557);
  assign tmp17544 = ~(s9 ? tmp17545 : tmp17546);
  assign tmp17397 = s10 ? tmp17398 : tmp17544;
  assign tmp17567 = ~(s6 ? tmp17529 : tmp17532);
  assign tmp17566 = s7 ? tmp17401 : tmp17567;
  assign tmp17568 = ~(s6 ? tmp17465 : tmp17471);
  assign tmp17565 = ~(s8 ? tmp17566 : tmp17568);
  assign tmp17564 = ~(s9 ? tmp17545 : tmp17565);
  assign tmp17563 = s10 ? tmp17398 : tmp17564;
  assign tmp17396 = ~(s11 ? tmp17397 : tmp17563);
  assign tmp17395 = s12 ? 1 : tmp17396;
  assign tmp17578 = l1 ? tmp16690 : tmp16693;
  assign tmp17580 = ~(l1 ? tmp16690 : tmp16693);
  assign tmp17579 = ~(s0 ? 1 : tmp17580);
  assign tmp17577 = s1 ? tmp17578 : tmp17579;
  assign tmp17583 = s0 ? tmp17578 : 0;
  assign tmp17582 = s1 ? tmp17583 : tmp17578;
  assign tmp17581 = s2 ? tmp17578 : tmp17582;
  assign tmp17576 = s3 ? tmp17577 : tmp17581;
  assign tmp17586 = s1 ? tmp17583 : 0;
  assign tmp17585 = s2 ? tmp17582 : tmp17586;
  assign tmp17589 = s0 ? 1 : tmp17578;
  assign tmp17588 = ~(s1 ? tmp17578 : tmp17589);
  assign tmp17587 = ~(s2 ? tmp16868 : tmp17588);
  assign tmp17584 = s3 ? tmp17585 : tmp17587;
  assign tmp17575 = s4 ? tmp17576 : tmp17584;
  assign tmp17594 = s1 ? tmp17583 : tmp17579;
  assign tmp17596 = s0 ? 1 : tmp17580;
  assign tmp17597 = ~(s0 ? tmp17578 : 0);
  assign tmp17595 = ~(s1 ? tmp17596 : tmp17597);
  assign tmp17593 = s2 ? tmp17594 : tmp17595;
  assign tmp17599 = ~(s1 ? 1 : tmp17578);
  assign tmp17598 = ~(s2 ? tmp17596 : tmp17599);
  assign tmp17592 = s3 ? tmp17593 : tmp17598;
  assign tmp17602 = s1 ? tmp17589 : 0;
  assign tmp17603 = ~(s1 ? 1 : tmp17597);
  assign tmp17601 = s2 ? tmp17602 : tmp17603;
  assign tmp17605 = s1 ? tmp17578 : tmp16887;
  assign tmp17604 = s2 ? tmp17605 : 1;
  assign tmp17600 = s3 ? tmp17601 : tmp17604;
  assign tmp17591 = s4 ? tmp17592 : tmp17600;
  assign tmp17611 = l1 ? 1 : tmp16693;
  assign tmp17610 = s0 ? tmp17578 : tmp17611;
  assign tmp17609 = s1 ? tmp17610 : 1;
  assign tmp17612 = s1 ? tmp17589 : tmp17578;
  assign tmp17608 = s2 ? tmp17609 : tmp17612;
  assign tmp17607 = s3 ? tmp17608 : tmp16893;
  assign tmp17616 = s0 ? tmp17611 : tmp17578;
  assign tmp17615 = s1 ? tmp17616 : tmp17578;
  assign tmp17614 = s2 ? tmp16690 : tmp17615;
  assign tmp17613 = s3 ? tmp17614 : tmp16733;
  assign tmp17606 = s4 ? tmp17607 : tmp17613;
  assign tmp17590 = s5 ? tmp17591 : tmp17606;
  assign tmp17574 = s6 ? tmp17575 : tmp17590;
  assign tmp17620 = ~(s2 ? tmp16901 : tmp17588);
  assign tmp17619 = s3 ? tmp17585 : tmp17620;
  assign tmp17618 = s4 ? tmp17576 : tmp17619;
  assign tmp17625 = s1 ? tmp17578 : tmp17583;
  assign tmp17624 = s2 ? tmp17582 : tmp17625;
  assign tmp17627 = s1 ? 1 : tmp17578;
  assign tmp17626 = s2 ? tmp17578 : tmp17627;
  assign tmp17623 = s3 ? tmp17624 : tmp17626;
  assign tmp17629 = s2 ? tmp17602 : tmp17578;
  assign tmp17631 = s1 ? tmp17578 : tmp16690;
  assign tmp17630 = s2 ? tmp17631 : 1;
  assign tmp17628 = s3 ? tmp17629 : tmp17630;
  assign tmp17622 = s4 ? tmp17623 : tmp17628;
  assign tmp17634 = s2 ? tmp17609 : tmp17631;
  assign tmp17633 = s3 ? tmp17634 : tmp16753;
  assign tmp17636 = s2 ? 1 : tmp17578;
  assign tmp17635 = s3 ? tmp17636 : tmp16690;
  assign tmp17632 = s4 ? tmp17633 : tmp17635;
  assign tmp17621 = s5 ? tmp17622 : tmp17632;
  assign tmp17617 = s6 ? tmp17618 : tmp17621;
  assign tmp17573 = s7 ? tmp17574 : tmp17617;
  assign tmp17643 = s1 ? tmp17578 : tmp16691;
  assign tmp17642 = s2 ? tmp17643 : 1;
  assign tmp17641 = s3 ? tmp17601 : tmp17642;
  assign tmp17640 = s4 ? tmp17592 : tmp17641;
  assign tmp17646 = s2 ? tmp16971 : tmp17615;
  assign tmp17645 = s3 ? tmp17646 : tmp16733;
  assign tmp17644 = s4 ? tmp17607 : tmp17645;
  assign tmp17639 = s5 ? tmp17640 : tmp17644;
  assign tmp17638 = s6 ? tmp17575 : tmp17639;
  assign tmp17637 = s7 ? tmp17638 : tmp17617;
  assign tmp17572 = s8 ? tmp17573 : tmp17637;
  assign tmp17652 = ~(s2 ? tmp16868 : tmp16860);
  assign tmp17651 = s3 ? tmp16865 : tmp17652;
  assign tmp17650 = s4 ? tmp16856 : tmp17651;
  assign tmp17657 = ~(s1 ? tmp16781 : tmp16858);
  assign tmp17656 = ~(s2 ? tmp16877 : tmp17657);
  assign tmp17655 = s3 ? tmp16874 : tmp17656;
  assign tmp17654 = s4 ? tmp17655 : tmp16881;
  assign tmp17662 = s0 ? tmp16858 : tmp16692;
  assign tmp17661 = s1 ? tmp17662 : tmp16692;
  assign tmp17660 = s2 ? tmp17661 : tmp16858;
  assign tmp17659 = s3 ? tmp17660 : tmp16893;
  assign tmp17665 = s1 ? tmp16690 : tmp16692;
  assign tmp17667 = s0 ? tmp16692 : tmp16858;
  assign tmp17666 = s1 ? tmp17667 : tmp16858;
  assign tmp17664 = s2 ? tmp17665 : tmp17666;
  assign tmp17669 = s1 ? tmp16692 : tmp16705;
  assign tmp17668 = s2 ? tmp17669 : tmp16735;
  assign tmp17663 = s3 ? tmp17664 : tmp17668;
  assign tmp17658 = s4 ? tmp17659 : tmp17663;
  assign tmp17653 = s5 ? tmp17654 : tmp17658;
  assign tmp17649 = s6 ? tmp17650 : tmp17653;
  assign tmp17673 = ~(s2 ? tmp16901 : tmp16860);
  assign tmp17672 = s3 ? tmp16865 : tmp17673;
  assign tmp17671 = s4 ? tmp16856 : tmp17672;
  assign tmp17678 = s1 ? tmp16781 : tmp16858;
  assign tmp17677 = s2 ? tmp16858 : tmp17678;
  assign tmp17676 = s3 ? tmp16905 : tmp17677;
  assign tmp17675 = s4 ? tmp17676 : tmp16909;
  assign tmp17680 = s3 ? tmp17660 : tmp17013;
  assign tmp17682 = s2 ? tmp16692 : tmp16858;
  assign tmp17681 = s3 ? tmp17682 : tmp16690;
  assign tmp17679 = s4 ? tmp17680 : tmp17681;
  assign tmp17674 = s5 ? tmp17675 : tmp17679;
  assign tmp17670 = s6 ? tmp17671 : tmp17674;
  assign tmp17648 = s7 ? tmp17649 : tmp17670;
  assign tmp17647 = s8 ? tmp17637 : tmp17648;
  assign tmp17571 = s9 ? tmp17572 : tmp17647;
  assign tmp17691 = s0 ? tmp16692 : tmp17578;
  assign tmp17690 = ~(s1 ? tmp17578 : tmp17691);
  assign tmp17689 = ~(s2 ? tmp16868 : tmp17690);
  assign tmp17688 = s3 ? tmp17585 : tmp17689;
  assign tmp17687 = s4 ? tmp17576 : tmp17688;
  assign tmp17696 = ~(s1 ? tmp16781 : tmp17578);
  assign tmp17695 = ~(s2 ? tmp17596 : tmp17696);
  assign tmp17694 = s3 ? tmp17593 : tmp17695;
  assign tmp17693 = s4 ? tmp17694 : tmp17600;
  assign tmp17700 = s1 ? tmp17610 : tmp16692;
  assign tmp17701 = s1 ? tmp17691 : tmp17578;
  assign tmp17699 = s2 ? tmp17700 : tmp17701;
  assign tmp17698 = s3 ? tmp17699 : tmp16893;
  assign tmp17703 = s2 ? tmp17665 : tmp17615;
  assign tmp17702 = s3 ? tmp17703 : tmp17668;
  assign tmp17697 = s4 ? tmp17698 : tmp17702;
  assign tmp17692 = s5 ? tmp17693 : tmp17697;
  assign tmp17686 = s6 ? tmp17687 : tmp17692;
  assign tmp17707 = ~(s2 ? tmp16901 : tmp17690);
  assign tmp17706 = s3 ? tmp17585 : tmp17707;
  assign tmp17705 = s4 ? tmp17576 : tmp17706;
  assign tmp17712 = s1 ? tmp16781 : tmp17578;
  assign tmp17711 = s2 ? tmp17578 : tmp17712;
  assign tmp17710 = s3 ? tmp17624 : tmp17711;
  assign tmp17709 = s4 ? tmp17710 : tmp17628;
  assign tmp17715 = s2 ? tmp17700 : tmp17631;
  assign tmp17714 = s3 ? tmp17715 : tmp16753;
  assign tmp17717 = s2 ? tmp16692 : tmp17578;
  assign tmp17716 = s3 ? tmp17717 : tmp16690;
  assign tmp17713 = s4 ? tmp17714 : tmp17716;
  assign tmp17708 = s5 ? tmp17709 : tmp17713;
  assign tmp17704 = s6 ? tmp17705 : tmp17708;
  assign tmp17685 = s7 ? tmp17686 : tmp17704;
  assign tmp17684 = s8 ? tmp17685 : tmp17686;
  assign tmp17719 = s7 ? tmp17617 : tmp17670;
  assign tmp17718 = s8 ? tmp17719 : tmp17704;
  assign tmp17683 = s9 ? tmp17684 : tmp17718;
  assign tmp17570 = s10 ? tmp17571 : tmp17683;
  assign tmp17728 = s3 ? tmp17056 : tmp16753;
  assign tmp17727 = s4 ? tmp17728 : tmp17164;
  assign tmp17726 = s5 ? tmp17065 : tmp17727;
  assign tmp17725 = s6 ? tmp17061 : tmp17726;
  assign tmp17724 = s7 ? tmp17038 : tmp17725;
  assign tmp17733 = s3 ? tmp17137 : tmp16753;
  assign tmp17732 = s4 ? tmp17733 : tmp17169;
  assign tmp17731 = s5 ? tmp17126 : tmp17732;
  assign tmp17730 = s6 ? tmp17120 : tmp17731;
  assign tmp17729 = s7 ? tmp17074 : tmp17730;
  assign tmp17723 = s8 ? tmp17724 : tmp17729;
  assign tmp17734 = s8 ? tmp17729 : tmp17142;
  assign tmp17722 = s9 ? tmp17723 : tmp17734;
  assign tmp17739 = s5 ? tmp17150 : tmp17727;
  assign tmp17738 = s6 ? tmp17061 : tmp17739;
  assign tmp17737 = s7 ? tmp17143 : tmp17738;
  assign tmp17736 = s8 ? tmp17737 : tmp17143;
  assign tmp17744 = s4 ? tmp17154 : tmp17164;
  assign tmp17743 = s5 ? tmp17150 : tmp17744;
  assign tmp17742 = s6 ? tmp17061 : tmp17743;
  assign tmp17741 = s7 ? tmp17725 : tmp17742;
  assign tmp17745 = s7 ? tmp17730 : tmp17738;
  assign tmp17740 = s8 ? tmp17741 : tmp17745;
  assign tmp17735 = s9 ? tmp17736 : tmp17740;
  assign tmp17721 = s10 ? tmp17722 : tmp17735;
  assign tmp17749 = s7 ? tmp17725 : tmp17148;
  assign tmp17748 = s8 ? tmp17749 : tmp17745;
  assign tmp17747 = s9 ? tmp17736 : tmp17748;
  assign tmp17746 = s10 ? tmp17722 : tmp17747;
  assign tmp17720 = s11 ? tmp17721 : tmp17746;
  assign tmp17569 = ~(s12 ? tmp17570 : tmp17720);
  assign tmp17394 = s13 ? tmp17395 : tmp17569;
  assign tmp17393 = s14 ? 1 : tmp17394;
  assign tmp17764 = ~(s0 ? tmp17189 : tmp16718);
  assign tmp17763 = ~(s1 ? tmp17210 : tmp17764);
  assign tmp17762 = s2 ? tmp17208 : tmp17763;
  assign tmp17766 = s0 ? tmp16692 : tmp17193;
  assign tmp17765 = ~(s2 ? tmp17766 : tmp17213);
  assign tmp17761 = s3 ? tmp17762 : tmp17765;
  assign tmp17760 = s4 ? tmp17761 : tmp17214;
  assign tmp17759 = s5 ? tmp17760 : tmp17220;
  assign tmp17758 = s6 ? tmp17186 : tmp17759;
  assign tmp17773 = s0 ? tmp17189 : tmp16718;
  assign tmp17772 = s1 ? tmp17189 : tmp17773;
  assign tmp17771 = s2 ? tmp17243 : tmp17772;
  assign tmp17770 = s3 ? tmp17771 : tmp17245;
  assign tmp17769 = s4 ? tmp17770 : tmp17247;
  assign tmp17776 = s2 ? 1 : tmp17254;
  assign tmp17775 = s3 ? tmp17252 : tmp17776;
  assign tmp17778 = s2 ? tmp17101 : tmp17189;
  assign tmp17777 = s3 ? tmp17778 : tmp17254;
  assign tmp17774 = s4 ? tmp17775 : tmp17777;
  assign tmp17768 = s5 ? tmp17769 : tmp17774;
  assign tmp17767 = s6 ? tmp17234 : tmp17768;
  assign tmp17757 = s7 ? tmp17758 : tmp17767;
  assign tmp17784 = s1 ? tmp17203 : tmp17189;
  assign tmp17783 = s2 ? tmp17784 : tmp17246;
  assign tmp17782 = s3 ? tmp17188 : tmp17783;
  assign tmp17781 = s4 ? tmp17782 : tmp17196;
  assign tmp17780 = s6 ? tmp17781 : tmp17263;
  assign tmp17786 = s4 ? tmp17782 : tmp17235;
  assign tmp17789 = s3 ? tmp17296 : tmp17776;
  assign tmp17791 = s2 ? 1 : tmp17189;
  assign tmp17790 = s3 ? tmp17791 : tmp17254;
  assign tmp17788 = s4 ? tmp17789 : tmp17790;
  assign tmp17787 = s5 ? tmp17285 : tmp17788;
  assign tmp17785 = s6 ? tmp17786 : tmp17787;
  assign tmp17779 = s7 ? tmp17780 : tmp17785;
  assign tmp17756 = s8 ? tmp17757 : tmp17779;
  assign tmp17798 = s2 ? tmp17309 : tmp17096;
  assign tmp17799 = s2 ? tmp17100 : tmp17082;
  assign tmp17797 = s3 ? tmp17798 : tmp17799;
  assign tmp17796 = s4 ? tmp17797 : tmp17313;
  assign tmp17795 = s5 ? tmp17796 : tmp17318;
  assign tmp17794 = s6 ? tmp17302 : tmp17795;
  assign tmp17804 = s2 ? tmp17335 : tmp17129;
  assign tmp17803 = s3 ? tmp17804 : tmp17081;
  assign tmp17802 = s4 ? tmp17803 : tmp17337;
  assign tmp17801 = s5 ? tmp17802 : tmp17340;
  assign tmp17800 = s6 ? tmp17330 : tmp17801;
  assign tmp17793 = s7 ? tmp17794 : tmp17800;
  assign tmp17792 = s8 ? tmp17779 : tmp17793;
  assign tmp17755 = s9 ? tmp17756 : tmp17792;
  assign tmp17812 = s2 ? tmp17208 : tmp17268;
  assign tmp17813 = s2 ? tmp17217 : tmp17246;
  assign tmp17811 = s3 ? tmp17812 : tmp17813;
  assign tmp17810 = s4 ? tmp17811 : tmp17214;
  assign tmp17809 = s5 ? tmp17810 : tmp17220;
  assign tmp17808 = s6 ? tmp17186 : tmp17809;
  assign tmp17818 = s2 ? tmp17243 : tmp17289;
  assign tmp17817 = s3 ? tmp17818 : tmp17245;
  assign tmp17816 = s4 ? tmp17817 : tmp17366;
  assign tmp17815 = s5 ? tmp17816 : tmp17774;
  assign tmp17814 = s6 ? tmp17234 : tmp17815;
  assign tmp17807 = s7 ? tmp17808 : tmp17814;
  assign tmp17806 = s8 ? tmp17807 : tmp17808;
  assign tmp17823 = s4 ? tmp17770 : tmp17373;
  assign tmp17822 = s5 ? tmp17823 : tmp17774;
  assign tmp17821 = s6 ? tmp17234 : tmp17822;
  assign tmp17825 = s5 ? tmp17802 : tmp17378;
  assign tmp17824 = s6 ? tmp17330 : tmp17825;
  assign tmp17820 = s7 ? tmp17821 : tmp17824;
  assign tmp17826 = s7 ? tmp17785 : tmp17814;
  assign tmp17819 = s8 ? tmp17820 : tmp17826;
  assign tmp17805 = s9 ? tmp17806 : tmp17819;
  assign tmp17754 = s10 ? tmp17755 : tmp17805;
  assign tmp17830 = s7 ? tmp17767 : tmp17800;
  assign tmp17829 = s8 ? tmp17830 : tmp17826;
  assign tmp17828 = s9 ? tmp17806 : tmp17829;
  assign tmp17827 = s10 ? tmp17755 : tmp17828;
  assign tmp17753 = s11 ? tmp17754 : tmp17827;
  assign tmp17840 = s1 ? tmp16793 : 1;
  assign tmp17839 = s2 ? tmp17840 : 1;
  assign tmp17838 = s3 ? tmp17839 : 1;
  assign tmp17837 = s4 ? 1 : tmp17838;
  assign tmp17846 = s0 ? 1 : tmp17611;
  assign tmp17845 = s1 ? tmp17846 : 1;
  assign tmp17848 = s0 ? tmp17611 : 1;
  assign tmp17847 = s1 ? tmp17848 : 1;
  assign tmp17844 = s2 ? tmp17845 : tmp17847;
  assign tmp17843 = s3 ? tmp17844 : 1;
  assign tmp17851 = s1 ? 1 : tmp16781;
  assign tmp17852 = s1 ? tmp16781 : tmp16793;
  assign tmp17850 = s2 ? tmp17851 : tmp17852;
  assign tmp17849 = s3 ? tmp17850 : 1;
  assign tmp17842 = s4 ? tmp17843 : tmp17849;
  assign tmp17841 = s5 ? tmp17842 : 1;
  assign tmp17836 = s6 ? tmp17837 : tmp17841;
  assign tmp17857 = s2 ? tmp17845 : 1;
  assign tmp17856 = s3 ? tmp17857 : 1;
  assign tmp17859 = s2 ? tmp17851 : 1;
  assign tmp17858 = s3 ? tmp17859 : 1;
  assign tmp17855 = s4 ? tmp17856 : tmp17858;
  assign tmp17854 = s5 ? tmp17855 : 1;
  assign tmp17853 = s6 ? tmp17837 : tmp17854;
  assign tmp17835 = s7 ? tmp17836 : tmp17853;
  assign tmp17865 = ~(l2 ? tmp17411 : 0);
  assign tmp17864 = l1 ? 1 : tmp17865;
  assign tmp17868 = s0 ? 1 : tmp17864;
  assign tmp17867 = s1 ? tmp17868 : tmp17864;
  assign tmp17866 = s2 ? tmp17867 : tmp17864;
  assign tmp17863 = s3 ? tmp17864 : tmp17866;
  assign tmp17872 = s0 ? tmp17864 : 0;
  assign tmp17871 = s1 ? tmp17872 : tmp17864;
  assign tmp17873 = s0 ? tmp17864 : 1;
  assign tmp17870 = s2 ? tmp17871 : tmp17873;
  assign tmp17875 = s1 ? tmp17411 : 0;
  assign tmp17876 = ~(l1 ? 1 : tmp17865);
  assign tmp17874 = ~(s2 ? tmp17875 : tmp17876);
  assign tmp17869 = s3 ? tmp17870 : tmp17874;
  assign tmp17862 = s4 ? tmp17863 : tmp17869;
  assign tmp17882 = s0 ? tmp17864 : tmp17611;
  assign tmp17881 = s1 ? tmp17882 : 1;
  assign tmp17884 = s0 ? tmp17611 : tmp17864;
  assign tmp17883 = s1 ? tmp17884 : tmp17864;
  assign tmp17880 = s2 ? tmp17881 : tmp17883;
  assign tmp17888 = l1 ? 1 : tmp17191;
  assign tmp17887 = s0 ? tmp17888 : 1;
  assign tmp17886 = s1 ? tmp17887 : tmp17864;
  assign tmp17885 = s2 ? tmp17864 : tmp17886;
  assign tmp17879 = s3 ? tmp17880 : tmp17885;
  assign tmp17892 = ~(s0 ? 1 : tmp17411);
  assign tmp17891 = s1 ? tmp17868 : tmp17892;
  assign tmp17894 = s0 ? 1 : tmp17411;
  assign tmp17895 = ~(s0 ? tmp17864 : 0);
  assign tmp17893 = ~(s1 ? tmp17894 : tmp17895);
  assign tmp17890 = s2 ? tmp17891 : tmp17893;
  assign tmp17898 = ~(s0 ? tmp17411 : 0);
  assign tmp17897 = s1 ? tmp17864 : tmp17898;
  assign tmp17896 = s2 ? tmp17897 : 1;
  assign tmp17889 = s3 ? tmp17890 : tmp17896;
  assign tmp17878 = s4 ? tmp17879 : tmp17889;
  assign tmp17903 = s0 ? 1 : tmp17888;
  assign tmp17902 = s1 ? tmp17873 : tmp17903;
  assign tmp17904 = s1 ? tmp17887 : 1;
  assign tmp17901 = s2 ? tmp17902 : tmp17904;
  assign tmp17900 = s3 ? tmp17901 : 1;
  assign tmp17907 = s1 ? 1 : tmp17903;
  assign tmp17908 = s1 ? tmp17868 : 1;
  assign tmp17906 = s2 ? tmp17907 : tmp17908;
  assign tmp17909 = s2 ? tmp17904 : 1;
  assign tmp17905 = s3 ? tmp17906 : tmp17909;
  assign tmp17899 = s4 ? tmp17900 : tmp17905;
  assign tmp17877 = s5 ? tmp17878 : tmp17899;
  assign tmp17861 = s6 ? tmp17862 : tmp17877;
  assign tmp17914 = s2 ? tmp17881 : tmp17864;
  assign tmp17913 = s3 ? tmp17914 : tmp17885;
  assign tmp17916 = s2 ? tmp17891 : tmp17864;
  assign tmp17918 = s1 ? tmp17864 : 1;
  assign tmp17917 = s2 ? tmp17918 : 1;
  assign tmp17915 = s3 ? tmp17916 : tmp17917;
  assign tmp17912 = s4 ? tmp17913 : tmp17915;
  assign tmp17922 = s1 ? tmp17873 : tmp17888;
  assign tmp17921 = s2 ? tmp17922 : tmp17904;
  assign tmp17920 = s3 ? tmp17921 : 1;
  assign tmp17925 = s1 ? 1 : tmp17888;
  assign tmp17924 = s2 ? tmp17925 : tmp17864;
  assign tmp17923 = s3 ? tmp17924 : tmp17904;
  assign tmp17919 = s4 ? tmp17920 : tmp17923;
  assign tmp17911 = s5 ? tmp17912 : tmp17919;
  assign tmp17910 = s6 ? tmp17862 : tmp17911;
  assign tmp17860 = s7 ? tmp17861 : tmp17910;
  assign tmp17834 = s8 ? tmp17835 : tmp17860;
  assign tmp17932 = s1 ? tmp17882 : tmp17864;
  assign tmp17931 = s2 ? tmp17932 : tmp17873;
  assign tmp17930 = s3 ? tmp17931 : tmp17874;
  assign tmp17929 = s4 ? tmp17863 : tmp17930;
  assign tmp17938 = ~(s0 ? tmp17864 : tmp17611);
  assign tmp17937 = ~(s1 ? tmp17894 : tmp17938);
  assign tmp17936 = s2 ? tmp17891 : tmp17937;
  assign tmp17935 = s3 ? tmp17936 : tmp17896;
  assign tmp17934 = s4 ? tmp17879 : tmp17935;
  assign tmp17933 = s5 ? tmp17934 : tmp17899;
  assign tmp17928 = s6 ? tmp17929 : tmp17933;
  assign tmp17939 = s6 ? tmp17929 : tmp17911;
  assign tmp17927 = s7 ? tmp17928 : tmp17939;
  assign tmp17946 = s0 ? tmp17888 : tmp16692;
  assign tmp17945 = s1 ? tmp17946 : tmp17888;
  assign tmp17944 = s2 ? tmp17945 : tmp17887;
  assign tmp17948 = ~(l1 ? 1 : tmp17191);
  assign tmp17947 = ~(s2 ? tmp17875 : tmp17948);
  assign tmp17943 = s3 ? tmp17944 : tmp17947;
  assign tmp17942 = s4 ? tmp17888 : tmp17943;
  assign tmp17953 = s1 ? tmp17946 : tmp16692;
  assign tmp17955 = s0 ? tmp16692 : tmp17888;
  assign tmp17954 = s1 ? tmp17955 : tmp17888;
  assign tmp17952 = s2 ? tmp17953 : tmp17954;
  assign tmp17957 = s1 ? tmp17887 : tmp17888;
  assign tmp17956 = s2 ? tmp17888 : tmp17957;
  assign tmp17951 = s3 ? tmp17952 : tmp17956;
  assign tmp17960 = s1 ? tmp17903 : tmp17892;
  assign tmp17962 = ~(s0 ? tmp17888 : tmp16692);
  assign tmp17961 = ~(s1 ? tmp17894 : tmp17962);
  assign tmp17959 = s2 ? tmp17960 : tmp17961;
  assign tmp17964 = s1 ? tmp17888 : tmp17898;
  assign tmp17963 = s2 ? tmp17964 : 1;
  assign tmp17958 = s3 ? tmp17959 : tmp17963;
  assign tmp17950 = s4 ? tmp17951 : tmp17958;
  assign tmp17968 = s1 ? tmp17887 : tmp17903;
  assign tmp17969 = s1 ? tmp17888 : tmp16793;
  assign tmp17967 = s2 ? tmp17968 : tmp17969;
  assign tmp17966 = s3 ? tmp17967 : 1;
  assign tmp17972 = s1 ? tmp17903 : tmp16781;
  assign tmp17971 = s2 ? tmp17907 : tmp17972;
  assign tmp17970 = s3 ? tmp17971 : tmp17909;
  assign tmp17965 = s4 ? tmp17966 : tmp17970;
  assign tmp17949 = s5 ? tmp17950 : tmp17965;
  assign tmp17941 = s6 ? tmp17942 : tmp17949;
  assign tmp17977 = s2 ? tmp17953 : tmp17888;
  assign tmp17976 = s3 ? tmp17977 : tmp17956;
  assign tmp17979 = s2 ? tmp17960 : tmp17888;
  assign tmp17981 = s1 ? tmp17888 : 1;
  assign tmp17980 = s2 ? tmp17981 : 1;
  assign tmp17978 = s3 ? tmp17979 : tmp17980;
  assign tmp17975 = s4 ? tmp17976 : tmp17978;
  assign tmp17984 = s2 ? tmp17957 : tmp17981;
  assign tmp17983 = s3 ? tmp17984 : 1;
  assign tmp17986 = s2 ? tmp17925 : tmp17888;
  assign tmp17985 = s3 ? tmp17986 : tmp17904;
  assign tmp17982 = s4 ? tmp17983 : tmp17985;
  assign tmp17974 = s5 ? tmp17975 : tmp17982;
  assign tmp17973 = s6 ? tmp17942 : tmp17974;
  assign tmp17940 = s7 ? tmp17941 : tmp17973;
  assign tmp17926 = s8 ? tmp17927 : tmp17940;
  assign tmp17833 = s9 ? tmp17834 : tmp17926;
  assign tmp17991 = s4 ? tmp17864 : tmp17930;
  assign tmp17996 = s1 ? tmp17882 : tmp17611;
  assign tmp17995 = s2 ? tmp17996 : tmp17883;
  assign tmp17994 = s3 ? tmp17995 : tmp17885;
  assign tmp17993 = s4 ? tmp17994 : tmp17935;
  assign tmp18000 = s1 ? tmp17864 : tmp17846;
  assign tmp17999 = s2 ? tmp17902 : tmp18000;
  assign tmp17998 = s3 ? tmp17999 : 1;
  assign tmp18003 = s1 ? tmp17868 : tmp17848;
  assign tmp18002 = s2 ? tmp17907 : tmp18003;
  assign tmp18001 = s3 ? tmp18002 : tmp17909;
  assign tmp17997 = s4 ? tmp17998 : tmp18001;
  assign tmp17992 = s5 ? tmp17993 : tmp17997;
  assign tmp17990 = s6 ? tmp17991 : tmp17992;
  assign tmp18008 = s2 ? tmp17996 : tmp17864;
  assign tmp18007 = s3 ? tmp18008 : tmp17885;
  assign tmp18006 = s4 ? tmp18007 : tmp17915;
  assign tmp18011 = s2 ? tmp17922 : tmp17918;
  assign tmp18010 = s3 ? tmp18011 : 1;
  assign tmp18009 = s4 ? tmp18010 : tmp17923;
  assign tmp18005 = s5 ? tmp18006 : tmp18009;
  assign tmp18004 = s6 ? tmp17991 : tmp18005;
  assign tmp17989 = s7 ? tmp17990 : tmp18004;
  assign tmp17988 = s8 ? tmp17989 : tmp17990;
  assign tmp18017 = s3 ? tmp17986 : 1;
  assign tmp18016 = s4 ? tmp17983 : tmp18017;
  assign tmp18015 = s5 ? tmp17975 : tmp18016;
  assign tmp18014 = s6 ? tmp17942 : tmp18015;
  assign tmp18013 = s7 ? tmp17853 : tmp18014;
  assign tmp18021 = s3 ? tmp17924 : 1;
  assign tmp18020 = s4 ? tmp18010 : tmp18021;
  assign tmp18019 = s5 ? tmp18006 : tmp18020;
  assign tmp18018 = s6 ? tmp17991 : tmp18019;
  assign tmp18012 = s8 ? tmp18013 : tmp18018;
  assign tmp17987 = s9 ? tmp17988 : tmp18012;
  assign tmp17832 = s10 ? tmp17833 : tmp17987;
  assign tmp18025 = s7 ? tmp17853 : tmp17973;
  assign tmp18024 = s8 ? tmp18025 : tmp18004;
  assign tmp18023 = s9 ? tmp17988 : tmp18024;
  assign tmp18022 = s10 ? tmp17833 : tmp18023;
  assign tmp17831 = s11 ? tmp17832 : tmp18022;
  assign tmp17752 = s12 ? tmp17753 : tmp17831;
  assign tmp17751 = s13 ? tmp17752 : 1;
  assign tmp17750 = ~(s14 ? 1 : tmp17751);
  assign tmp17392 = s15 ? tmp17393 : tmp17750;
  assign tmp16676 = s16 ? tmp16677 : tmp17392;
  assign tmp18041 = s1 ? tmp16793 : tmp16781;
  assign tmp18040 = s2 ? tmp16791 : tmp18041;
  assign tmp18042 = s2 ? tmp16793 : tmp16795;
  assign tmp18039 = s3 ? tmp18040 : tmp18042;
  assign tmp18038 = s4 ? tmp18039 : tmp16796;
  assign tmp18037 = s5 ? tmp18038 : tmp16801;
  assign tmp18036 = s6 ? tmp16777 : tmp18037;
  assign tmp18048 = s1 ? tmp16692 : tmp16781;
  assign tmp18047 = s2 ? tmp16791 : tmp18048;
  assign tmp18046 = s3 ? tmp18047 : tmp16794;
  assign tmp18045 = s4 ? tmp18046 : tmp16796;
  assign tmp18044 = s5 ? tmp18045 : tmp16823;
  assign tmp18043 = s6 ? tmp16816 : tmp18044;
  assign tmp18035 = s7 ? tmp18036 : tmp18043;
  assign tmp18034 = ~(s8 ? tmp17489 : tmp18035);
  assign tmp18033 = s9 ? tmp17399 : tmp18034;
  assign tmp18050 = s8 ? tmp16756 : tmp16757;
  assign tmp18053 = ~(s6 ? tmp16816 : tmp18044);
  assign tmp18052 = s7 ? tmp17548 : tmp18053;
  assign tmp18055 = s6 ? tmp17465 : tmp17558;
  assign tmp18056 = ~(s6 ? tmp16737 : tmp16766);
  assign tmp18054 = ~(s7 ? tmp18055 : tmp18056);
  assign tmp18051 = s8 ? tmp18052 : tmp18054;
  assign tmp18049 = s9 ? tmp18050 : tmp18051;
  assign tmp18032 = s10 ? tmp18033 : tmp18049;
  assign tmp18060 = s7 ? tmp17401 : tmp18053;
  assign tmp18061 = ~(s7 ? tmp17464 : tmp18056);
  assign tmp18059 = s8 ? tmp18060 : tmp18061;
  assign tmp18058 = s9 ? tmp18050 : tmp18059;
  assign tmp18057 = s10 ? tmp18033 : tmp18058;
  assign tmp18031 = ~(s11 ? tmp18032 : tmp18057);
  assign tmp18030 = s12 ? 1 : tmp18031;
  assign tmp18072 = s1 ? tmp17667 : 0;
  assign tmp18071 = s2 ? tmp18072 : tmp16884;
  assign tmp18070 = s3 ? tmp18071 : tmp16885;
  assign tmp18069 = s4 ? tmp16873 : tmp18070;
  assign tmp18076 = s1 ? tmp17662 : 1;
  assign tmp18075 = s2 ? tmp18076 : tmp16858;
  assign tmp18074 = s3 ? tmp18075 : tmp16893;
  assign tmp18078 = s2 ? tmp16690 : tmp17666;
  assign tmp18077 = s3 ? tmp18078 : tmp16733;
  assign tmp18073 = s4 ? tmp18074 : tmp18077;
  assign tmp18068 = s5 ? tmp18069 : tmp18073;
  assign tmp18067 = s6 ? tmp16855 : tmp18068;
  assign tmp18083 = s2 ? tmp18072 : tmp16858;
  assign tmp18082 = s3 ? tmp18083 : tmp16911;
  assign tmp18081 = s4 ? tmp16904 : tmp18082;
  assign tmp18085 = s3 ? tmp18075 : tmp16915;
  assign tmp18084 = s4 ? tmp18085 : tmp16916;
  assign tmp18080 = s5 ? tmp18081 : tmp18084;
  assign tmp18079 = s6 ? tmp16898 : tmp18080;
  assign tmp18066 = s7 ? tmp18067 : tmp18079;
  assign tmp18092 = s1 ? tmp16858 : tmp16691;
  assign tmp18091 = s2 ? tmp18092 : 1;
  assign tmp18090 = s3 ? tmp18071 : tmp18091;
  assign tmp18089 = s4 ? tmp16873 : tmp18090;
  assign tmp18095 = s2 ? tmp18076 : tmp16896;
  assign tmp18094 = s3 ? tmp18095 : tmp16893;
  assign tmp18097 = s2 ? tmp16971 : tmp17666;
  assign tmp18096 = s3 ? tmp18097 : tmp16733;
  assign tmp18093 = s4 ? tmp18094 : tmp18096;
  assign tmp18088 = s5 ? tmp18089 : tmp18093;
  assign tmp18087 = s6 ? tmp16855 : tmp18088;
  assign tmp18086 = s7 ? tmp18087 : tmp18079;
  assign tmp18065 = s8 ? tmp18066 : tmp18086;
  assign tmp18104 = s2 ? tmp18076 : tmp17006;
  assign tmp18103 = s3 ? tmp18104 : tmp16893;
  assign tmp18102 = s4 ? tmp18103 : tmp18077;
  assign tmp18101 = s5 ? tmp18069 : tmp18102;
  assign tmp18100 = s6 ? tmp16855 : tmp18101;
  assign tmp18109 = s2 ? tmp18076 : tmp16912;
  assign tmp18108 = s3 ? tmp18109 : tmp17013;
  assign tmp18107 = s4 ? tmp18108 : tmp16916;
  assign tmp18106 = s5 ? tmp18081 : tmp18107;
  assign tmp18105 = s6 ? tmp16898 : tmp18106;
  assign tmp18099 = s7 ? tmp18100 : tmp18105;
  assign tmp18098 = s8 ? tmp18086 : tmp18099;
  assign tmp18064 = s9 ? tmp18065 : tmp18098;
  assign tmp18116 = s3 ? tmp18109 : tmp16915;
  assign tmp18115 = s4 ? tmp18116 : tmp16916;
  assign tmp18114 = s5 ? tmp18081 : tmp18115;
  assign tmp18113 = s6 ? tmp16898 : tmp18114;
  assign tmp18112 = s7 ? tmp18067 : tmp18113;
  assign tmp18111 = s8 ? tmp18112 : tmp18067;
  assign tmp18117 = s7 ? tmp18079 : tmp18113;
  assign tmp18110 = s9 ? tmp18111 : tmp18117;
  assign tmp18063 = s10 ? tmp18064 : tmp18110;
  assign tmp18062 = ~(s12 ? tmp18063 : tmp17033);
  assign tmp18029 = s13 ? tmp18030 : tmp18062;
  assign tmp18028 = s14 ? 1 : tmp18029;
  assign tmp18130 = s2 ? tmp17840 : tmp16791;
  assign tmp18129 = s3 ? tmp18130 : 1;
  assign tmp18128 = s4 ? tmp18129 : tmp17849;
  assign tmp18127 = s5 ? tmp18128 : 1;
  assign tmp18126 = s6 ? tmp17837 : tmp18127;
  assign tmp18133 = s4 ? tmp17838 : tmp17858;
  assign tmp18132 = s5 ? tmp18133 : 1;
  assign tmp18131 = s6 ? tmp17837 : tmp18132;
  assign tmp18125 = s7 ? tmp18126 : tmp18131;
  assign tmp18124 = s8 ? tmp17927 : tmp18125;
  assign tmp18123 = s9 ? tmp17834 : tmp18124;
  assign tmp18138 = s4 ? 1 : tmp17856;
  assign tmp18143 = s1 ? tmp16781 : tmp17846;
  assign tmp18142 = s2 ? tmp17851 : tmp18143;
  assign tmp18141 = s3 ? tmp18142 : 1;
  assign tmp18140 = s4 ? tmp17843 : tmp18141;
  assign tmp18139 = s5 ? tmp18140 : 1;
  assign tmp18137 = s6 ? tmp18138 : tmp18139;
  assign tmp18144 = s6 ? tmp18138 : tmp17854;
  assign tmp18136 = s7 ? tmp18137 : tmp18144;
  assign tmp18135 = s8 ? tmp18136 : tmp18137;
  assign tmp18146 = s7 ? tmp17853 : tmp18131;
  assign tmp18150 = s4 ? tmp17920 : tmp18021;
  assign tmp18149 = s5 ? tmp17912 : tmp18150;
  assign tmp18148 = s6 ? tmp17929 : tmp18149;
  assign tmp18147 = s7 ? tmp18148 : tmp18144;
  assign tmp18145 = s8 ? tmp18146 : tmp18147;
  assign tmp18134 = s9 ? tmp18135 : tmp18145;
  assign tmp18122 = s10 ? tmp18123 : tmp18134;
  assign tmp18154 = s7 ? tmp17939 : tmp18144;
  assign tmp18153 = s8 ? tmp18146 : tmp18154;
  assign tmp18152 = s9 ? tmp18135 : tmp18153;
  assign tmp18151 = s10 ? tmp18123 : tmp18152;
  assign tmp18121 = s11 ? tmp18122 : tmp18151;
  assign tmp18120 = s12 ? tmp17180 : tmp18121;
  assign tmp18119 = s13 ? tmp18120 : 1;
  assign tmp18118 = ~(s14 ? 1 : tmp18119);
  assign tmp18027 = s15 ? tmp18028 : tmp18118;
  assign tmp18167 = ~(s1 ? tmp16858 : tmp17667);
  assign tmp18166 = ~(s2 ? tmp16868 : tmp18167);
  assign tmp18165 = s3 ? tmp16865 : tmp18166;
  assign tmp18164 = s4 ? tmp16856 : tmp18165;
  assign tmp18169 = s4 ? tmp17655 : tmp18070;
  assign tmp18173 = s1 ? tmp16690 : tmp16858;
  assign tmp18172 = s2 ? tmp18173 : tmp17666;
  assign tmp18171 = s3 ? tmp18172 : tmp17668;
  assign tmp18170 = s4 ? tmp17659 : tmp18171;
  assign tmp18168 = s5 ? tmp18169 : tmp18170;
  assign tmp18163 = s6 ? tmp18164 : tmp18168;
  assign tmp18177 = ~(s2 ? tmp16901 : tmp18167);
  assign tmp18176 = s3 ? tmp16865 : tmp18177;
  assign tmp18175 = s4 ? tmp16856 : tmp18176;
  assign tmp18179 = s4 ? tmp17676 : tmp18082;
  assign tmp18181 = s3 ? tmp17660 : tmp16915;
  assign tmp18180 = s4 ? tmp18181 : tmp17681;
  assign tmp18178 = s5 ? tmp18179 : tmp18180;
  assign tmp18174 = s6 ? tmp18175 : tmp18178;
  assign tmp18162 = s7 ? tmp18163 : tmp18174;
  assign tmp18187 = s2 ? tmp17661 : tmp17666;
  assign tmp18186 = s3 ? tmp18187 : tmp16893;
  assign tmp18185 = s4 ? tmp18186 : tmp17663;
  assign tmp18184 = s5 ? tmp18169 : tmp18185;
  assign tmp18183 = s6 ? tmp18164 : tmp18184;
  assign tmp18182 = s7 ? tmp18183 : tmp18174;
  assign tmp18161 = s8 ? tmp18162 : tmp18182;
  assign tmp18160 = s9 ? tmp18161 : tmp18182;
  assign tmp18189 = s8 ? tmp18182 : tmp18183;
  assign tmp18188 = s9 ? tmp18189 : tmp18174;
  assign tmp18159 = s10 ? tmp18160 : tmp18188;
  assign tmp18158 = ~(s12 ? tmp18159 : tmp17033);
  assign tmp18157 = s13 ? tmp17395 : tmp18158;
  assign tmp18156 = s14 ? 1 : tmp18157;
  assign tmp18192 = s12 ? tmp17180 : tmp17831;
  assign tmp18191 = s13 ? tmp18192 : 1;
  assign tmp18190 = ~(s14 ? 1 : tmp18191);
  assign tmp18155 = s15 ? tmp18156 : tmp18190;
  assign tmp18026 = s16 ? tmp18027 : tmp18155;
  assign tmp16675 = s17 ? tmp16676 : tmp18026;
  assign s15n = tmp16675;

  assign tmp18208 = l3 ? 1 : 0;
  assign tmp18209 = l2 ? 1 : 0;
  assign tmp18207 = l1 ? tmp18208 : tmp18209;
  assign tmp18211 = l1 ? tmp18208 : 1;
  assign tmp18210 = s0 ? tmp18211 : tmp18207;
  assign tmp18206 = s1 ? tmp18207 : tmp18210;
  assign tmp18214 = s0 ? tmp18207 : 1;
  assign tmp18213 = s1 ? tmp18214 : tmp18207;
  assign tmp18212 = s2 ? tmp18207 : tmp18213;
  assign tmp18205 = s3 ? tmp18206 : tmp18212;
  assign tmp18218 = s0 ? tmp18207 : tmp18211;
  assign tmp18217 = s1 ? tmp18218 : tmp18207;
  assign tmp18220 = s0 ? tmp18211 : 1;
  assign tmp18219 = s1 ? tmp18214 : tmp18220;
  assign tmp18216 = s2 ? tmp18217 : tmp18219;
  assign tmp18223 = s0 ? 1 : 0;
  assign tmp18222 = s1 ? tmp18211 : tmp18223;
  assign tmp18225 = s0 ? tmp18207 : tmp18209;
  assign tmp18227 = ~(l1 ? tmp18208 : tmp18209);
  assign tmp18226 = ~(s0 ? 1 : tmp18227);
  assign tmp18224 = s1 ? tmp18225 : tmp18226;
  assign tmp18221 = s2 ? tmp18222 : tmp18224;
  assign tmp18215 = s3 ? tmp18216 : tmp18221;
  assign tmp18204 = s4 ? tmp18205 : tmp18215;
  assign tmp18233 = s0 ? 1 : tmp18207;
  assign tmp18232 = s1 ? tmp18214 : tmp18233;
  assign tmp18235 = s0 ? tmp18209 : 1;
  assign tmp18234 = s1 ? tmp18233 : tmp18235;
  assign tmp18231 = s2 ? tmp18232 : tmp18234;
  assign tmp18237 = s0 ? 1 : tmp18209;
  assign tmp18239 = ~(s0 ? tmp18207 : 0);
  assign tmp18238 = ~(s1 ? 1 : tmp18239);
  assign tmp18236 = s2 ? tmp18237 : tmp18238;
  assign tmp18230 = s3 ? tmp18231 : tmp18236;
  assign tmp18243 = s0 ? 1 : tmp18227;
  assign tmp18244 = ~(s0 ? tmp18211 : 0);
  assign tmp18242 = s1 ? tmp18243 : tmp18244;
  assign tmp18246 = s0 ? tmp18211 : 0;
  assign tmp18245 = ~(s1 ? tmp18246 : tmp18218);
  assign tmp18241 = s2 ? tmp18242 : tmp18245;
  assign tmp18248 = s1 ? tmp18209 : 0;
  assign tmp18247 = ~(s2 ? tmp18248 : 0);
  assign tmp18240 = ~(s3 ? tmp18241 : tmp18247);
  assign tmp18229 = s4 ? tmp18230 : tmp18240;
  assign tmp18253 = s0 ? tmp18209 : 0;
  assign tmp18252 = s1 ? tmp18253 : 0;
  assign tmp18256 = ~(l2 ? 1 : 0);
  assign tmp18255 = s0 ? 1 : tmp18256;
  assign tmp18254 = ~(s1 ? tmp18255 : tmp18256);
  assign tmp18251 = s2 ? tmp18252 : tmp18254;
  assign tmp18250 = s3 ? tmp18251 : 0;
  assign tmp18259 = s1 ? tmp18255 : tmp18256;
  assign tmp18258 = s2 ? 1 : tmp18259;
  assign tmp18257 = ~(s3 ? tmp18258 : 1);
  assign tmp18249 = s4 ? tmp18250 : tmp18257;
  assign tmp18228 = s5 ? tmp18229 : tmp18249;
  assign tmp18203 = s6 ? tmp18204 : tmp18228;
  assign tmp18264 = s1 ? tmp18214 : tmp18211;
  assign tmp18263 = s2 ? tmp18217 : tmp18264;
  assign tmp18266 = s1 ? tmp18211 : 0;
  assign tmp18265 = s2 ? tmp18266 : tmp18224;
  assign tmp18262 = s3 ? tmp18263 : tmp18265;
  assign tmp18261 = s4 ? tmp18205 : tmp18262;
  assign tmp18271 = s1 ? tmp18207 : tmp18235;
  assign tmp18270 = s2 ? tmp18213 : tmp18271;
  assign tmp18272 = s2 ? tmp18209 : tmp18238;
  assign tmp18269 = s3 ? tmp18270 : tmp18272;
  assign tmp18275 = ~(s1 ? tmp18211 : tmp18218);
  assign tmp18274 = s2 ? tmp18242 : tmp18275;
  assign tmp18273 = ~(s3 ? tmp18274 : tmp18247);
  assign tmp18268 = s4 ? tmp18269 : tmp18273;
  assign tmp18278 = s2 ? tmp18252 : tmp18248;
  assign tmp18277 = s3 ? tmp18278 : 0;
  assign tmp18280 = s2 ? 1 : tmp18256;
  assign tmp18279 = ~(s3 ? tmp18280 : 1);
  assign tmp18276 = s4 ? tmp18277 : tmp18279;
  assign tmp18267 = s5 ? tmp18268 : tmp18276;
  assign tmp18260 = s6 ? tmp18261 : tmp18267;
  assign tmp18202 = s7 ? tmp18203 : tmp18260;
  assign tmp18287 = l2 ? 1 : tmp18208;
  assign tmp18286 = l1 ? tmp18287 : tmp18209;
  assign tmp18289 = l1 ? tmp18287 : 1;
  assign tmp18288 = s0 ? tmp18289 : tmp18286;
  assign tmp18285 = s1 ? tmp18286 : tmp18288;
  assign tmp18292 = s0 ? tmp18286 : 1;
  assign tmp18291 = s1 ? tmp18292 : tmp18286;
  assign tmp18290 = s2 ? tmp18286 : tmp18291;
  assign tmp18284 = s3 ? tmp18285 : tmp18290;
  assign tmp18296 = s0 ? tmp18286 : tmp18289;
  assign tmp18295 = s1 ? tmp18296 : tmp18286;
  assign tmp18298 = s0 ? tmp18289 : 1;
  assign tmp18297 = s1 ? tmp18292 : tmp18298;
  assign tmp18294 = s2 ? tmp18295 : tmp18297;
  assign tmp18300 = s1 ? tmp18289 : tmp18223;
  assign tmp18302 = s0 ? tmp18286 : tmp18209;
  assign tmp18304 = ~(l1 ? tmp18287 : tmp18209);
  assign tmp18303 = ~(s0 ? 1 : tmp18304);
  assign tmp18301 = s1 ? tmp18302 : tmp18303;
  assign tmp18299 = s2 ? tmp18300 : tmp18301;
  assign tmp18293 = s3 ? tmp18294 : tmp18299;
  assign tmp18283 = s4 ? tmp18284 : tmp18293;
  assign tmp18310 = s0 ? 1 : tmp18286;
  assign tmp18309 = s1 ? tmp18292 : tmp18310;
  assign tmp18311 = s1 ? tmp18310 : tmp18235;
  assign tmp18308 = s2 ? tmp18309 : tmp18311;
  assign tmp18315 = l1 ? tmp18209 : 0;
  assign tmp18314 = ~(s0 ? tmp18286 : tmp18315);
  assign tmp18313 = ~(s1 ? 1 : tmp18314);
  assign tmp18312 = s2 ? tmp18237 : tmp18313;
  assign tmp18307 = s3 ? tmp18308 : tmp18312;
  assign tmp18319 = s0 ? 1 : tmp18304;
  assign tmp18320 = ~(s0 ? tmp18289 : tmp18209);
  assign tmp18318 = s1 ? tmp18319 : tmp18320;
  assign tmp18322 = s0 ? tmp18289 : tmp18209;
  assign tmp18321 = ~(s1 ? tmp18322 : tmp18296);
  assign tmp18317 = s2 ? tmp18318 : tmp18321;
  assign tmp18325 = s0 ? tmp18209 : tmp18315;
  assign tmp18324 = s1 ? tmp18325 : tmp18253;
  assign tmp18323 = ~(s2 ? tmp18324 : 0);
  assign tmp18316 = ~(s3 ? tmp18317 : tmp18323);
  assign tmp18306 = s4 ? tmp18307 : tmp18316;
  assign tmp18305 = s5 ? tmp18306 : tmp18249;
  assign tmp18282 = s6 ? tmp18283 : tmp18305;
  assign tmp18330 = s1 ? tmp18292 : tmp18289;
  assign tmp18329 = s2 ? tmp18295 : tmp18330;
  assign tmp18332 = s1 ? tmp18289 : 0;
  assign tmp18331 = s2 ? tmp18332 : tmp18301;
  assign tmp18328 = s3 ? tmp18329 : tmp18331;
  assign tmp18327 = s4 ? tmp18284 : tmp18328;
  assign tmp18337 = s1 ? tmp18286 : tmp18235;
  assign tmp18336 = s2 ? tmp18291 : tmp18337;
  assign tmp18338 = s2 ? tmp18209 : tmp18313;
  assign tmp18335 = s3 ? tmp18336 : tmp18338;
  assign tmp18340 = s2 ? tmp18318 : tmp18304;
  assign tmp18342 = s1 ? tmp18325 : 0;
  assign tmp18341 = ~(s2 ? tmp18342 : 0);
  assign tmp18339 = ~(s3 ? tmp18340 : tmp18341);
  assign tmp18334 = s4 ? tmp18335 : tmp18339;
  assign tmp18333 = s5 ? tmp18334 : tmp18276;
  assign tmp18326 = s6 ? tmp18327 : tmp18333;
  assign tmp18281 = s7 ? tmp18282 : tmp18326;
  assign tmp18201 = s8 ? tmp18202 : tmp18281;
  assign tmp18348 = s2 ? tmp18211 : tmp18220;
  assign tmp18352 = ~(l1 ? 1 : 0);
  assign tmp18351 = s0 ? tmp18211 : tmp18352;
  assign tmp18354 = ~(l1 ? tmp18208 : 1);
  assign tmp18353 = ~(s0 ? 1 : tmp18354);
  assign tmp18350 = s1 ? tmp18351 : tmp18353;
  assign tmp18349 = s2 ? tmp18222 : tmp18350;
  assign tmp18347 = s3 ? tmp18348 : tmp18349;
  assign tmp18346 = s4 ? tmp18211 : tmp18347;
  assign tmp18361 = l1 ? 1 : 0;
  assign tmp18360 = ~(s0 ? tmp18361 : 0);
  assign tmp18359 = s1 ? tmp18211 : tmp18360;
  assign tmp18358 = s2 ? tmp18211 : tmp18359;
  assign tmp18363 = s0 ? 1 : tmp18352;
  assign tmp18364 = ~(s1 ? 1 : tmp18244);
  assign tmp18362 = s2 ? tmp18363 : tmp18364;
  assign tmp18357 = s3 ? tmp18358 : tmp18362;
  assign tmp18368 = s0 ? 1 : tmp18354;
  assign tmp18367 = s1 ? tmp18368 : tmp18244;
  assign tmp18369 = ~(s1 ? tmp18246 : tmp18211);
  assign tmp18366 = s2 ? tmp18367 : tmp18369;
  assign tmp18370 = s2 ? tmp18361 : 1;
  assign tmp18365 = ~(s3 ? tmp18366 : tmp18370);
  assign tmp18356 = s4 ? tmp18357 : tmp18365;
  assign tmp18375 = s0 ? tmp18361 : 1;
  assign tmp18374 = s1 ? tmp18375 : 1;
  assign tmp18377 = s0 ? 1 : tmp18361;
  assign tmp18376 = s1 ? tmp18377 : tmp18361;
  assign tmp18373 = s2 ? tmp18374 : tmp18376;
  assign tmp18372 = s3 ? tmp18373 : 1;
  assign tmp18379 = s2 ? 1 : tmp18376;
  assign tmp18378 = s3 ? tmp18379 : 1;
  assign tmp18371 = ~(s4 ? tmp18372 : tmp18378);
  assign tmp18355 = s5 ? tmp18356 : tmp18371;
  assign tmp18345 = s6 ? tmp18346 : tmp18355;
  assign tmp18384 = s1 ? tmp18220 : tmp18211;
  assign tmp18383 = s2 ? tmp18211 : tmp18384;
  assign tmp18385 = s2 ? tmp18266 : tmp18350;
  assign tmp18382 = s3 ? tmp18383 : tmp18385;
  assign tmp18381 = s4 ? tmp18211 : tmp18382;
  assign tmp18390 = s1 ? 1 : tmp18244;
  assign tmp18389 = ~(s2 ? tmp18361 : tmp18390);
  assign tmp18388 = s3 ? tmp18358 : tmp18389;
  assign tmp18392 = s2 ? tmp18367 : tmp18354;
  assign tmp18394 = s1 ? tmp18361 : 1;
  assign tmp18393 = s2 ? tmp18394 : 1;
  assign tmp18391 = ~(s3 ? tmp18392 : tmp18393);
  assign tmp18387 = s4 ? tmp18388 : tmp18391;
  assign tmp18397 = s2 ? tmp18374 : tmp18394;
  assign tmp18396 = s3 ? tmp18397 : 1;
  assign tmp18399 = s2 ? 1 : tmp18361;
  assign tmp18398 = s3 ? tmp18399 : 1;
  assign tmp18395 = ~(s4 ? tmp18396 : tmp18398);
  assign tmp18386 = s5 ? tmp18387 : tmp18395;
  assign tmp18380 = s6 ? tmp18381 : tmp18386;
  assign tmp18344 = s7 ? tmp18345 : tmp18380;
  assign tmp18343 = s8 ? tmp18281 : tmp18344;
  assign tmp18200 = s9 ? tmp18201 : tmp18343;
  assign tmp18407 = s2 ? tmp18242 : tmp18227;
  assign tmp18406 = ~(s3 ? tmp18407 : tmp18247);
  assign tmp18405 = s4 ? tmp18269 : tmp18406;
  assign tmp18404 = s5 ? tmp18405 : tmp18276;
  assign tmp18403 = s6 ? tmp18261 : tmp18404;
  assign tmp18402 = s7 ? tmp18203 : tmp18403;
  assign tmp18401 = s8 ? tmp18402 : tmp18203;
  assign tmp18415 = ~(s1 ? tmp18211 : tmp18207);
  assign tmp18414 = s2 ? tmp18242 : tmp18415;
  assign tmp18413 = ~(s3 ? tmp18414 : tmp18247);
  assign tmp18412 = s4 ? tmp18269 : tmp18413;
  assign tmp18411 = s5 ? tmp18412 : tmp18276;
  assign tmp18410 = s6 ? tmp18261 : tmp18411;
  assign tmp18409 = s7 ? tmp18410 : tmp18380;
  assign tmp18416 = s7 ? tmp18326 : tmp18403;
  assign tmp18408 = s8 ? tmp18409 : tmp18416;
  assign tmp18400 = s9 ? tmp18401 : tmp18408;
  assign tmp18199 = s10 ? tmp18200 : tmp18400;
  assign tmp18420 = s7 ? tmp18260 : tmp18380;
  assign tmp18419 = s8 ? tmp18420 : tmp18416;
  assign tmp18418 = s9 ? tmp18401 : tmp18419;
  assign tmp18417 = s10 ? tmp18200 : tmp18418;
  assign tmp18198 = s11 ? tmp18199 : tmp18417;
  assign tmp18197 = s13 ? tmp18198 : 1;
  assign tmp18422 = s12 ? 1 : 0;
  assign tmp18433 = l1 ? 1 : tmp18256;
  assign tmp18434 = s0 ? tmp18361 : tmp18433;
  assign tmp18432 = s1 ? tmp18433 : tmp18434;
  assign tmp18437 = s0 ? tmp18433 : 0;
  assign tmp18436 = s1 ? tmp18437 : tmp18433;
  assign tmp18435 = s2 ? tmp18433 : tmp18436;
  assign tmp18431 = s3 ? tmp18432 : tmp18435;
  assign tmp18441 = s0 ? tmp18433 : tmp18361;
  assign tmp18440 = s1 ? tmp18441 : tmp18433;
  assign tmp18443 = s0 ? tmp18361 : 0;
  assign tmp18442 = s1 ? tmp18437 : tmp18443;
  assign tmp18439 = s2 ? tmp18440 : tmp18442;
  assign tmp18446 = ~(s0 ? 1 : 0);
  assign tmp18445 = s1 ? tmp18361 : tmp18446;
  assign tmp18448 = s0 ? 1 : tmp18433;
  assign tmp18447 = s1 ? tmp18433 : tmp18448;
  assign tmp18444 = s2 ? tmp18445 : tmp18447;
  assign tmp18438 = s3 ? tmp18439 : tmp18444;
  assign tmp18430 = s4 ? tmp18431 : tmp18438;
  assign tmp18455 = ~(l1 ? 1 : tmp18256);
  assign tmp18454 = ~(s0 ? 1 : tmp18455);
  assign tmp18453 = s1 ? tmp18437 : tmp18454;
  assign tmp18457 = s0 ? 1 : tmp18455;
  assign tmp18458 = ~(s0 ? tmp18433 : 0);
  assign tmp18456 = ~(s1 ? tmp18457 : tmp18458);
  assign tmp18452 = s2 ? tmp18453 : tmp18456;
  assign tmp18461 = s0 ? tmp18433 : 1;
  assign tmp18460 = ~(s1 ? 1 : tmp18461);
  assign tmp18459 = ~(s2 ? tmp18457 : tmp18460);
  assign tmp18451 = s3 ? tmp18452 : tmp18459;
  assign tmp18464 = s1 ? tmp18448 : tmp18375;
  assign tmp18465 = s1 ? tmp18375 : tmp18441;
  assign tmp18463 = s2 ? tmp18464 : tmp18465;
  assign tmp18467 = s1 ? tmp18461 : 1;
  assign tmp18466 = s2 ? tmp18467 : 1;
  assign tmp18462 = s3 ? tmp18463 : tmp18466;
  assign tmp18450 = s4 ? tmp18451 : tmp18462;
  assign tmp18470 = s2 ? tmp18467 : tmp18448;
  assign tmp18469 = s3 ? tmp18470 : 1;
  assign tmp18473 = s1 ? tmp18448 : tmp18461;
  assign tmp18472 = s2 ? 1 : tmp18473;
  assign tmp18471 = s3 ? tmp18472 : 1;
  assign tmp18468 = s4 ? tmp18469 : tmp18471;
  assign tmp18449 = s5 ? tmp18450 : tmp18468;
  assign tmp18429 = s6 ? tmp18430 : tmp18449;
  assign tmp18478 = s1 ? tmp18437 : tmp18361;
  assign tmp18477 = s2 ? tmp18440 : tmp18478;
  assign tmp18479 = s2 ? tmp18394 : tmp18447;
  assign tmp18476 = s3 ? tmp18477 : tmp18479;
  assign tmp18475 = s4 ? tmp18431 : tmp18476;
  assign tmp18484 = s1 ? tmp18433 : tmp18437;
  assign tmp18483 = s2 ? tmp18436 : tmp18484;
  assign tmp18486 = s1 ? 1 : tmp18461;
  assign tmp18485 = s2 ? tmp18433 : tmp18486;
  assign tmp18482 = s3 ? tmp18483 : tmp18485;
  assign tmp18488 = s2 ? tmp18464 : tmp18433;
  assign tmp18487 = s3 ? tmp18488 : tmp18466;
  assign tmp18481 = s4 ? tmp18482 : tmp18487;
  assign tmp18492 = s1 ? tmp18433 : tmp18461;
  assign tmp18491 = s2 ? 1 : tmp18492;
  assign tmp18490 = s3 ? tmp18491 : 1;
  assign tmp18489 = s4 ? tmp18469 : tmp18490;
  assign tmp18480 = s5 ? tmp18481 : tmp18489;
  assign tmp18474 = s6 ? tmp18475 : tmp18480;
  assign tmp18428 = s7 ? tmp18429 : tmp18474;
  assign tmp18498 = ~(l3 ? 1 : 0);
  assign tmp18497 = l1 ? 1 : tmp18498;
  assign tmp18501 = s0 ? tmp18497 : tmp18498;
  assign tmp18500 = s1 ? tmp18501 : tmp18497;
  assign tmp18499 = s2 ? tmp18497 : tmp18500;
  assign tmp18496 = s3 ? tmp18497 : tmp18499;
  assign tmp18505 = s0 ? tmp18497 : tmp18361;
  assign tmp18504 = s1 ? tmp18505 : tmp18497;
  assign tmp18506 = s0 ? tmp18497 : 0;
  assign tmp18503 = s2 ? tmp18504 : tmp18506;
  assign tmp18508 = s1 ? tmp18497 : tmp18446;
  assign tmp18510 = s0 ? 1 : tmp18497;
  assign tmp18509 = s1 ? tmp18497 : tmp18510;
  assign tmp18507 = s2 ? tmp18508 : tmp18509;
  assign tmp18502 = s3 ? tmp18503 : tmp18507;
  assign tmp18495 = s4 ? tmp18496 : tmp18502;
  assign tmp18517 = ~(l1 ? 1 : tmp18498);
  assign tmp18516 = ~(s0 ? 1 : tmp18517);
  assign tmp18515 = s1 ? tmp18506 : tmp18516;
  assign tmp18519 = s0 ? 1 : tmp18517;
  assign tmp18520 = ~(s0 ? tmp18497 : tmp18498);
  assign tmp18518 = ~(s1 ? tmp18519 : tmp18520);
  assign tmp18514 = s2 ? tmp18515 : tmp18518;
  assign tmp18522 = s0 ? tmp18208 : tmp18517;
  assign tmp18523 = ~(s1 ? 1 : tmp18497);
  assign tmp18521 = ~(s2 ? tmp18522 : tmp18523);
  assign tmp18513 = s3 ? tmp18514 : tmp18521;
  assign tmp18526 = s1 ? tmp18510 : tmp18375;
  assign tmp18527 = s1 ? tmp18375 : tmp18505;
  assign tmp18525 = s2 ? tmp18526 : tmp18527;
  assign tmp18529 = s1 ? tmp18497 : 1;
  assign tmp18528 = s2 ? tmp18529 : 1;
  assign tmp18524 = s3 ? tmp18525 : tmp18528;
  assign tmp18512 = s4 ? tmp18513 : tmp18524;
  assign tmp18534 = s0 ? tmp18497 : 1;
  assign tmp18533 = s1 ? tmp18534 : 1;
  assign tmp18532 = s2 ? tmp18533 : tmp18510;
  assign tmp18531 = s3 ? tmp18532 : 1;
  assign tmp18537 = s1 ? tmp18510 : tmp18534;
  assign tmp18536 = s2 ? 1 : tmp18537;
  assign tmp18535 = s3 ? tmp18536 : 1;
  assign tmp18530 = s4 ? tmp18531 : tmp18535;
  assign tmp18511 = s5 ? tmp18512 : tmp18530;
  assign tmp18494 = s6 ? tmp18495 : tmp18511;
  assign tmp18542 = s1 ? tmp18506 : tmp18497;
  assign tmp18541 = s2 ? tmp18504 : tmp18542;
  assign tmp18543 = s2 ? tmp18529 : tmp18509;
  assign tmp18540 = s3 ? tmp18541 : tmp18543;
  assign tmp18539 = s4 ? tmp18496 : tmp18540;
  assign tmp18548 = s1 ? tmp18497 : tmp18501;
  assign tmp18547 = s2 ? tmp18542 : tmp18548;
  assign tmp18550 = s1 ? 1 : tmp18497;
  assign tmp18549 = s2 ? tmp18497 : tmp18550;
  assign tmp18546 = s3 ? tmp18547 : tmp18549;
  assign tmp18552 = s2 ? tmp18526 : tmp18497;
  assign tmp18551 = s3 ? tmp18552 : tmp18528;
  assign tmp18545 = s4 ? tmp18546 : tmp18551;
  assign tmp18555 = s2 ? tmp18533 : tmp18529;
  assign tmp18554 = s3 ? tmp18555 : 1;
  assign tmp18557 = s2 ? 1 : tmp18529;
  assign tmp18556 = s3 ? tmp18557 : 1;
  assign tmp18553 = s4 ? tmp18554 : tmp18556;
  assign tmp18544 = s5 ? tmp18545 : tmp18553;
  assign tmp18538 = s6 ? tmp18539 : tmp18544;
  assign tmp18493 = s7 ? tmp18494 : tmp18538;
  assign tmp18427 = s8 ? tmp18428 : tmp18493;
  assign tmp18564 = s1 ? tmp18443 : tmp18361;
  assign tmp18563 = s2 ? tmp18361 : tmp18564;
  assign tmp18562 = s3 ? tmp18361 : tmp18563;
  assign tmp18566 = s2 ? tmp18361 : tmp18443;
  assign tmp18568 = s1 ? tmp18361 : tmp18377;
  assign tmp18567 = s2 ? tmp18445 : tmp18568;
  assign tmp18565 = s3 ? tmp18566 : tmp18567;
  assign tmp18561 = s4 ? tmp18562 : tmp18565;
  assign tmp18574 = ~(s0 ? 1 : tmp18352);
  assign tmp18573 = s1 ? tmp18443 : tmp18574;
  assign tmp18575 = ~(s1 ? tmp18363 : tmp18360);
  assign tmp18572 = s2 ? tmp18573 : tmp18575;
  assign tmp18577 = ~(s1 ? 1 : tmp18434);
  assign tmp18576 = ~(s2 ? tmp18363 : tmp18577);
  assign tmp18571 = s3 ? tmp18572 : tmp18576;
  assign tmp18580 = s1 ? tmp18377 : tmp18375;
  assign tmp18581 = s1 ? tmp18375 : tmp18361;
  assign tmp18579 = s2 ? tmp18580 : tmp18581;
  assign tmp18583 = s1 ? tmp18434 : 1;
  assign tmp18582 = s2 ? tmp18583 : 1;
  assign tmp18578 = s3 ? tmp18579 : tmp18582;
  assign tmp18570 = s4 ? tmp18571 : tmp18578;
  assign tmp18587 = s1 ? tmp18377 : tmp18441;
  assign tmp18586 = s2 ? tmp18374 : tmp18587;
  assign tmp18585 = s3 ? tmp18586 : 1;
  assign tmp18590 = s1 ? tmp18377 : tmp18434;
  assign tmp18589 = s2 ? 1 : tmp18590;
  assign tmp18588 = s3 ? tmp18589 : 1;
  assign tmp18584 = s4 ? tmp18585 : tmp18588;
  assign tmp18569 = s5 ? tmp18570 : tmp18584;
  assign tmp18560 = s6 ? tmp18561 : tmp18569;
  assign tmp18594 = s2 ? tmp18394 : tmp18568;
  assign tmp18593 = s3 ? tmp18563 : tmp18594;
  assign tmp18592 = s4 ? tmp18562 : tmp18593;
  assign tmp18599 = s1 ? tmp18361 : tmp18443;
  assign tmp18598 = s2 ? tmp18564 : tmp18599;
  assign tmp18601 = s1 ? 1 : tmp18434;
  assign tmp18600 = s2 ? tmp18361 : tmp18601;
  assign tmp18597 = s3 ? tmp18598 : tmp18600;
  assign tmp18603 = s2 ? tmp18580 : tmp18361;
  assign tmp18602 = s3 ? tmp18603 : tmp18582;
  assign tmp18596 = s4 ? tmp18597 : tmp18602;
  assign tmp18607 = s1 ? tmp18361 : tmp18433;
  assign tmp18606 = s2 ? 1 : tmp18607;
  assign tmp18605 = s3 ? tmp18606 : 1;
  assign tmp18604 = s4 ? tmp18396 : tmp18605;
  assign tmp18595 = s5 ? tmp18596 : tmp18604;
  assign tmp18591 = s6 ? tmp18592 : tmp18595;
  assign tmp18559 = s7 ? tmp18560 : tmp18591;
  assign tmp18558 = s8 ? tmp18493 : tmp18559;
  assign tmp18426 = s9 ? tmp18427 : tmp18558;
  assign tmp18616 = s1 ? tmp18433 : 1;
  assign tmp18615 = s2 ? tmp18467 : tmp18616;
  assign tmp18614 = s3 ? tmp18615 : 1;
  assign tmp18618 = s2 ? 1 : tmp18616;
  assign tmp18617 = s3 ? tmp18618 : 1;
  assign tmp18613 = s4 ? tmp18614 : tmp18617;
  assign tmp18612 = s5 ? tmp18481 : tmp18613;
  assign tmp18611 = s6 ? tmp18475 : tmp18612;
  assign tmp18610 = s7 ? tmp18429 : tmp18611;
  assign tmp18609 = s8 ? tmp18610 : tmp18429;
  assign tmp18625 = s2 ? 1 : tmp18433;
  assign tmp18624 = s3 ? tmp18625 : 1;
  assign tmp18623 = s4 ? tmp18469 : tmp18624;
  assign tmp18622 = s5 ? tmp18481 : tmp18623;
  assign tmp18621 = s6 ? tmp18475 : tmp18622;
  assign tmp18628 = s4 ? tmp18396 : tmp18398;
  assign tmp18627 = s5 ? tmp18596 : tmp18628;
  assign tmp18626 = s6 ? tmp18592 : tmp18627;
  assign tmp18620 = s7 ? tmp18621 : tmp18626;
  assign tmp18634 = s2 ? 1 : tmp18497;
  assign tmp18633 = s3 ? tmp18634 : 1;
  assign tmp18632 = s4 ? tmp18554 : tmp18633;
  assign tmp18631 = s5 ? tmp18545 : tmp18632;
  assign tmp18630 = s6 ? tmp18539 : tmp18631;
  assign tmp18637 = s4 ? tmp18614 : tmp18624;
  assign tmp18636 = s5 ? tmp18481 : tmp18637;
  assign tmp18635 = s6 ? tmp18475 : tmp18636;
  assign tmp18629 = s7 ? tmp18630 : tmp18635;
  assign tmp18619 = s8 ? tmp18620 : tmp18629;
  assign tmp18608 = s9 ? tmp18609 : tmp18619;
  assign tmp18425 = s10 ? tmp18426 : tmp18608;
  assign tmp18641 = s7 ? tmp18474 : tmp18591;
  assign tmp18642 = s7 ? tmp18538 : tmp18611;
  assign tmp18640 = s8 ? tmp18641 : tmp18642;
  assign tmp18639 = s9 ? tmp18609 : tmp18640;
  assign tmp18638 = s10 ? tmp18426 : tmp18639;
  assign tmp18424 = s11 ? tmp18425 : tmp18638;
  assign tmp18423 = ~(s12 ? tmp18424 : 1);
  assign tmp18421 = s13 ? tmp18422 : tmp18423;
  assign tmp18196 = s14 ? tmp18197 : tmp18421;
  assign tmp18653 = ~(l2 ? 1 : tmp18498);
  assign tmp18652 = l1 ? 1 : tmp18653;
  assign tmp18651 = s1 ? tmp18652 : tmp18574;
  assign tmp18657 = ~(l1 ? 1 : tmp18653);
  assign tmp18656 = s0 ? 1 : tmp18657;
  assign tmp18658 = ~(s0 ? tmp18361 : tmp18652);
  assign tmp18655 = s1 ? tmp18656 : tmp18658;
  assign tmp18659 = ~(s1 ? tmp18443 : tmp18652);
  assign tmp18654 = ~(s2 ? tmp18655 : tmp18659);
  assign tmp18650 = s3 ? tmp18651 : tmp18654;
  assign tmp18662 = s1 ? 1 : tmp18657;
  assign tmp18664 = s0 ? tmp18652 : 0;
  assign tmp18663 = ~(s1 ? tmp18664 : 0);
  assign tmp18661 = s2 ? tmp18662 : tmp18663;
  assign tmp18666 = s1 ? 1 : tmp18656;
  assign tmp18665 = s2 ? tmp18666 : tmp18657;
  assign tmp18660 = ~(s3 ? tmp18661 : tmp18665);
  assign tmp18649 = s4 ? tmp18650 : tmp18660;
  assign tmp18671 = s1 ? tmp18443 : 0;
  assign tmp18673 = ~(s0 ? tmp18652 : 0);
  assign tmp18672 = ~(s1 ? tmp18363 : tmp18673);
  assign tmp18670 = s2 ? tmp18671 : tmp18672;
  assign tmp18675 = s1 ? tmp18363 : tmp18656;
  assign tmp18674 = ~(s2 ? tmp18675 : tmp18657);
  assign tmp18669 = s3 ? tmp18670 : tmp18674;
  assign tmp18678 = s1 ? tmp18652 : 0;
  assign tmp18677 = s2 ? tmp18678 : 0;
  assign tmp18679 = ~(s2 ? tmp18656 : tmp18657);
  assign tmp18676 = s3 ? tmp18677 : tmp18679;
  assign tmp18668 = s4 ? tmp18669 : tmp18676;
  assign tmp18684 = s0 ? tmp18652 : tmp18361;
  assign tmp18683 = s1 ? tmp18684 : tmp18377;
  assign tmp18682 = s2 ? tmp18683 : tmp18671;
  assign tmp18687 = s0 ? 1 : tmp18498;
  assign tmp18688 = ~(s0 ? tmp18208 : 1);
  assign tmp18686 = s1 ? tmp18687 : tmp18688;
  assign tmp18689 = ~(s1 ? tmp18652 : tmp18664);
  assign tmp18685 = ~(s2 ? tmp18686 : tmp18689);
  assign tmp18681 = s3 ? tmp18682 : tmp18685;
  assign tmp18692 = s1 ? tmp18363 : tmp18658;
  assign tmp18693 = ~(s1 ? tmp18377 : 0);
  assign tmp18691 = s2 ? tmp18692 : tmp18693;
  assign tmp18697 = l1 ? 1 : tmp18208;
  assign tmp18696 = s0 ? tmp18361 : tmp18697;
  assign tmp18695 = s1 ? tmp18696 : tmp18652;
  assign tmp18699 = s0 ? tmp18208 : tmp18361;
  assign tmp18698 = s1 ? tmp18664 : tmp18699;
  assign tmp18694 = ~(s2 ? tmp18695 : tmp18698);
  assign tmp18690 = ~(s3 ? tmp18691 : tmp18694);
  assign tmp18680 = s4 ? tmp18681 : tmp18690;
  assign tmp18667 = s5 ? tmp18668 : tmp18680;
  assign tmp18648 = s6 ? tmp18649 : tmp18667;
  assign tmp18703 = s2 ? tmp18662 : tmp18657;
  assign tmp18702 = ~(s3 ? tmp18661 : tmp18703);
  assign tmp18701 = s4 ? tmp18650 : tmp18702;
  assign tmp18708 = s1 ? tmp18361 : tmp18664;
  assign tmp18707 = s2 ? tmp18671 : tmp18708;
  assign tmp18710 = s1 ? tmp18361 : tmp18652;
  assign tmp18709 = s2 ? tmp18710 : tmp18652;
  assign tmp18706 = s3 ? tmp18707 : tmp18709;
  assign tmp18705 = s4 ? tmp18706 : tmp18676;
  assign tmp18714 = s1 ? tmp18684 : tmp18361;
  assign tmp18713 = s2 ? tmp18714 : 0;
  assign tmp18716 = s1 ? tmp18208 : 1;
  assign tmp18717 = s1 ? tmp18652 : tmp18664;
  assign tmp18715 = s2 ? tmp18716 : tmp18717;
  assign tmp18712 = s3 ? tmp18713 : tmp18715;
  assign tmp18719 = s2 ? tmp18710 : tmp18361;
  assign tmp18718 = s3 ? tmp18719 : tmp18652;
  assign tmp18711 = s4 ? tmp18712 : tmp18718;
  assign tmp18704 = s5 ? tmp18705 : tmp18711;
  assign tmp18700 = s6 ? tmp18701 : tmp18704;
  assign tmp18647 = s7 ? tmp18648 : tmp18700;
  assign tmp18721 = s8 ? tmp18647 : tmp18648;
  assign tmp18720 = s9 ? tmp18721 : tmp18700;
  assign tmp18646 = s10 ? tmp18647 : tmp18720;
  assign tmp18730 = s0 ? 1 : tmp18208;
  assign tmp18729 = s1 ? 1 : tmp18730;
  assign tmp18732 = s0 ? 1 : tmp18211;
  assign tmp18733 = s1 ? 1 : tmp18211;
  assign tmp18731 = s2 ? tmp18732 : tmp18733;
  assign tmp18728 = s3 ? tmp18729 : tmp18731;
  assign tmp18735 = s2 ? tmp18733 : 1;
  assign tmp18736 = s2 ? tmp18733 : tmp18211;
  assign tmp18734 = s3 ? tmp18735 : tmp18736;
  assign tmp18727 = s4 ? tmp18728 : tmp18734;
  assign tmp18741 = s1 ? tmp18208 : tmp18220;
  assign tmp18740 = s2 ? tmp18716 : tmp18741;
  assign tmp18743 = s1 ? 1 : tmp18732;
  assign tmp18742 = s2 ? tmp18743 : tmp18211;
  assign tmp18739 = s3 ? tmp18740 : tmp18742;
  assign tmp18746 = s1 ? tmp18211 : 1;
  assign tmp18745 = s2 ? tmp18746 : 1;
  assign tmp18748 = s1 ? 1 : tmp18220;
  assign tmp18747 = s2 ? tmp18743 : tmp18748;
  assign tmp18744 = s3 ? tmp18745 : tmp18747;
  assign tmp18738 = s4 ? tmp18739 : tmp18744;
  assign tmp18751 = s2 ? tmp18211 : 1;
  assign tmp18754 = s0 ? tmp18361 : tmp18354;
  assign tmp18753 = s1 ? tmp18361 : tmp18754;
  assign tmp18755 = ~(s1 ? tmp18211 : 1);
  assign tmp18752 = ~(s2 ? tmp18753 : tmp18755);
  assign tmp18750 = s3 ? tmp18751 : tmp18752;
  assign tmp18758 = s1 ? tmp18730 : tmp18211;
  assign tmp18759 = s1 ? tmp18730 : 1;
  assign tmp18757 = s2 ? tmp18758 : tmp18759;
  assign tmp18761 = s1 ? tmp18732 : tmp18211;
  assign tmp18763 = ~(s0 ? tmp18361 : tmp18498);
  assign tmp18762 = s1 ? 1 : tmp18763;
  assign tmp18760 = s2 ? tmp18761 : tmp18762;
  assign tmp18756 = s3 ? tmp18757 : tmp18760;
  assign tmp18749 = s4 ? tmp18750 : tmp18756;
  assign tmp18737 = s5 ? tmp18738 : tmp18749;
  assign tmp18726 = s6 ? tmp18727 : tmp18737;
  assign tmp18767 = s3 ? tmp18740 : tmp18736;
  assign tmp18768 = s3 ? tmp18745 : tmp18733;
  assign tmp18766 = s4 ? tmp18767 : tmp18768;
  assign tmp18772 = s1 ? tmp18361 : tmp18354;
  assign tmp18771 = ~(s2 ? tmp18772 : tmp18755);
  assign tmp18770 = s3 ? tmp18745 : tmp18771;
  assign tmp18774 = s2 ? tmp18211 : tmp18208;
  assign tmp18773 = s3 ? tmp18774 : tmp18211;
  assign tmp18769 = s4 ? tmp18770 : tmp18773;
  assign tmp18765 = s5 ? tmp18766 : tmp18769;
  assign tmp18764 = s6 ? tmp18727 : tmp18765;
  assign tmp18725 = s7 ? tmp18726 : tmp18764;
  assign tmp18778 = s3 ? tmp18735 : tmp18742;
  assign tmp18777 = s4 ? tmp18728 : tmp18778;
  assign tmp18776 = s6 ? tmp18777 : tmp18737;
  assign tmp18775 = s7 ? tmp18776 : tmp18764;
  assign tmp18724 = s8 ? tmp18725 : tmp18775;
  assign tmp18723 = s9 ? tmp18724 : tmp18775;
  assign tmp18780 = s8 ? tmp18775 : tmp18776;
  assign tmp18779 = s9 ? tmp18780 : tmp18764;
  assign tmp18722 = s10 ? tmp18723 : tmp18779;
  assign tmp18645 = s12 ? tmp18646 : tmp18722;
  assign tmp18644 = s13 ? 1 : tmp18645;
  assign tmp18792 = l1 ? tmp18209 : 1;
  assign tmp18791 = s0 ? 1 : tmp18792;
  assign tmp18794 = s1 ? tmp18791 : tmp18792;
  assign tmp18796 = s0 ? tmp18792 : 1;
  assign tmp18795 = s1 ? tmp18796 : tmp18792;
  assign tmp18793 = s2 ? tmp18794 : tmp18795;
  assign tmp18790 = s3 ? tmp18791 : tmp18793;
  assign tmp18799 = s1 ? 1 : tmp18792;
  assign tmp18800 = s1 ? tmp18796 : 1;
  assign tmp18798 = s2 ? tmp18799 : tmp18800;
  assign tmp18802 = s1 ? 1 : tmp18363;
  assign tmp18801 = s2 ? tmp18802 : tmp18792;
  assign tmp18797 = s3 ? tmp18798 : tmp18801;
  assign tmp18789 = s4 ? tmp18790 : tmp18797;
  assign tmp18807 = s1 ? tmp18791 : tmp18796;
  assign tmp18806 = s2 ? tmp18800 : tmp18807;
  assign tmp18810 = s0 ? tmp18792 : 0;
  assign tmp18809 = s1 ? tmp18810 : tmp18792;
  assign tmp18808 = s2 ? tmp18791 : tmp18809;
  assign tmp18805 = s3 ? tmp18806 : tmp18808;
  assign tmp18815 = ~(l1 ? tmp18209 : 1);
  assign tmp18814 = s0 ? tmp18361 : tmp18815;
  assign tmp18813 = s1 ? tmp18814 : 0;
  assign tmp18812 = s2 ? tmp18813 : 0;
  assign tmp18817 = s1 ? tmp18792 : tmp18791;
  assign tmp18818 = ~(s1 ? 1 : tmp18375);
  assign tmp18816 = ~(s2 ? tmp18817 : tmp18818);
  assign tmp18811 = ~(s3 ? tmp18812 : tmp18816);
  assign tmp18804 = s4 ? tmp18805 : tmp18811;
  assign tmp18823 = ~(s0 ? 1 : tmp18815);
  assign tmp18822 = s1 ? tmp18810 : tmp18823;
  assign tmp18821 = s2 ? tmp18822 : tmp18800;
  assign tmp18825 = s1 ? tmp18223 : 0;
  assign tmp18826 = ~(s1 ? tmp18361 : tmp18443);
  assign tmp18824 = s2 ? tmp18825 : tmp18826;
  assign tmp18820 = s3 ? tmp18821 : tmp18824;
  assign tmp18829 = s1 ? tmp18237 : tmp18792;
  assign tmp18831 = s0 ? 1 : tmp18815;
  assign tmp18830 = ~(s1 ? tmp18831 : 0);
  assign tmp18828 = s2 ? tmp18829 : tmp18830;
  assign tmp18833 = s1 ? tmp18792 : tmp18823;
  assign tmp18834 = ~(s1 ? tmp18443 : tmp18255);
  assign tmp18832 = s2 ? tmp18833 : tmp18834;
  assign tmp18827 = s3 ? tmp18828 : tmp18832;
  assign tmp18819 = s4 ? tmp18820 : tmp18827;
  assign tmp18803 = s5 ? tmp18804 : tmp18819;
  assign tmp18788 = s6 ? tmp18789 : tmp18803;
  assign tmp18839 = s1 ? 1 : tmp18352;
  assign tmp18838 = s2 ? tmp18839 : tmp18792;
  assign tmp18837 = s3 ? tmp18798 : tmp18838;
  assign tmp18836 = s4 ? tmp18790 : tmp18837;
  assign tmp18844 = s1 ? tmp18792 : tmp18796;
  assign tmp18843 = s2 ? tmp18800 : tmp18844;
  assign tmp18845 = s2 ? tmp18792 : tmp18809;
  assign tmp18842 = s3 ? tmp18843 : tmp18845;
  assign tmp18848 = ~(s1 ? 1 : tmp18361);
  assign tmp18847 = ~(s2 ? tmp18792 : tmp18848);
  assign tmp18846 = ~(s3 ? tmp18812 : tmp18847);
  assign tmp18841 = s4 ? tmp18842 : tmp18846;
  assign tmp18851 = s2 ? tmp18809 : tmp18800;
  assign tmp18853 = s1 ? tmp18361 : 0;
  assign tmp18852 = ~(s2 ? 1 : tmp18853);
  assign tmp18850 = s3 ? tmp18851 : tmp18852;
  assign tmp18849 = s4 ? tmp18850 : tmp18792;
  assign tmp18840 = s5 ? tmp18841 : tmp18849;
  assign tmp18835 = s6 ? tmp18836 : tmp18840;
  assign tmp18787 = s7 ? tmp18788 : tmp18835;
  assign tmp18861 = s0 ? tmp18209 : tmp18792;
  assign tmp18860 = s1 ? tmp18237 : tmp18861;
  assign tmp18859 = s2 ? tmp18860 : tmp18830;
  assign tmp18864 = s0 ? tmp18792 : tmp18209;
  assign tmp18863 = s1 ? tmp18864 : tmp18823;
  assign tmp18862 = s2 ? tmp18863 : tmp18834;
  assign tmp18858 = s3 ? tmp18859 : tmp18862;
  assign tmp18857 = s4 ? tmp18820 : tmp18858;
  assign tmp18856 = s5 ? tmp18804 : tmp18857;
  assign tmp18855 = s6 ? tmp18789 : tmp18856;
  assign tmp18869 = s2 ? tmp18809 : 1;
  assign tmp18868 = s3 ? tmp18869 : tmp18852;
  assign tmp18872 = s1 ? tmp18209 : tmp18792;
  assign tmp18871 = s2 ? tmp18872 : tmp18792;
  assign tmp18870 = s3 ? tmp18871 : tmp18872;
  assign tmp18867 = s4 ? tmp18868 : tmp18870;
  assign tmp18866 = s5 ? tmp18841 : tmp18867;
  assign tmp18865 = s6 ? tmp18836 : tmp18866;
  assign tmp18854 = s7 ? tmp18855 : tmp18865;
  assign tmp18786 = s8 ? tmp18787 : tmp18854;
  assign tmp18877 = s4 ? tmp18868 : tmp18792;
  assign tmp18876 = s5 ? tmp18841 : tmp18877;
  assign tmp18875 = s6 ? tmp18836 : tmp18876;
  assign tmp18874 = s7 ? tmp18788 : tmp18875;
  assign tmp18873 = s8 ? tmp18854 : tmp18874;
  assign tmp18785 = s9 ? tmp18786 : tmp18873;
  assign tmp18884 = s3 ? tmp18792 : tmp18872;
  assign tmp18883 = s4 ? tmp18868 : tmp18884;
  assign tmp18882 = s5 ? tmp18841 : tmp18883;
  assign tmp18881 = s6 ? tmp18836 : tmp18882;
  assign tmp18880 = s7 ? tmp18788 : tmp18881;
  assign tmp18879 = s8 ? tmp18880 : tmp18788;
  assign tmp18889 = s4 ? tmp18850 : tmp18884;
  assign tmp18888 = s5 ? tmp18841 : tmp18889;
  assign tmp18887 = s6 ? tmp18836 : tmp18888;
  assign tmp18886 = s7 ? tmp18887 : tmp18875;
  assign tmp18890 = s7 ? tmp18865 : tmp18881;
  assign tmp18885 = s8 ? tmp18886 : tmp18890;
  assign tmp18878 = s9 ? tmp18879 : tmp18885;
  assign tmp18784 = s10 ? tmp18785 : tmp18878;
  assign tmp18894 = s7 ? tmp18835 : tmp18875;
  assign tmp18893 = s8 ? tmp18894 : tmp18890;
  assign tmp18892 = s9 ? tmp18879 : tmp18893;
  assign tmp18891 = s10 ? tmp18785 : tmp18892;
  assign tmp18783 = s11 ? tmp18784 : tmp18891;
  assign tmp18782 = s12 ? 1 : tmp18783;
  assign tmp18901 = s1 ? tmp18208 : 0;
  assign tmp18902 = ~(s2 ? tmp18510 : tmp18550);
  assign tmp18900 = s3 ? tmp18901 : tmp18902;
  assign tmp18906 = s0 ? tmp18208 : 0;
  assign tmp18905 = ~(s1 ? tmp18906 : 0);
  assign tmp18904 = s2 ? tmp18550 : tmp18905;
  assign tmp18908 = s1 ? 1 : tmp18510;
  assign tmp18907 = s2 ? tmp18908 : tmp18497;
  assign tmp18903 = ~(s3 ? tmp18904 : tmp18907);
  assign tmp18899 = s4 ? tmp18900 : tmp18903;
  assign tmp18913 = s1 ? 1 : tmp18534;
  assign tmp18912 = s2 ? 1 : tmp18913;
  assign tmp18911 = s3 ? tmp18912 : tmp18907;
  assign tmp18915 = s2 ? tmp18510 : tmp18497;
  assign tmp18914 = s3 ? tmp18528 : tmp18915;
  assign tmp18910 = s4 ? tmp18911 : tmp18914;
  assign tmp18919 = s1 ? tmp18506 : tmp18446;
  assign tmp18918 = s2 ? tmp18919 : 1;
  assign tmp18921 = s1 ? tmp18510 : tmp18497;
  assign tmp18923 = ~(s0 ? tmp18208 : 0);
  assign tmp18922 = s1 ? tmp18497 : tmp18923;
  assign tmp18920 = s2 ? tmp18921 : tmp18922;
  assign tmp18917 = s3 ? tmp18918 : tmp18920;
  assign tmp18926 = ~(s1 ? tmp18223 : 0);
  assign tmp18925 = s2 ? tmp18908 : tmp18926;
  assign tmp18927 = s2 ? tmp18921 : tmp18534;
  assign tmp18924 = s3 ? tmp18925 : tmp18927;
  assign tmp18916 = s4 ? tmp18917 : tmp18924;
  assign tmp18909 = ~(s5 ? tmp18910 : tmp18916);
  assign tmp18898 = s6 ? tmp18899 : tmp18909;
  assign tmp18931 = s2 ? tmp18550 : tmp18497;
  assign tmp18930 = ~(s3 ? tmp18904 : tmp18931);
  assign tmp18929 = s4 ? tmp18900 : tmp18930;
  assign tmp18934 = s3 ? tmp18912 : tmp18931;
  assign tmp18933 = s4 ? tmp18934 : tmp18914;
  assign tmp18938 = s1 ? tmp18506 : 1;
  assign tmp18937 = s2 ? tmp18938 : 1;
  assign tmp18940 = ~(s1 ? tmp18208 : 0);
  assign tmp18939 = s2 ? tmp18497 : tmp18940;
  assign tmp18936 = s3 ? tmp18937 : tmp18939;
  assign tmp18942 = s2 ? tmp18550 : 1;
  assign tmp18941 = s3 ? tmp18942 : tmp18497;
  assign tmp18935 = s4 ? tmp18936 : tmp18941;
  assign tmp18932 = ~(s5 ? tmp18933 : tmp18935);
  assign tmp18928 = s6 ? tmp18929 : tmp18932;
  assign tmp18897 = s7 ? tmp18898 : tmp18928;
  assign tmp18944 = s8 ? tmp18897 : tmp18898;
  assign tmp18943 = s9 ? tmp18944 : tmp18928;
  assign tmp18896 = s10 ? tmp18897 : tmp18943;
  assign tmp18954 = l2 ? 1 : tmp18498;
  assign tmp18953 = l1 ? tmp18954 : 1;
  assign tmp18952 = s0 ? 1 : tmp18953;
  assign tmp18956 = s1 ? tmp18952 : tmp18953;
  assign tmp18957 = s1 ? tmp18792 : tmp18953;
  assign tmp18955 = s2 ? tmp18956 : tmp18957;
  assign tmp18951 = s3 ? tmp18952 : tmp18955;
  assign tmp18960 = s1 ? 1 : tmp18953;
  assign tmp18959 = s2 ? tmp18960 : tmp18800;
  assign tmp18964 = ~(l1 ? tmp18208 : 0);
  assign tmp18963 = s0 ? 1 : tmp18964;
  assign tmp18962 = s1 ? 1 : tmp18963;
  assign tmp18961 = s2 ? tmp18962 : tmp18953;
  assign tmp18958 = s3 ? tmp18959 : tmp18961;
  assign tmp18950 = s4 ? tmp18951 : tmp18958;
  assign tmp18970 = s0 ? tmp18953 : 1;
  assign tmp18969 = s1 ? tmp18970 : 1;
  assign tmp18975 = ~(l4 ? 1 : 0);
  assign tmp18974 = ~(l2 ? 1 : tmp18975);
  assign tmp18973 = l1 ? tmp18209 : tmp18974;
  assign tmp18972 = s0 ? tmp18953 : tmp18973;
  assign tmp18971 = s1 ? tmp18952 : tmp18972;
  assign tmp18968 = s2 ? tmp18969 : tmp18971;
  assign tmp18977 = s0 ? tmp18973 : tmp18953;
  assign tmp18976 = s2 ? tmp18977 : tmp18953;
  assign tmp18967 = s3 ? tmp18968 : tmp18976;
  assign tmp18980 = s1 ? tmp18953 : 1;
  assign tmp18979 = s2 ? tmp18980 : 1;
  assign tmp18984 = l1 ? tmp18208 : 0;
  assign tmp18983 = s0 ? tmp18984 : 1;
  assign tmp18982 = ~(s1 ? 1 : tmp18983);
  assign tmp18981 = s2 ? tmp18952 : tmp18982;
  assign tmp18978 = s3 ? tmp18979 : tmp18981;
  assign tmp18966 = s4 ? tmp18967 : tmp18978;
  assign tmp18987 = s2 ? tmp18953 : tmp18800;
  assign tmp18989 = s1 ? 1 : tmp18687;
  assign tmp18990 = ~(s1 ? tmp18984 : tmp18443);
  assign tmp18988 = s2 ? tmp18989 : tmp18990;
  assign tmp18986 = s3 ? tmp18987 : tmp18988;
  assign tmp18992 = s2 ? tmp18956 : tmp18980;
  assign tmp18995 = ~(s0 ? 1 : tmp18953);
  assign tmp18994 = ~(s1 ? tmp18443 : tmp18995);
  assign tmp18993 = s2 ? tmp18953 : tmp18994;
  assign tmp18991 = s3 ? tmp18992 : tmp18993;
  assign tmp18985 = s4 ? tmp18986 : tmp18991;
  assign tmp18965 = s5 ? tmp18966 : tmp18985;
  assign tmp18949 = s6 ? tmp18950 : tmp18965;
  assign tmp19000 = s1 ? 1 : tmp18964;
  assign tmp18999 = s2 ? tmp19000 : tmp18953;
  assign tmp18998 = s3 ? tmp18959 : tmp18999;
  assign tmp18997 = s4 ? tmp18951 : tmp18998;
  assign tmp19005 = s1 ? tmp18953 : tmp18972;
  assign tmp19004 = s2 ? tmp18969 : tmp19005;
  assign tmp19003 = s3 ? tmp19004 : tmp18953;
  assign tmp19008 = ~(s1 ? 1 : tmp18984);
  assign tmp19007 = s2 ? tmp18952 : tmp19008;
  assign tmp19006 = s3 ? tmp18979 : tmp19007;
  assign tmp19002 = s4 ? tmp19003 : tmp19006;
  assign tmp19012 = s1 ? tmp18953 : tmp18792;
  assign tmp19011 = s2 ? tmp19012 : 1;
  assign tmp19014 = s1 ? 1 : tmp18498;
  assign tmp19015 = ~(s1 ? tmp18361 : 0);
  assign tmp19013 = s2 ? tmp19014 : tmp19015;
  assign tmp19010 = s3 ? tmp19011 : tmp19013;
  assign tmp19009 = s4 ? tmp19010 : tmp18953;
  assign tmp19001 = s5 ? tmp19002 : tmp19009;
  assign tmp18996 = s6 ? tmp18997 : tmp19001;
  assign tmp18948 = s7 ? tmp18949 : tmp18996;
  assign tmp19021 = s1 ? tmp18796 : tmp18953;
  assign tmp19020 = s2 ? tmp18956 : tmp19021;
  assign tmp19019 = s3 ? tmp18952 : tmp19020;
  assign tmp19028 = l3 ? 1 : tmp18975;
  assign tmp19027 = l2 ? tmp19028 : 1;
  assign tmp19026 = l1 ? 1 : tmp19027;
  assign tmp19025 = s0 ? tmp18792 : tmp19026;
  assign tmp19024 = s1 ? tmp19025 : 1;
  assign tmp19023 = s2 ? tmp18960 : tmp19024;
  assign tmp19022 = s3 ? tmp19023 : tmp18961;
  assign tmp19018 = s4 ? tmp19019 : tmp19022;
  assign tmp19033 = s1 ? tmp18952 : tmp18970;
  assign tmp19032 = s2 ? tmp18969 : tmp19033;
  assign tmp19034 = s2 ? tmp18952 : tmp18953;
  assign tmp19031 = s3 ? tmp19032 : tmp19034;
  assign tmp19030 = s4 ? tmp19031 : tmp18978;
  assign tmp19029 = s5 ? tmp19030 : tmp18985;
  assign tmp19017 = s6 ? tmp19018 : tmp19029;
  assign tmp19037 = s3 ? tmp19023 : tmp18999;
  assign tmp19036 = s4 ? tmp19019 : tmp19037;
  assign tmp19042 = s1 ? tmp18953 : tmp18970;
  assign tmp19041 = s2 ? tmp18969 : tmp19042;
  assign tmp19040 = s3 ? tmp19041 : tmp18953;
  assign tmp19039 = s4 ? tmp19040 : tmp19006;
  assign tmp19038 = s5 ? tmp19039 : tmp19009;
  assign tmp19035 = s6 ? tmp19036 : tmp19038;
  assign tmp19016 = s7 ? tmp19017 : tmp19035;
  assign tmp18947 = s8 ? tmp18948 : tmp19016;
  assign tmp19046 = s4 ? tmp19019 : tmp18958;
  assign tmp19045 = s6 ? tmp19046 : tmp19029;
  assign tmp19048 = s4 ? tmp19019 : tmp18998;
  assign tmp19047 = s6 ? tmp19048 : tmp19038;
  assign tmp19044 = s7 ? tmp19045 : tmp19047;
  assign tmp19043 = s8 ? tmp19016 : tmp19044;
  assign tmp18946 = s9 ? tmp18947 : tmp19043;
  assign tmp19059 = l1 ? 1 : tmp18975;
  assign tmp19058 = s0 ? tmp19059 : tmp18953;
  assign tmp19057 = s1 ? tmp18791 : tmp19058;
  assign tmp19056 = s2 ? tmp19057 : tmp18982;
  assign tmp19055 = s3 ? tmp18979 : tmp19056;
  assign tmp19054 = s4 ? tmp19031 : tmp19055;
  assign tmp19053 = s5 ? tmp19054 : tmp18985;
  assign tmp19052 = s6 ? tmp19046 : tmp19053;
  assign tmp19051 = s7 ? tmp19052 : tmp19047;
  assign tmp19050 = s8 ? tmp19051 : tmp19052;
  assign tmp19061 = s7 ? tmp18996 : tmp19047;
  assign tmp19062 = s7 ? tmp19035 : tmp19047;
  assign tmp19060 = s8 ? tmp19061 : tmp19062;
  assign tmp19049 = s9 ? tmp19050 : tmp19060;
  assign tmp18945 = ~(s10 ? tmp18946 : tmp19049);
  assign tmp18895 = ~(s12 ? tmp18896 : tmp18945);
  assign tmp18781 = ~(s13 ? tmp18782 : tmp18895);
  assign tmp18643 = s14 ? tmp18644 : tmp18781;
  assign tmp18195 = s15 ? tmp18196 : tmp18643;
  assign tmp19077 = s0 ? tmp18209 : tmp18352;
  assign tmp19076 = s1 ? tmp18310 : tmp19077;
  assign tmp19075 = s2 ? tmp18309 : tmp19076;
  assign tmp19079 = s0 ? tmp18361 : tmp18256;
  assign tmp19080 = s1 ? 1 : tmp18314;
  assign tmp19078 = ~(s2 ? tmp19079 : tmp19080);
  assign tmp19074 = s3 ? tmp19075 : tmp19078;
  assign tmp19073 = s4 ? tmp19074 : tmp18316;
  assign tmp19072 = s5 ? tmp19073 : tmp18249;
  assign tmp19071 = s6 ? tmp18283 : tmp19072;
  assign tmp19086 = s1 ? tmp18286 : tmp19077;
  assign tmp19085 = s2 ? tmp18291 : tmp19086;
  assign tmp19084 = s3 ? tmp19085 : tmp18338;
  assign tmp19090 = l1 ? tmp18954 : 0;
  assign tmp19092 = ~(l1 ? tmp18954 : 0);
  assign tmp19091 = ~(s0 ? tmp18286 : tmp19092);
  assign tmp19089 = s1 ? tmp19090 : tmp19091;
  assign tmp19088 = s2 ? tmp18318 : tmp19089;
  assign tmp19087 = ~(s3 ? tmp19088 : tmp18341);
  assign tmp19083 = s4 ? tmp19084 : tmp19087;
  assign tmp19082 = s5 ? tmp19083 : tmp18276;
  assign tmp19081 = s6 ? tmp18327 : tmp19082;
  assign tmp19070 = s7 ? tmp19071 : tmp19081;
  assign tmp19069 = s8 ? tmp18202 : tmp19070;
  assign tmp19099 = s0 ? tmp19090 : tmp18792;
  assign tmp19098 = s2 ? tmp19090 : tmp19099;
  assign tmp19101 = s1 ? tmp19090 : tmp18796;
  assign tmp19103 = s0 ? tmp19090 : tmp18361;
  assign tmp19104 = s0 ? 1 : tmp19090;
  assign tmp19102 = s1 ? tmp19103 : tmp19104;
  assign tmp19100 = s2 ? tmp19101 : tmp19102;
  assign tmp19097 = s3 ? tmp19098 : tmp19100;
  assign tmp19096 = s4 ? tmp19090 : tmp19097;
  assign tmp19109 = s1 ? tmp19090 : tmp18361;
  assign tmp19108 = s2 ? tmp19090 : tmp19109;
  assign tmp19112 = s0 ? tmp19090 : 1;
  assign tmp19111 = s1 ? 1 : tmp19112;
  assign tmp19110 = s2 ? tmp18361 : tmp19111;
  assign tmp19107 = s3 ? tmp19108 : tmp19110;
  assign tmp19115 = s1 ? tmp19104 : tmp19112;
  assign tmp19116 = s1 ? tmp19112 : tmp19090;
  assign tmp19114 = s2 ? tmp19115 : tmp19116;
  assign tmp19117 = s2 ? tmp18374 : 1;
  assign tmp19113 = s3 ? tmp19114 : tmp19117;
  assign tmp19106 = s4 ? tmp19107 : tmp19113;
  assign tmp19118 = s4 ? tmp18372 : tmp18378;
  assign tmp19105 = s5 ? tmp19106 : tmp19118;
  assign tmp19095 = s6 ? tmp19096 : tmp19105;
  assign tmp19123 = s1 ? tmp19099 : tmp19090;
  assign tmp19122 = s2 ? tmp19090 : tmp19123;
  assign tmp19125 = s1 ? tmp19090 : 1;
  assign tmp19124 = s2 ? tmp19125 : tmp19102;
  assign tmp19121 = s3 ? tmp19122 : tmp19124;
  assign tmp19120 = s4 ? tmp19090 : tmp19121;
  assign tmp19129 = s2 ? tmp19115 : tmp19090;
  assign tmp19128 = s3 ? tmp19129 : tmp19117;
  assign tmp19127 = s4 ? tmp19107 : tmp19128;
  assign tmp19126 = s5 ? tmp19127 : tmp18628;
  assign tmp19119 = s6 ? tmp19120 : tmp19126;
  assign tmp19094 = ~(s7 ? tmp19095 : tmp19119);
  assign tmp19093 = s8 ? tmp19070 : tmp19094;
  assign tmp19068 = s9 ? tmp19069 : tmp19093;
  assign tmp19137 = l1 ? tmp18954 : tmp18256;
  assign tmp19138 = s0 ? tmp19090 : tmp19137;
  assign tmp19136 = s1 ? tmp19137 : tmp19138;
  assign tmp19141 = s0 ? tmp19137 : tmp18315;
  assign tmp19140 = s1 ? tmp19141 : tmp19137;
  assign tmp19139 = s2 ? tmp19137 : tmp19140;
  assign tmp19135 = s3 ? tmp19136 : tmp19139;
  assign tmp19145 = s0 ? tmp19137 : tmp19090;
  assign tmp19144 = s1 ? tmp19145 : tmp19137;
  assign tmp19147 = s0 ? tmp19137 : tmp18792;
  assign tmp19146 = s1 ? tmp19147 : tmp19099;
  assign tmp19143 = s2 ? tmp19144 : tmp19146;
  assign tmp19150 = s0 ? tmp19137 : tmp18433;
  assign tmp19151 = s0 ? 1 : tmp19137;
  assign tmp19149 = s1 ? tmp19150 : tmp19151;
  assign tmp19148 = s2 ? tmp19101 : tmp19149;
  assign tmp19142 = s3 ? tmp19143 : tmp19148;
  assign tmp19134 = s4 ? tmp19135 : tmp19142;
  assign tmp19157 = s0 ? tmp19137 : 0;
  assign tmp19159 = ~(l1 ? tmp18954 : tmp18256);
  assign tmp19158 = ~(s0 ? 1 : tmp19159);
  assign tmp19156 = s1 ? tmp19157 : tmp19158;
  assign tmp19161 = s0 ? 1 : tmp19159;
  assign tmp19162 = ~(s0 ? tmp18433 : tmp18361);
  assign tmp19160 = ~(s1 ? tmp19161 : tmp19162);
  assign tmp19155 = s2 ? tmp19156 : tmp19160;
  assign tmp19164 = s1 ? tmp18434 : tmp19079;
  assign tmp19166 = s0 ? tmp19137 : 1;
  assign tmp19165 = s1 ? 1 : tmp19166;
  assign tmp19163 = s2 ? tmp19164 : tmp19165;
  assign tmp19154 = s3 ? tmp19155 : tmp19163;
  assign tmp19169 = s1 ? tmp19151 : tmp19112;
  assign tmp19170 = s1 ? tmp19112 : tmp19145;
  assign tmp19168 = s2 ? tmp19169 : tmp19170;
  assign tmp19171 = ~(s2 ? tmp18252 : 0);
  assign tmp19167 = s3 ? tmp19168 : tmp19171;
  assign tmp19153 = s4 ? tmp19154 : tmp19167;
  assign tmp19172 = ~(s4 ? tmp18250 : tmp18257);
  assign tmp19152 = s5 ? tmp19153 : tmp19172;
  assign tmp19133 = s6 ? tmp19134 : tmp19152;
  assign tmp19177 = s1 ? tmp19147 : tmp19090;
  assign tmp19176 = s2 ? tmp19144 : tmp19177;
  assign tmp19178 = s2 ? tmp19125 : tmp19149;
  assign tmp19175 = s3 ? tmp19176 : tmp19178;
  assign tmp19174 = s4 ? tmp19135 : tmp19175;
  assign tmp19183 = s1 ? tmp19157 : tmp19137;
  assign tmp19184 = s1 ? tmp19137 : tmp18441;
  assign tmp19182 = s2 ? tmp19183 : tmp19184;
  assign tmp19186 = s1 ? tmp18433 : tmp18256;
  assign tmp19185 = s2 ? tmp19186 : tmp19165;
  assign tmp19181 = s3 ? tmp19182 : tmp19185;
  assign tmp19189 = s1 ? tmp19090 : tmp19145;
  assign tmp19188 = s2 ? tmp19169 : tmp19189;
  assign tmp19187 = s3 ? tmp19188 : tmp19171;
  assign tmp19180 = s4 ? tmp19181 : tmp19187;
  assign tmp19190 = ~(s4 ? tmp18277 : tmp18279);
  assign tmp19179 = s5 ? tmp19180 : tmp19190;
  assign tmp19173 = s6 ? tmp19174 : tmp19179;
  assign tmp19132 = s7 ? tmp19133 : tmp19173;
  assign tmp19131 = s8 ? tmp19132 : tmp19133;
  assign tmp19193 = ~(s6 ? tmp19120 : tmp19126);
  assign tmp19192 = s7 ? tmp18410 : tmp19193;
  assign tmp19200 = s1 ? tmp19090 : tmp18304;
  assign tmp19199 = s2 ? tmp18318 : tmp19200;
  assign tmp19198 = ~(s3 ? tmp19199 : tmp18341);
  assign tmp19197 = s4 ? tmp19084 : tmp19198;
  assign tmp19196 = s5 ? tmp19197 : tmp18276;
  assign tmp19195 = s6 ? tmp18327 : tmp19196;
  assign tmp19206 = s1 ? tmp19090 : tmp19137;
  assign tmp19205 = s2 ? tmp19169 : tmp19206;
  assign tmp19204 = s3 ? tmp19205 : tmp19171;
  assign tmp19203 = s4 ? tmp19181 : tmp19204;
  assign tmp19202 = s5 ? tmp19203 : tmp19190;
  assign tmp19201 = ~(s6 ? tmp19174 : tmp19202);
  assign tmp19194 = s7 ? tmp19195 : tmp19201;
  assign tmp19191 = ~(s8 ? tmp19192 : tmp19194);
  assign tmp19130 = ~(s9 ? tmp19131 : tmp19191);
  assign tmp19067 = s10 ? tmp19068 : tmp19130;
  assign tmp19210 = s7 ? tmp18260 : tmp19193;
  assign tmp19212 = ~(s6 ? tmp19174 : tmp19179);
  assign tmp19211 = s7 ? tmp19081 : tmp19212;
  assign tmp19209 = ~(s8 ? tmp19210 : tmp19211);
  assign tmp19208 = ~(s9 ? tmp19131 : tmp19209);
  assign tmp19207 = s10 ? tmp19068 : tmp19208;
  assign tmp19066 = s11 ? tmp19067 : tmp19207;
  assign tmp19223 = s1 ? 1 : tmp18223;
  assign tmp19224 = s1 ? 1 : tmp18446;
  assign tmp19222 = s2 ? tmp19223 : tmp19224;
  assign tmp19221 = s3 ? 1 : tmp19222;
  assign tmp19220 = s4 ? 1 : tmp19221;
  assign tmp19229 = ~(s1 ? 1 : tmp18446);
  assign tmp19228 = s2 ? tmp19223 : tmp19229;
  assign tmp19227 = s3 ? 1 : tmp19228;
  assign tmp19232 = s1 ? tmp18223 : tmp18446;
  assign tmp19233 = ~(s1 ? tmp18223 : 1);
  assign tmp19231 = s2 ? tmp19232 : tmp19233;
  assign tmp19230 = ~(s3 ? tmp19231 : 1);
  assign tmp19226 = s4 ? tmp19227 : tmp19230;
  assign tmp19225 = s5 ? tmp19226 : 0;
  assign tmp19219 = s6 ? tmp19220 : tmp19225;
  assign tmp19239 = s1 ? 1 : 0;
  assign tmp19238 = s2 ? tmp19239 : tmp19229;
  assign tmp19237 = s3 ? 1 : tmp19238;
  assign tmp19241 = s2 ? tmp19232 : 0;
  assign tmp19240 = ~(s3 ? tmp19241 : 1);
  assign tmp19236 = s4 ? tmp19237 : tmp19240;
  assign tmp19235 = s5 ? tmp19236 : 0;
  assign tmp19234 = s6 ? tmp19220 : tmp19235;
  assign tmp19218 = s7 ? tmp19219 : tmp19234;
  assign tmp19248 = ~(s1 ? 1 : 0);
  assign tmp19247 = s2 ? tmp19223 : tmp19248;
  assign tmp19246 = s3 ? 1 : tmp19247;
  assign tmp19250 = s2 ? tmp18825 : 0;
  assign tmp19249 = ~(s3 ? tmp19250 : 1);
  assign tmp19245 = s4 ? tmp19246 : tmp19249;
  assign tmp19244 = s5 ? tmp19245 : 0;
  assign tmp19243 = s6 ? tmp19220 : tmp19244;
  assign tmp19257 = ~(l1 ? tmp18209 : 0);
  assign tmp19256 = s0 ? 1 : tmp19257;
  assign tmp19255 = s1 ? 1 : tmp19256;
  assign tmp19254 = s2 ? 1 : tmp19255;
  assign tmp19260 = ~(s0 ? tmp18315 : 1);
  assign tmp19259 = s1 ? 1 : tmp19260;
  assign tmp19258 = s2 ? tmp19259 : tmp19224;
  assign tmp19253 = s3 ? tmp19254 : tmp19258;
  assign tmp19252 = s4 ? 1 : tmp19253;
  assign tmp19264 = s2 ? tmp19239 : tmp19248;
  assign tmp19263 = s3 ? 1 : tmp19264;
  assign tmp19262 = s4 ? tmp19263 : tmp19249;
  assign tmp19261 = s5 ? tmp19262 : 0;
  assign tmp19251 = s6 ? tmp19252 : tmp19261;
  assign tmp19242 = s7 ? tmp19243 : tmp19251;
  assign tmp19217 = s8 ? tmp19218 : tmp19242;
  assign tmp19272 = s0 ? tmp18315 : 1;
  assign tmp19271 = s1 ? tmp18315 : tmp19272;
  assign tmp19274 = s0 ? 1 : tmp18315;
  assign tmp19273 = s1 ? tmp18315 : tmp19274;
  assign tmp19270 = s2 ? tmp19271 : tmp19273;
  assign tmp19269 = s3 ? tmp18315 : tmp19270;
  assign tmp19268 = s4 ? tmp18315 : tmp19269;
  assign tmp19280 = s0 ? tmp18315 : 0;
  assign tmp19281 = ~(s0 ? 1 : tmp19257);
  assign tmp19279 = s1 ? tmp19280 : tmp19281;
  assign tmp19282 = ~(s1 ? tmp18255 : tmp18352);
  assign tmp19278 = s2 ? tmp19279 : tmp19282;
  assign tmp19284 = s1 ? tmp18361 : tmp18375;
  assign tmp19285 = s1 ? 1 : tmp18209;
  assign tmp19283 = s2 ? tmp19284 : tmp19285;
  assign tmp19277 = s3 ? tmp19278 : tmp19283;
  assign tmp19288 = s1 ? tmp18237 : tmp18209;
  assign tmp19287 = s2 ? tmp19288 : tmp18209;
  assign tmp19286 = s3 ? tmp19287 : 1;
  assign tmp19276 = s4 ? tmp19277 : tmp19286;
  assign tmp19275 = s5 ? tmp19276 : 1;
  assign tmp19267 = s6 ? tmp19268 : tmp19275;
  assign tmp19294 = s1 ? tmp19280 : tmp18315;
  assign tmp19295 = s1 ? tmp18209 : tmp18361;
  assign tmp19293 = s2 ? tmp19294 : tmp19295;
  assign tmp19296 = s2 ? tmp18394 : tmp19285;
  assign tmp19292 = s3 ? tmp19293 : tmp19296;
  assign tmp19291 = s4 ? tmp19292 : tmp19286;
  assign tmp19290 = s5 ? tmp19291 : 1;
  assign tmp19289 = s6 ? tmp19268 : tmp19290;
  assign tmp19266 = ~(s7 ? tmp19267 : tmp19289);
  assign tmp19265 = s8 ? tmp19242 : tmp19266;
  assign tmp19216 = s9 ? tmp19217 : tmp19265;
  assign tmp19299 = s7 ? tmp19267 : tmp19289;
  assign tmp19298 = s8 ? tmp19299 : tmp19267;
  assign tmp19305 = s2 ? tmp19239 : tmp19224;
  assign tmp19304 = s3 ? 1 : tmp19305;
  assign tmp19303 = s4 ? 1 : tmp19304;
  assign tmp19302 = s6 ? tmp19303 : tmp19235;
  assign tmp19310 = s1 ? tmp18315 : 1;
  assign tmp19309 = s2 ? tmp19310 : tmp19273;
  assign tmp19308 = s3 ? tmp18315 : tmp19309;
  assign tmp19307 = s4 ? tmp18315 : tmp19308;
  assign tmp19306 = ~(s6 ? tmp19307 : tmp19290);
  assign tmp19301 = s7 ? tmp19302 : tmp19306;
  assign tmp19314 = s3 ? tmp19254 : tmp19305;
  assign tmp19313 = s4 ? 1 : tmp19314;
  assign tmp19312 = s6 ? tmp19313 : tmp19261;
  assign tmp19311 = s7 ? tmp19312 : tmp19306;
  assign tmp19300 = ~(s8 ? tmp19301 : tmp19311);
  assign tmp19297 = ~(s9 ? tmp19298 : tmp19300);
  assign tmp19215 = s10 ? tmp19216 : tmp19297;
  assign tmp19319 = ~(s6 ? tmp19268 : tmp19290);
  assign tmp19318 = s7 ? tmp19234 : tmp19319;
  assign tmp19320 = s7 ? tmp19251 : tmp19319;
  assign tmp19317 = ~(s8 ? tmp19318 : tmp19320);
  assign tmp19316 = ~(s9 ? tmp19298 : tmp19317);
  assign tmp19315 = s10 ? tmp19216 : tmp19316;
  assign tmp19214 = s11 ? tmp19215 : tmp19315;
  assign tmp19213 = s12 ? 1 : tmp19214;
  assign tmp19065 = s13 ? tmp19066 : tmp19213;
  assign tmp19330 = s2 ? tmp19284 : tmp18568;
  assign tmp19329 = s3 ? tmp18361 : tmp19330;
  assign tmp19328 = s4 ? tmp18361 : tmp19329;
  assign tmp19334 = ~(s1 ? tmp18223 : tmp18352);
  assign tmp19333 = s2 ? tmp18573 : tmp19334;
  assign tmp19332 = s3 ? tmp19333 : tmp18370;
  assign tmp19331 = s4 ? tmp19332 : 1;
  assign tmp19327 = s6 ? tmp19328 : tmp19331;
  assign tmp19338 = s2 ? tmp18361 : tmp18394;
  assign tmp19337 = s3 ? tmp19338 : tmp18594;
  assign tmp19336 = s4 ? tmp18361 : tmp19337;
  assign tmp19342 = s1 ? 1 : tmp18361;
  assign tmp19341 = s2 ? tmp18564 : tmp19342;
  assign tmp19344 = l1 ? 1 : tmp18209;
  assign tmp19343 = s2 ? tmp19344 : 1;
  assign tmp19340 = s3 ? tmp19341 : tmp19343;
  assign tmp19339 = s4 ? tmp19340 : 1;
  assign tmp19335 = s6 ? tmp19336 : tmp19339;
  assign tmp19326 = ~(s7 ? tmp19327 : tmp19335);
  assign tmp19325 = s8 ? 1 : tmp19326;
  assign tmp19324 = s9 ? tmp19325 : tmp19326;
  assign tmp19347 = s7 ? tmp19327 : tmp19335;
  assign tmp19346 = s8 ? tmp19347 : tmp19327;
  assign tmp19350 = ~(s6 ? tmp19336 : tmp19339);
  assign tmp19349 = s7 ? 1 : tmp19350;
  assign tmp19348 = ~(s8 ? tmp19349 : tmp19350);
  assign tmp19345 = ~(s9 ? tmp19346 : tmp19348);
  assign tmp19323 = s10 ? tmp19324 : tmp19345;
  assign tmp19322 = s12 ? tmp19323 : 0;
  assign tmp19359 = ~(l2 ? tmp18208 : 0);
  assign tmp19358 = l1 ? 1 : tmp19359;
  assign tmp19362 = s0 ? tmp19358 : 0;
  assign tmp19361 = s2 ? tmp19358 : tmp19362;
  assign tmp19365 = s0 ? 1 : tmp19358;
  assign tmp19364 = s1 ? tmp19358 : tmp19365;
  assign tmp19363 = s2 ? tmp18508 : tmp19364;
  assign tmp19360 = s3 ? tmp19361 : tmp19363;
  assign tmp19357 = s4 ? tmp19358 : tmp19360;
  assign tmp19371 = s0 ? tmp19358 : 1;
  assign tmp19370 = s1 ? 1 : tmp19371;
  assign tmp19369 = s2 ? tmp19358 : tmp19370;
  assign tmp19368 = s3 ? tmp19358 : tmp19369;
  assign tmp19374 = s1 ? tmp19365 : tmp18375;
  assign tmp19375 = s1 ? tmp18375 : tmp19358;
  assign tmp19373 = s2 ? tmp19374 : tmp19375;
  assign tmp19377 = s1 ? tmp19371 : 1;
  assign tmp19376 = s2 ? tmp19377 : 1;
  assign tmp19372 = s3 ? tmp19373 : tmp19376;
  assign tmp19367 = s4 ? tmp19368 : tmp19372;
  assign tmp19380 = s2 ? tmp19377 : tmp19365;
  assign tmp19379 = s3 ? tmp19380 : 1;
  assign tmp19383 = s1 ? tmp19365 : tmp19371;
  assign tmp19382 = s2 ? 1 : tmp19383;
  assign tmp19381 = s3 ? tmp19382 : 1;
  assign tmp19378 = s4 ? tmp19379 : tmp19381;
  assign tmp19366 = s5 ? tmp19367 : tmp19378;
  assign tmp19356 = s6 ? tmp19357 : tmp19366;
  assign tmp19388 = s1 ? tmp19362 : tmp18497;
  assign tmp19387 = s2 ? tmp19358 : tmp19388;
  assign tmp19389 = s2 ? tmp18529 : tmp19364;
  assign tmp19386 = s3 ? tmp19387 : tmp19389;
  assign tmp19385 = s4 ? tmp19358 : tmp19386;
  assign tmp19393 = s2 ? tmp19374 : tmp19358;
  assign tmp19392 = s3 ? tmp19393 : tmp19376;
  assign tmp19391 = s4 ? tmp19368 : tmp19392;
  assign tmp19397 = s1 ? tmp19358 : 1;
  assign tmp19396 = s2 ? tmp19377 : tmp19397;
  assign tmp19395 = s3 ? tmp19396 : 1;
  assign tmp19399 = s2 ? 1 : tmp19358;
  assign tmp19398 = s3 ? tmp19399 : 1;
  assign tmp19394 = s4 ? tmp19395 : tmp19398;
  assign tmp19390 = s5 ? tmp19391 : tmp19394;
  assign tmp19384 = s6 ? tmp19385 : tmp19390;
  assign tmp19355 = s7 ? tmp19356 : tmp19384;
  assign tmp19405 = s2 ? tmp18497 : tmp18506;
  assign tmp19404 = s3 ? tmp19405 : tmp18507;
  assign tmp19403 = s4 ? tmp18497 : tmp19404;
  assign tmp19409 = s2 ? tmp18497 : tmp18913;
  assign tmp19408 = s3 ? tmp18497 : tmp19409;
  assign tmp19412 = s1 ? tmp18375 : tmp18497;
  assign tmp19411 = s2 ? tmp18526 : tmp19412;
  assign tmp19413 = s2 ? tmp18533 : 1;
  assign tmp19410 = s3 ? tmp19411 : tmp19413;
  assign tmp19407 = s4 ? tmp19408 : tmp19410;
  assign tmp19406 = s5 ? tmp19407 : tmp18530;
  assign tmp19402 = s6 ? tmp19403 : tmp19406;
  assign tmp19417 = s2 ? tmp18497 : tmp18542;
  assign tmp19416 = s3 ? tmp19417 : tmp18543;
  assign tmp19415 = s4 ? tmp18497 : tmp19416;
  assign tmp19420 = s3 ? tmp18552 : tmp19413;
  assign tmp19419 = s4 ? tmp19408 : tmp19420;
  assign tmp19424 = s1 ? tmp18497 : tmp18534;
  assign tmp19423 = s2 ? 1 : tmp19424;
  assign tmp19422 = s3 ? tmp19423 : 1;
  assign tmp19421 = s4 ? tmp18531 : tmp19422;
  assign tmp19418 = s5 ? tmp19419 : tmp19421;
  assign tmp19414 = s6 ? tmp19415 : tmp19418;
  assign tmp19401 = s7 ? tmp19402 : tmp19414;
  assign tmp19400 = s8 ? tmp19355 : tmp19401;
  assign tmp19354 = s9 ? tmp19355 : tmp19400;
  assign tmp19426 = s8 ? tmp19355 : tmp19356;
  assign tmp19432 = s2 ? tmp18433 : tmp18478;
  assign tmp19431 = s3 ? tmp19432 : tmp18479;
  assign tmp19430 = s4 ? tmp18433 : tmp19431;
  assign tmp19435 = s3 ? tmp18433 : tmp18485;
  assign tmp19434 = s4 ? tmp19435 : tmp18487;
  assign tmp19433 = s5 ? tmp19434 : tmp18637;
  assign tmp19429 = s6 ? tmp19430 : tmp19433;
  assign tmp19438 = s4 ? tmp18531 : tmp18633;
  assign tmp19437 = s5 ? tmp19419 : tmp19438;
  assign tmp19436 = s6 ? tmp19415 : tmp19437;
  assign tmp19428 = s7 ? tmp19429 : tmp19436;
  assign tmp19427 = s8 ? tmp19428 : tmp19384;
  assign tmp19425 = s9 ? tmp19426 : tmp19427;
  assign tmp19353 = s10 ? tmp19354 : tmp19425;
  assign tmp19442 = s7 ? tmp19429 : tmp19414;
  assign tmp19441 = s8 ? tmp19442 : tmp19384;
  assign tmp19440 = s9 ? tmp19426 : tmp19441;
  assign tmp19439 = s10 ? tmp19354 : tmp19440;
  assign tmp19352 = s11 ? tmp19353 : tmp19439;
  assign tmp19351 = ~(s12 ? tmp19352 : 1);
  assign tmp19321 = s13 ? tmp19322 : tmp19351;
  assign tmp19064 = s14 ? tmp19065 : tmp19321;
  assign tmp19454 = s2 ? tmp18792 : tmp18795;
  assign tmp19453 = s3 ? tmp18791 : tmp19454;
  assign tmp19452 = s4 ? tmp19453 : tmp18797;
  assign tmp19458 = s2 ? tmp18822 : tmp18792;
  assign tmp19457 = s3 ? tmp19458 : tmp18824;
  assign tmp19456 = s4 ? tmp19457 : tmp18827;
  assign tmp19455 = s5 ? tmp18804 : tmp19456;
  assign tmp19451 = s6 ? tmp19452 : tmp19455;
  assign tmp19460 = s4 ? tmp19453 : tmp18837;
  assign tmp19465 = s1 ? tmp18792 : 1;
  assign tmp19464 = s2 ? tmp18809 : tmp19465;
  assign tmp19463 = s3 ? tmp19464 : tmp18852;
  assign tmp19462 = s4 ? tmp19463 : tmp18792;
  assign tmp19461 = s5 ? tmp18841 : tmp19462;
  assign tmp19459 = s6 ? tmp19460 : tmp19461;
  assign tmp19450 = s7 ? tmp19451 : tmp19459;
  assign tmp19449 = s8 ? tmp18787 : tmp19450;
  assign tmp19448 = s9 ? tmp18787 : tmp19449;
  assign tmp19469 = s6 ? tmp19452 : tmp18803;
  assign tmp19470 = s6 ? tmp19460 : tmp18840;
  assign tmp19468 = s7 ? tmp19469 : tmp19470;
  assign tmp19467 = s8 ? tmp19468 : tmp19469;
  assign tmp19472 = s7 ? tmp18887 : tmp19459;
  assign tmp19473 = s6 ? tmp19460 : tmp18888;
  assign tmp19471 = s8 ? tmp19472 : tmp19473;
  assign tmp19466 = s9 ? tmp19467 : tmp19471;
  assign tmp19447 = s10 ? tmp19448 : tmp19466;
  assign tmp19477 = s7 ? tmp18835 : tmp19459;
  assign tmp19476 = s8 ? tmp19477 : tmp19470;
  assign tmp19475 = s9 ? tmp19467 : tmp19476;
  assign tmp19474 = s10 ? tmp19448 : tmp19475;
  assign tmp19446 = s11 ? tmp19447 : tmp19474;
  assign tmp19445 = s12 ? 1 : tmp19446;
  assign tmp19444 = ~(s13 ? tmp19445 : tmp18895);
  assign tmp19443 = s14 ? tmp18644 : tmp19444;
  assign tmp19063 = s15 ? tmp19064 : tmp19443;
  assign tmp18194 = s16 ? tmp18195 : tmp19063;
  assign tmp19485 = s8 ? tmp19070 : tmp18344;
  assign tmp19484 = s9 ? tmp19069 : tmp19485;
  assign tmp19488 = s7 ? tmp19195 : tmp18403;
  assign tmp19487 = s8 ? tmp18409 : tmp19488;
  assign tmp19486 = s9 ? tmp18401 : tmp19487;
  assign tmp19483 = s10 ? tmp19484 : tmp19486;
  assign tmp19492 = s7 ? tmp19081 : tmp18403;
  assign tmp19491 = s8 ? tmp18420 : tmp19492;
  assign tmp19490 = s9 ? tmp18401 : tmp19491;
  assign tmp19489 = s10 ? tmp19484 : tmp19490;
  assign tmp19482 = s11 ? tmp19483 : tmp19489;
  assign tmp19498 = s7 ? tmp19219 : tmp19302;
  assign tmp19497 = s8 ? tmp19242 : tmp19498;
  assign tmp19496 = s9 ? tmp19217 : tmp19497;
  assign tmp19500 = s8 ? tmp19498 : tmp19219;
  assign tmp19502 = s7 ? tmp19312 : tmp19302;
  assign tmp19501 = s8 ? tmp19302 : tmp19502;
  assign tmp19499 = s9 ? tmp19500 : tmp19501;
  assign tmp19495 = s10 ? tmp19496 : tmp19499;
  assign tmp19506 = s7 ? tmp19234 : tmp19302;
  assign tmp19507 = s7 ? tmp19251 : tmp19302;
  assign tmp19505 = s8 ? tmp19506 : tmp19507;
  assign tmp19504 = s9 ? tmp19500 : tmp19505;
  assign tmp19503 = s10 ? tmp19496 : tmp19504;
  assign tmp19494 = s11 ? tmp19495 : tmp19503;
  assign tmp19493 = s12 ? 1 : tmp19494;
  assign tmp19481 = s13 ? tmp19482 : tmp19493;
  assign tmp19512 = ~(s8 ? tmp19347 : 0);
  assign tmp19511 = s9 ? tmp19325 : tmp19512;
  assign tmp19515 = ~(s7 ? tmp19335 : 0);
  assign tmp19514 = s8 ? 1 : tmp19515;
  assign tmp19513 = s9 ? 1 : tmp19514;
  assign tmp19510 = s10 ? tmp19511 : tmp19513;
  assign tmp19509 = s12 ? tmp19510 : 0;
  assign tmp19526 = s1 ? tmp19358 : tmp19371;
  assign tmp19525 = s2 ? 1 : tmp19526;
  assign tmp19524 = s3 ? tmp19525 : 1;
  assign tmp19523 = s4 ? tmp19379 : tmp19524;
  assign tmp19522 = s5 ? tmp19391 : tmp19523;
  assign tmp19521 = s6 ? tmp19385 : tmp19522;
  assign tmp19520 = s7 ? tmp19356 : tmp19521;
  assign tmp19530 = s4 ? tmp18361 : tmp18565;
  assign tmp19535 = s1 ? 1 : tmp18375;
  assign tmp19534 = s2 ? tmp18361 : tmp19535;
  assign tmp19533 = s3 ? tmp18361 : tmp19534;
  assign tmp19536 = s3 ? tmp18579 : tmp19117;
  assign tmp19532 = s4 ? tmp19533 : tmp19536;
  assign tmp19539 = s2 ? tmp18374 : tmp18377;
  assign tmp19538 = s3 ? tmp19539 : 1;
  assign tmp19541 = s2 ? 1 : tmp18580;
  assign tmp19540 = s3 ? tmp19541 : 1;
  assign tmp19537 = s4 ? tmp19538 : tmp19540;
  assign tmp19531 = s5 ? tmp19532 : tmp19537;
  assign tmp19529 = s6 ? tmp19530 : tmp19531;
  assign tmp19543 = s4 ? tmp18361 : tmp18593;
  assign tmp19546 = s3 ? tmp18603 : tmp19117;
  assign tmp19545 = s4 ? tmp19533 : tmp19546;
  assign tmp19549 = s2 ? 1 : tmp18394;
  assign tmp19548 = s3 ? tmp19549 : 1;
  assign tmp19547 = s4 ? tmp18396 : tmp19548;
  assign tmp19544 = s5 ? tmp19545 : tmp19547;
  assign tmp19542 = s6 ? tmp19543 : tmp19544;
  assign tmp19528 = s7 ? tmp19529 : tmp19542;
  assign tmp19527 = s8 ? tmp19520 : tmp19528;
  assign tmp19519 = s9 ? tmp19520 : tmp19527;
  assign tmp19556 = s2 ? tmp18433 : tmp18437;
  assign tmp19555 = s3 ? tmp19556 : tmp18444;
  assign tmp19554 = s4 ? tmp18433 : tmp19555;
  assign tmp19561 = s1 ? tmp18375 : tmp18433;
  assign tmp19560 = s2 ? tmp18464 : tmp19561;
  assign tmp19559 = s3 ? tmp19560 : tmp18466;
  assign tmp19558 = s4 ? tmp19435 : tmp19559;
  assign tmp19557 = s5 ? tmp19558 : tmp18468;
  assign tmp19553 = s6 ? tmp19554 : tmp19557;
  assign tmp19563 = s5 ? tmp19434 : tmp18613;
  assign tmp19562 = s6 ? tmp19430 : tmp19563;
  assign tmp19552 = s7 ? tmp19553 : tmp19562;
  assign tmp19551 = s8 ? tmp19552 : tmp19553;
  assign tmp19567 = s4 ? tmp19379 : tmp19398;
  assign tmp19566 = s5 ? tmp19391 : tmp19567;
  assign tmp19565 = s6 ? tmp19385 : tmp19566;
  assign tmp19564 = s7 ? tmp19565 : tmp19429;
  assign tmp19550 = s9 ? tmp19551 : tmp19564;
  assign tmp19518 = s10 ? tmp19519 : tmp19550;
  assign tmp19570 = s7 ? tmp19521 : tmp19562;
  assign tmp19569 = s9 ? tmp19551 : tmp19570;
  assign tmp19568 = s10 ? tmp19519 : tmp19569;
  assign tmp19517 = s11 ? tmp19518 : tmp19568;
  assign tmp19516 = ~(s12 ? tmp19517 : 1);
  assign tmp19508 = s13 ? tmp19509 : tmp19516;
  assign tmp19480 = s14 ? tmp19481 : tmp19508;
  assign tmp19577 = s8 ? tmp18787 : tmp18874;
  assign tmp19576 = s9 ? tmp18787 : tmp19577;
  assign tmp19580 = s7 ? tmp18887 : tmp18881;
  assign tmp19579 = s8 ? tmp18886 : tmp19580;
  assign tmp19578 = s9 ? tmp18879 : tmp19579;
  assign tmp19575 = s10 ? tmp19576 : tmp19578;
  assign tmp19584 = s7 ? tmp18835 : tmp18881;
  assign tmp19583 = s8 ? tmp18894 : tmp19584;
  assign tmp19582 = s9 ? tmp18879 : tmp19583;
  assign tmp19581 = s10 ? tmp19576 : tmp19582;
  assign tmp19574 = s11 ? tmp19575 : tmp19581;
  assign tmp19573 = s12 ? 1 : tmp19574;
  assign tmp19572 = ~(s13 ? tmp19573 : tmp18895);
  assign tmp19571 = s14 ? tmp18644 : tmp19572;
  assign tmp19479 = s15 ? tmp19480 : tmp19571;
  assign tmp19592 = s8 ? tmp19520 : tmp19401;
  assign tmp19591 = s9 ? tmp19520 : tmp19592;
  assign tmp19594 = s8 ? tmp19520 : tmp19356;
  assign tmp19593 = s9 ? tmp19594 : tmp19565;
  assign tmp19590 = s10 ? tmp19591 : tmp19593;
  assign tmp19596 = s9 ? tmp19594 : tmp19521;
  assign tmp19595 = s10 ? tmp19591 : tmp19596;
  assign tmp19589 = s11 ? tmp19590 : tmp19595;
  assign tmp19588 = ~(s12 ? tmp19589 : 1);
  assign tmp19587 = s13 ? tmp19322 : tmp19588;
  assign tmp19586 = s14 ? tmp19065 : tmp19587;
  assign tmp19585 = s15 ? tmp19586 : tmp19443;
  assign tmp19478 = s16 ? tmp19479 : tmp19585;
  assign tmp18193 = s17 ? tmp18194 : tmp19478;
  assign s14n = tmp18193;

  assign tmp19612 = ~(l2 ? 1 : 0);
  assign tmp19611 = l1 ? 1 : tmp19612;
  assign tmp19614 = l1 ? 1 : 0;
  assign tmp19613 = s0 ? tmp19614 : tmp19611;
  assign tmp19610 = s1 ? tmp19611 : tmp19613;
  assign tmp19617 = s0 ? tmp19611 : tmp19614;
  assign tmp19616 = s1 ? tmp19617 : tmp19611;
  assign tmp19615 = s2 ? tmp19611 : tmp19616;
  assign tmp19609 = s3 ? tmp19610 : tmp19615;
  assign tmp19621 = s0 ? tmp19611 : 1;
  assign tmp19622 = s0 ? tmp19614 : 1;
  assign tmp19620 = s1 ? tmp19621 : tmp19622;
  assign tmp19619 = s2 ? tmp19616 : tmp19620;
  assign tmp19624 = s1 ? tmp19614 : 1;
  assign tmp19626 = s0 ? tmp19611 : tmp19612;
  assign tmp19627 = s0 ? 1 : tmp19611;
  assign tmp19625 = s1 ? tmp19626 : tmp19627;
  assign tmp19623 = s2 ? tmp19624 : tmp19625;
  assign tmp19618 = s3 ? tmp19619 : tmp19623;
  assign tmp19608 = s4 ? tmp19609 : tmp19618;
  assign tmp19632 = s1 ? tmp19617 : tmp19613;
  assign tmp19635 = l2 ? 1 : 0;
  assign tmp19634 = ~(s0 ? tmp19635 : 1);
  assign tmp19633 = s1 ? tmp19613 : tmp19634;
  assign tmp19631 = s2 ? tmp19632 : tmp19633;
  assign tmp19637 = s0 ? 1 : tmp19635;
  assign tmp19638 = ~(s1 ? 1 : tmp19621);
  assign tmp19636 = ~(s2 ? tmp19637 : tmp19638);
  assign tmp19630 = s3 ? tmp19631 : tmp19636;
  assign tmp19641 = s1 ? tmp19627 : tmp19622;
  assign tmp19642 = s1 ? tmp19622 : tmp19617;
  assign tmp19640 = s2 ? tmp19641 : tmp19642;
  assign tmp19644 = s1 ? tmp19635 : 0;
  assign tmp19643 = ~(s2 ? tmp19644 : 0);
  assign tmp19639 = s3 ? tmp19640 : tmp19643;
  assign tmp19629 = s4 ? tmp19630 : tmp19639;
  assign tmp19649 = s0 ? tmp19635 : 0;
  assign tmp19648 = s1 ? tmp19649 : 0;
  assign tmp19651 = s0 ? 1 : tmp19612;
  assign tmp19650 = ~(s1 ? tmp19651 : tmp19612);
  assign tmp19647 = s2 ? tmp19648 : tmp19650;
  assign tmp19646 = s3 ? tmp19647 : 0;
  assign tmp19654 = s1 ? tmp19651 : tmp19612;
  assign tmp19653 = s2 ? 1 : tmp19654;
  assign tmp19652 = ~(s3 ? tmp19653 : 1);
  assign tmp19645 = ~(s4 ? tmp19646 : tmp19652);
  assign tmp19628 = s5 ? tmp19629 : tmp19645;
  assign tmp19607 = s6 ? tmp19608 : tmp19628;
  assign tmp19659 = s1 ? tmp19621 : tmp19614;
  assign tmp19658 = s2 ? tmp19616 : tmp19659;
  assign tmp19657 = s3 ? tmp19658 : tmp19623;
  assign tmp19656 = s4 ? tmp19609 : tmp19657;
  assign tmp19664 = s1 ? tmp19611 : tmp19634;
  assign tmp19663 = s2 ? tmp19616 : tmp19664;
  assign tmp19665 = ~(s2 ? tmp19635 : tmp19638);
  assign tmp19662 = s3 ? tmp19663 : tmp19665;
  assign tmp19668 = s1 ? tmp19614 : tmp19617;
  assign tmp19667 = s2 ? tmp19641 : tmp19668;
  assign tmp19666 = s3 ? tmp19667 : tmp19643;
  assign tmp19661 = s4 ? tmp19662 : tmp19666;
  assign tmp19671 = s2 ? tmp19648 : tmp19644;
  assign tmp19670 = s3 ? tmp19671 : 0;
  assign tmp19673 = s2 ? 1 : tmp19612;
  assign tmp19672 = ~(s3 ? tmp19673 : 1);
  assign tmp19669 = ~(s4 ? tmp19670 : tmp19672);
  assign tmp19660 = s5 ? tmp19661 : tmp19669;
  assign tmp19655 = s6 ? tmp19656 : tmp19660;
  assign tmp19606 = s7 ? tmp19607 : tmp19655;
  assign tmp19679 = s1 ? tmp19611 : tmp19627;
  assign tmp19678 = s2 ? tmp19624 : tmp19679;
  assign tmp19677 = s3 ? tmp19619 : tmp19678;
  assign tmp19676 = s4 ? tmp19609 : tmp19677;
  assign tmp19684 = s1 ? tmp19613 : tmp19617;
  assign tmp19683 = s2 ? tmp19632 : tmp19684;
  assign tmp19687 = s0 ? tmp19614 : tmp19612;
  assign tmp19686 = s1 ? tmp19613 : tmp19687;
  assign tmp19688 = s1 ? 1 : tmp19621;
  assign tmp19685 = s2 ? tmp19686 : tmp19688;
  assign tmp19682 = s3 ? tmp19683 : tmp19685;
  assign tmp19690 = ~(s2 ? tmp19648 : 0);
  assign tmp19689 = s3 ? tmp19640 : tmp19690;
  assign tmp19681 = s4 ? tmp19682 : tmp19689;
  assign tmp19680 = s5 ? tmp19681 : tmp19645;
  assign tmp19675 = s6 ? tmp19676 : tmp19680;
  assign tmp19693 = s3 ? tmp19658 : tmp19678;
  assign tmp19692 = s4 ? tmp19609 : tmp19693;
  assign tmp19698 = s1 ? tmp19611 : tmp19617;
  assign tmp19697 = s2 ? tmp19616 : tmp19698;
  assign tmp19700 = s1 ? tmp19611 : tmp19612;
  assign tmp19699 = s2 ? tmp19700 : tmp19688;
  assign tmp19696 = s3 ? tmp19697 : tmp19699;
  assign tmp19702 = s2 ? tmp19641 : tmp19611;
  assign tmp19701 = s3 ? tmp19702 : tmp19690;
  assign tmp19695 = s4 ? tmp19696 : tmp19701;
  assign tmp19694 = s5 ? tmp19695 : tmp19669;
  assign tmp19691 = s6 ? tmp19692 : tmp19694;
  assign tmp19674 = s7 ? tmp19675 : tmp19691;
  assign tmp19605 = s8 ? tmp19606 : tmp19674;
  assign tmp19708 = s2 ? tmp19614 : tmp19622;
  assign tmp19711 = s0 ? 1 : tmp19614;
  assign tmp19710 = s1 ? tmp19614 : tmp19711;
  assign tmp19709 = s2 ? tmp19624 : tmp19710;
  assign tmp19707 = s3 ? tmp19708 : tmp19709;
  assign tmp19706 = s4 ? tmp19614 : tmp19707;
  assign tmp19717 = s0 ? tmp19614 : 0;
  assign tmp19716 = s1 ? tmp19614 : tmp19717;
  assign tmp19715 = s2 ? tmp19614 : tmp19716;
  assign tmp19720 = ~(l1 ? 1 : 0);
  assign tmp19719 = s0 ? 1 : tmp19720;
  assign tmp19721 = ~(s1 ? 1 : tmp19622);
  assign tmp19718 = ~(s2 ? tmp19719 : tmp19721);
  assign tmp19714 = s3 ? tmp19715 : tmp19718;
  assign tmp19724 = s1 ? tmp19711 : tmp19622;
  assign tmp19725 = s1 ? tmp19622 : tmp19614;
  assign tmp19723 = s2 ? tmp19724 : tmp19725;
  assign tmp19726 = s2 ? tmp19614 : 1;
  assign tmp19722 = s3 ? tmp19723 : tmp19726;
  assign tmp19713 = s4 ? tmp19714 : tmp19722;
  assign tmp19730 = s1 ? tmp19622 : 1;
  assign tmp19731 = s1 ? tmp19711 : tmp19614;
  assign tmp19729 = s2 ? tmp19730 : tmp19731;
  assign tmp19728 = s3 ? tmp19729 : 1;
  assign tmp19733 = s2 ? 1 : tmp19731;
  assign tmp19732 = s3 ? tmp19733 : 1;
  assign tmp19727 = s4 ? tmp19728 : tmp19732;
  assign tmp19712 = s5 ? tmp19713 : tmp19727;
  assign tmp19705 = s6 ? tmp19706 : tmp19712;
  assign tmp19739 = s1 ? 1 : tmp19622;
  assign tmp19738 = s2 ? tmp19614 : tmp19739;
  assign tmp19737 = s3 ? tmp19715 : tmp19738;
  assign tmp19741 = s2 ? tmp19724 : tmp19614;
  assign tmp19742 = s2 ? tmp19624 : 1;
  assign tmp19740 = s3 ? tmp19741 : tmp19742;
  assign tmp19736 = s4 ? tmp19737 : tmp19740;
  assign tmp19745 = s2 ? tmp19730 : tmp19624;
  assign tmp19744 = s3 ? tmp19745 : 1;
  assign tmp19747 = s2 ? 1 : tmp19614;
  assign tmp19746 = s3 ? tmp19747 : 1;
  assign tmp19743 = s4 ? tmp19744 : tmp19746;
  assign tmp19735 = s5 ? tmp19736 : tmp19743;
  assign tmp19734 = s6 ? tmp19706 : tmp19735;
  assign tmp19704 = s7 ? tmp19705 : tmp19734;
  assign tmp19703 = s8 ? tmp19674 : tmp19704;
  assign tmp19604 = s9 ? tmp19605 : tmp19703;
  assign tmp19754 = s3 ? tmp19702 : tmp19643;
  assign tmp19753 = s4 ? tmp19662 : tmp19754;
  assign tmp19752 = s5 ? tmp19753 : tmp19669;
  assign tmp19751 = s6 ? tmp19656 : tmp19752;
  assign tmp19750 = s7 ? tmp19607 : tmp19751;
  assign tmp19749 = s8 ? tmp19750 : tmp19607;
  assign tmp19762 = s1 ? tmp19614 : tmp19611;
  assign tmp19761 = s2 ? tmp19641 : tmp19762;
  assign tmp19760 = s3 ? tmp19761 : tmp19643;
  assign tmp19759 = s4 ? tmp19662 : tmp19760;
  assign tmp19758 = s5 ? tmp19759 : tmp19669;
  assign tmp19757 = s6 ? tmp19656 : tmp19758;
  assign tmp19756 = s7 ? tmp19757 : tmp19734;
  assign tmp19763 = s7 ? tmp19691 : tmp19751;
  assign tmp19755 = s8 ? tmp19756 : tmp19763;
  assign tmp19748 = s9 ? tmp19749 : tmp19755;
  assign tmp19603 = s10 ? tmp19604 : tmp19748;
  assign tmp19767 = s7 ? tmp19655 : tmp19734;
  assign tmp19766 = s8 ? tmp19767 : tmp19763;
  assign tmp19765 = s9 ? tmp19749 : tmp19766;
  assign tmp19764 = s10 ? tmp19604 : tmp19765;
  assign tmp19602 = s11 ? tmp19603 : tmp19764;
  assign tmp19777 = s2 ? tmp19611 : tmp19621;
  assign tmp19780 = s0 ? 1 : 0;
  assign tmp19779 = s1 ? tmp19611 : tmp19780;
  assign tmp19783 = ~(l1 ? 1 : tmp19612);
  assign tmp19782 = ~(s0 ? 1 : tmp19783);
  assign tmp19781 = s1 ? tmp19611 : tmp19782;
  assign tmp19778 = s2 ? tmp19779 : tmp19781;
  assign tmp19776 = s3 ? tmp19777 : tmp19778;
  assign tmp19775 = s4 ? tmp19611 : tmp19776;
  assign tmp19789 = ~(s0 ? tmp19614 : 0);
  assign tmp19788 = s1 ? 1 : tmp19789;
  assign tmp19787 = ~(s2 ? tmp19635 : tmp19788);
  assign tmp19786 = s3 ? tmp19611 : tmp19787;
  assign tmp19792 = s1 ? tmp19719 : tmp19789;
  assign tmp19793 = ~(s1 ? tmp19717 : tmp19614);
  assign tmp19791 = s2 ? tmp19792 : tmp19793;
  assign tmp19790 = ~(s3 ? tmp19791 : 1);
  assign tmp19785 = s4 ? tmp19786 : tmp19790;
  assign tmp19784 = s5 ? tmp19785 : 0;
  assign tmp19774 = s6 ? tmp19775 : tmp19784;
  assign tmp19798 = s2 ? tmp19792 : tmp19720;
  assign tmp19797 = ~(s3 ? tmp19798 : 1);
  assign tmp19796 = s4 ? tmp19786 : tmp19797;
  assign tmp19795 = s5 ? tmp19796 : 0;
  assign tmp19794 = s6 ? tmp19775 : tmp19795;
  assign tmp19773 = s7 ? tmp19774 : tmp19794;
  assign tmp19806 = ~(s0 ? tmp19614 : 1);
  assign tmp19805 = ~(s1 ? 1 : tmp19806);
  assign tmp19804 = s2 ? tmp19611 : tmp19805;
  assign tmp19803 = s3 ? tmp19611 : tmp19804;
  assign tmp19809 = s1 ? tmp19719 : tmp19806;
  assign tmp19810 = ~(s1 ? tmp19622 : tmp19614);
  assign tmp19808 = s2 ? tmp19809 : tmp19810;
  assign tmp19813 = ~(s0 ? 1 : 0);
  assign tmp19812 = s1 ? tmp19780 : tmp19813;
  assign tmp19811 = s2 ? tmp19812 : 1;
  assign tmp19807 = ~(s3 ? tmp19808 : tmp19811);
  assign tmp19802 = s4 ? tmp19803 : tmp19807;
  assign tmp19801 = s5 ? tmp19802 : 0;
  assign tmp19800 = s6 ? tmp19775 : tmp19801;
  assign tmp19818 = s1 ? tmp19611 : 0;
  assign tmp19817 = s2 ? tmp19818 : tmp19781;
  assign tmp19816 = s3 ? tmp19777 : tmp19817;
  assign tmp19815 = s4 ? tmp19611 : tmp19816;
  assign tmp19822 = s2 ? tmp19809 : tmp19720;
  assign tmp19824 = s1 ? tmp19780 : 1;
  assign tmp19823 = s2 ? tmp19824 : 1;
  assign tmp19821 = ~(s3 ? tmp19822 : tmp19823);
  assign tmp19820 = s4 ? tmp19803 : tmp19821;
  assign tmp19819 = s5 ? tmp19820 : 0;
  assign tmp19814 = s6 ? tmp19815 : tmp19819;
  assign tmp19799 = s7 ? tmp19800 : tmp19814;
  assign tmp19772 = s8 ? tmp19773 : tmp19799;
  assign tmp19830 = ~(s3 ? tmp19808 : 1);
  assign tmp19829 = s4 ? tmp19786 : tmp19830;
  assign tmp19828 = s5 ? tmp19829 : 0;
  assign tmp19827 = s6 ? tmp19775 : tmp19828;
  assign tmp19834 = ~(s3 ? tmp19822 : 1);
  assign tmp19833 = s4 ? tmp19786 : tmp19834;
  assign tmp19832 = s5 ? tmp19833 : 0;
  assign tmp19831 = s6 ? tmp19815 : tmp19832;
  assign tmp19826 = s7 ? tmp19827 : tmp19831;
  assign tmp19825 = s8 ? tmp19799 : tmp19826;
  assign tmp19771 = s9 ? tmp19772 : tmp19825;
  assign tmp19836 = s8 ? tmp19826 : tmp19827;
  assign tmp19844 = s1 ? tmp19614 : tmp19612;
  assign tmp19843 = s2 ? tmp19611 : tmp19844;
  assign tmp19846 = s1 ? tmp19635 : 1;
  assign tmp19845 = ~(s2 ? tmp19846 : tmp19788);
  assign tmp19842 = s3 ? tmp19843 : tmp19845;
  assign tmp19841 = s4 ? tmp19842 : tmp19797;
  assign tmp19840 = s5 ? tmp19841 : 0;
  assign tmp19839 = s6 ? tmp19815 : tmp19840;
  assign tmp19850 = s3 ? tmp19843 : tmp19787;
  assign tmp19849 = s4 ? tmp19850 : tmp19834;
  assign tmp19848 = s5 ? tmp19849 : 0;
  assign tmp19847 = s6 ? tmp19815 : tmp19848;
  assign tmp19838 = s7 ? tmp19839 : tmp19847;
  assign tmp19856 = s2 ? tmp19611 : tmp19762;
  assign tmp19855 = s3 ? tmp19856 : tmp19804;
  assign tmp19854 = s4 ? tmp19855 : tmp19821;
  assign tmp19853 = s5 ? tmp19854 : 0;
  assign tmp19852 = s6 ? tmp19815 : tmp19853;
  assign tmp19851 = s7 ? tmp19852 : tmp19847;
  assign tmp19837 = s8 ? tmp19838 : tmp19851;
  assign tmp19835 = s9 ? tmp19836 : tmp19837;
  assign tmp19770 = s10 ? tmp19771 : tmp19835;
  assign tmp19860 = s7 ? tmp19794 : tmp19831;
  assign tmp19861 = s7 ? tmp19814 : tmp19831;
  assign tmp19859 = s8 ? tmp19860 : tmp19861;
  assign tmp19858 = s9 ? tmp19836 : tmp19859;
  assign tmp19857 = s10 ? tmp19771 : tmp19858;
  assign tmp19769 = s11 ? tmp19770 : tmp19857;
  assign tmp19768 = s12 ? tmp19769 : 1;
  assign tmp19601 = s13 ? tmp19602 : tmp19768;
  assign tmp19872 = s2 ? tmp19635 : tmp19649;
  assign tmp19874 = s1 ? tmp19635 : tmp19813;
  assign tmp19875 = s1 ? tmp19635 : tmp19637;
  assign tmp19873 = s2 ? tmp19874 : tmp19875;
  assign tmp19871 = s3 ? tmp19872 : tmp19873;
  assign tmp19870 = s4 ? tmp19635 : tmp19871;
  assign tmp19879 = s2 ? tmp19635 : 1;
  assign tmp19878 = s3 ? tmp19635 : tmp19879;
  assign tmp19877 = s4 ? tmp19878 : 1;
  assign tmp19876 = s5 ? tmp19877 : 1;
  assign tmp19869 = s6 ? tmp19870 : tmp19876;
  assign tmp19883 = s2 ? tmp19846 : tmp19875;
  assign tmp19882 = s3 ? tmp19872 : tmp19883;
  assign tmp19881 = s4 ? tmp19635 : tmp19882;
  assign tmp19888 = s1 ? 1 : tmp19635;
  assign tmp19887 = s2 ? tmp19635 : tmp19888;
  assign tmp19886 = s3 ? tmp19887 : tmp19879;
  assign tmp19885 = s4 ? tmp19886 : 1;
  assign tmp19884 = s5 ? tmp19885 : 1;
  assign tmp19880 = s6 ? tmp19881 : tmp19884;
  assign tmp19868 = s7 ? tmp19869 : tmp19880;
  assign tmp19896 = s0 ? tmp19635 : 1;
  assign tmp19895 = s1 ? tmp19896 : tmp19635;
  assign tmp19894 = s2 ? tmp19635 : tmp19895;
  assign tmp19893 = s3 ? tmp19894 : tmp19879;
  assign tmp19892 = s4 ? tmp19893 : 1;
  assign tmp19891 = s5 ? tmp19892 : 1;
  assign tmp19890 = s6 ? tmp19870 : tmp19891;
  assign tmp19889 = s7 ? tmp19890 : tmp19880;
  assign tmp19867 = s8 ? tmp19868 : tmp19889;
  assign tmp19866 = s9 ? tmp19867 : tmp19889;
  assign tmp19898 = s8 ? tmp19889 : tmp19890;
  assign tmp19905 = s2 ? tmp19846 : 1;
  assign tmp19904 = s3 ? tmp19887 : tmp19905;
  assign tmp19903 = s4 ? tmp19904 : 1;
  assign tmp19902 = s5 ? tmp19903 : 1;
  assign tmp19901 = s6 ? tmp19881 : tmp19902;
  assign tmp19900 = s7 ? tmp19901 : tmp19880;
  assign tmp19899 = s8 ? tmp19900 : tmp19880;
  assign tmp19897 = s9 ? tmp19898 : tmp19899;
  assign tmp19865 = s10 ? tmp19866 : tmp19897;
  assign tmp19907 = s9 ? tmp19898 : tmp19880;
  assign tmp19906 = s10 ? tmp19866 : tmp19907;
  assign tmp19864 = s11 ? tmp19865 : tmp19906;
  assign tmp19917 = ~(s0 ? tmp19614 : tmp19612);
  assign tmp19916 = s1 ? tmp19635 : tmp19917;
  assign tmp19919 = s1 ? tmp19649 : tmp19635;
  assign tmp19918 = s2 ? tmp19635 : tmp19919;
  assign tmp19915 = s3 ? tmp19916 : tmp19918;
  assign tmp19922 = s1 ? tmp19649 : tmp19806;
  assign tmp19921 = s2 ? tmp19919 : tmp19922;
  assign tmp19924 = s1 ? tmp19614 : tmp19780;
  assign tmp19925 = ~(s1 ? tmp19635 : tmp19637);
  assign tmp19923 = ~(s2 ? tmp19924 : tmp19925);
  assign tmp19920 = s3 ? tmp19921 : tmp19923;
  assign tmp19914 = s4 ? tmp19915 : tmp19920;
  assign tmp19928 = s3 ? tmp19647 : tmp19887;
  assign tmp19931 = s1 ? tmp19637 : tmp19720;
  assign tmp19933 = ~(s0 ? tmp19635 : 0);
  assign tmp19932 = ~(s1 ? tmp19614 : tmp19933);
  assign tmp19930 = s2 ? tmp19931 : tmp19932;
  assign tmp19934 = s2 ? tmp19916 : 1;
  assign tmp19929 = s3 ? tmp19930 : tmp19934;
  assign tmp19927 = s4 ? tmp19928 : tmp19929;
  assign tmp19938 = s1 ? tmp19896 : 1;
  assign tmp19939 = s1 ? tmp19780 : 0;
  assign tmp19937 = s2 ? tmp19938 : tmp19939;
  assign tmp19941 = ~(s1 ? 1 : tmp19637);
  assign tmp19940 = ~(s2 ? tmp19939 : tmp19941);
  assign tmp19936 = s3 ? tmp19937 : tmp19940;
  assign tmp19944 = s1 ? tmp19637 : 0;
  assign tmp19943 = s2 ? tmp19938 : tmp19944;
  assign tmp19946 = s1 ? 1 : tmp19637;
  assign tmp19947 = s1 ? tmp19637 : 1;
  assign tmp19945 = s2 ? tmp19946 : tmp19947;
  assign tmp19942 = s3 ? tmp19943 : tmp19945;
  assign tmp19935 = s4 ? tmp19936 : tmp19942;
  assign tmp19926 = s5 ? tmp19927 : tmp19935;
  assign tmp19913 = s6 ? tmp19914 : tmp19926;
  assign tmp19952 = s1 ? tmp19649 : tmp19720;
  assign tmp19951 = s2 ? tmp19919 : tmp19952;
  assign tmp19954 = s1 ? tmp19614 : 0;
  assign tmp19953 = ~(s2 ? tmp19954 : tmp19925);
  assign tmp19950 = s3 ? tmp19951 : tmp19953;
  assign tmp19949 = s4 ? tmp19915 : tmp19950;
  assign tmp19958 = s2 ? tmp19648 : tmp19635;
  assign tmp19957 = s3 ? tmp19958 : tmp19887;
  assign tmp19961 = ~(s1 ? tmp19614 : tmp19612);
  assign tmp19960 = s2 ? tmp19931 : tmp19961;
  assign tmp19959 = s3 ? tmp19960 : tmp19934;
  assign tmp19956 = s4 ? tmp19957 : tmp19959;
  assign tmp19964 = s2 ? tmp19938 : 0;
  assign tmp19965 = s2 ? 1 : tmp19888;
  assign tmp19963 = s3 ? tmp19964 : tmp19965;
  assign tmp19967 = s2 ? 1 : tmp19635;
  assign tmp19966 = s3 ? tmp19967 : tmp19888;
  assign tmp19962 = s4 ? tmp19963 : tmp19966;
  assign tmp19955 = s5 ? tmp19956 : tmp19962;
  assign tmp19948 = s6 ? tmp19949 : tmp19955;
  assign tmp19912 = s7 ? tmp19913 : tmp19948;
  assign tmp19974 = ~(s1 ? tmp19651 : tmp19933);
  assign tmp19973 = s2 ? tmp19648 : tmp19974;
  assign tmp19976 = ~(s1 ? 1 : tmp19635);
  assign tmp19975 = ~(s2 ? tmp19651 : tmp19976);
  assign tmp19972 = s3 ? tmp19973 : tmp19975;
  assign tmp19971 = s4 ? tmp19972 : tmp19929;
  assign tmp19970 = s5 ? tmp19971 : tmp19935;
  assign tmp19969 = s6 ? tmp19914 : tmp19970;
  assign tmp19982 = s1 ? tmp19635 : tmp19649;
  assign tmp19981 = s2 ? tmp19648 : tmp19982;
  assign tmp19980 = s3 ? tmp19981 : tmp19887;
  assign tmp19984 = s2 ? tmp19931 : tmp19635;
  assign tmp19983 = s3 ? tmp19984 : tmp19879;
  assign tmp19979 = s4 ? tmp19980 : tmp19983;
  assign tmp19978 = s5 ? tmp19979 : tmp19962;
  assign tmp19977 = s6 ? tmp19949 : tmp19978;
  assign tmp19968 = s7 ? tmp19969 : tmp19977;
  assign tmp19911 = s8 ? tmp19912 : tmp19968;
  assign tmp19990 = s2 ? tmp19614 : tmp19725;
  assign tmp19989 = s3 ? tmp19614 : tmp19990;
  assign tmp19994 = ~(s0 ? 1 : tmp19720);
  assign tmp19993 = s1 ? tmp19614 : tmp19994;
  assign tmp19992 = s2 ? tmp19924 : tmp19993;
  assign tmp19991 = s3 ? tmp19708 : tmp19992;
  assign tmp19988 = s4 ? tmp19989 : tmp19991;
  assign tmp19999 = ~(s1 ? 1 : tmp19720);
  assign tmp19998 = s2 ? tmp19614 : tmp19999;
  assign tmp19997 = s3 ? tmp19729 : tmp19998;
  assign tmp20002 = s1 ? tmp19719 : tmp19720;
  assign tmp20001 = s2 ? tmp20002 : tmp19720;
  assign tmp20003 = ~(s2 ? tmp19614 : 0);
  assign tmp20000 = ~(s3 ? tmp20001 : tmp20003);
  assign tmp19996 = s4 ? tmp19997 : tmp20000;
  assign tmp20007 = s1 ? tmp19717 : 0;
  assign tmp20008 = ~(s1 ? tmp19780 : 0);
  assign tmp20006 = s2 ? tmp20007 : tmp20008;
  assign tmp20010 = ~(s1 ? 1 : tmp19719);
  assign tmp20009 = s2 ? tmp19939 : tmp20010;
  assign tmp20005 = s3 ? tmp20006 : tmp20009;
  assign tmp20013 = ~(s1 ? tmp19719 : 0);
  assign tmp20012 = s2 ? tmp20007 : tmp20013;
  assign tmp20015 = s1 ? 1 : tmp19719;
  assign tmp20016 = s1 ? tmp19719 : 1;
  assign tmp20014 = ~(s2 ? tmp20015 : tmp20016);
  assign tmp20011 = s3 ? tmp20012 : tmp20014;
  assign tmp20004 = s4 ? tmp20005 : tmp20011;
  assign tmp19995 = s5 ? tmp19996 : tmp20004;
  assign tmp19987 = s6 ? tmp19988 : tmp19995;
  assign tmp20020 = s2 ? tmp19954 : tmp19993;
  assign tmp20019 = s3 ? tmp19708 : tmp20020;
  assign tmp20018 = s4 ? tmp19989 : tmp20019;
  assign tmp20024 = s2 ? tmp19730 : tmp19614;
  assign tmp20023 = s3 ? tmp20024 : tmp19998;
  assign tmp20022 = s4 ? tmp20023 : tmp20000;
  assign tmp20027 = s2 ? tmp20007 : 1;
  assign tmp20029 = s1 ? 1 : tmp19720;
  assign tmp20028 = ~(s2 ? 1 : tmp20029);
  assign tmp20026 = s3 ? tmp20027 : tmp20028;
  assign tmp20031 = s2 ? 1 : tmp19720;
  assign tmp20030 = ~(s3 ? tmp20031 : tmp20029);
  assign tmp20025 = s4 ? tmp20026 : tmp20030;
  assign tmp20021 = s5 ? tmp20022 : tmp20025;
  assign tmp20017 = s6 ? tmp20018 : tmp20021;
  assign tmp19986 = ~(s7 ? tmp19987 : tmp20017);
  assign tmp19985 = s8 ? tmp19968 : tmp19986;
  assign tmp19910 = s9 ? tmp19911 : tmp19985;
  assign tmp20037 = s4 ? tmp19957 : tmp19983;
  assign tmp20036 = s5 ? tmp20037 : tmp19962;
  assign tmp20035 = s6 ? tmp19949 : tmp20036;
  assign tmp20034 = s7 ? tmp19913 : tmp20035;
  assign tmp20033 = s8 ? tmp20034 : tmp19913;
  assign tmp20043 = s3 ? tmp19960 : tmp19879;
  assign tmp20042 = s4 ? tmp19957 : tmp20043;
  assign tmp20041 = s5 ? tmp20042 : tmp19962;
  assign tmp20040 = s6 ? tmp19949 : tmp20041;
  assign tmp20044 = ~(s6 ? tmp20018 : tmp20021);
  assign tmp20039 = s7 ? tmp20040 : tmp20044;
  assign tmp20045 = s7 ? tmp19977 : tmp20035;
  assign tmp20038 = s8 ? tmp20039 : tmp20045;
  assign tmp20032 = s9 ? tmp20033 : tmp20038;
  assign tmp19909 = s10 ? tmp19910 : tmp20032;
  assign tmp20049 = s7 ? tmp19948 : tmp20044;
  assign tmp20048 = s8 ? tmp20049 : tmp20045;
  assign tmp20047 = s9 ? tmp20033 : tmp20048;
  assign tmp20046 = s10 ? tmp19910 : tmp20047;
  assign tmp19908 = s11 ? tmp19909 : tmp20046;
  assign tmp19863 = s12 ? tmp19864 : tmp19908;
  assign tmp20058 = s3 ? tmp19916 : tmp19894;
  assign tmp20062 = s0 ? tmp19635 : tmp19720;
  assign tmp20061 = s1 ? tmp20062 : tmp19635;
  assign tmp20063 = s1 ? tmp19896 : tmp19789;
  assign tmp20060 = s2 ? tmp20061 : tmp20063;
  assign tmp20059 = s3 ? tmp20060 : tmp19953;
  assign tmp20057 = s4 ? tmp20058 : tmp20059;
  assign tmp20068 = s1 ? tmp19896 : tmp19637;
  assign tmp20069 = s1 ? tmp19637 : tmp19896;
  assign tmp20067 = s2 ? tmp20068 : tmp20069;
  assign tmp20073 = l1 ? tmp19635 : 0;
  assign tmp20072 = s0 ? tmp19635 : tmp20073;
  assign tmp20071 = s1 ? 1 : tmp20072;
  assign tmp20070 = s2 ? tmp19637 : tmp20071;
  assign tmp20066 = s3 ? tmp20067 : tmp20070;
  assign tmp20076 = s1 ? tmp19637 : tmp19806;
  assign tmp20078 = ~(s0 ? tmp19635 : tmp19720);
  assign tmp20077 = ~(s1 ? tmp19622 : tmp20078);
  assign tmp20075 = s2 ? tmp20076 : tmp20077;
  assign tmp20081 = ~(s0 ? 1 : tmp19612);
  assign tmp20080 = s1 ? tmp20072 : tmp20081;
  assign tmp20079 = s2 ? tmp20080 : 1;
  assign tmp20074 = s3 ? tmp20075 : tmp20079;
  assign tmp20065 = s4 ? tmp20066 : tmp20074;
  assign tmp20085 = s0 ? tmp20073 : tmp19635;
  assign tmp20084 = s2 ? tmp19938 : tmp20085;
  assign tmp20086 = s2 ? tmp19938 : tmp19946;
  assign tmp20083 = s3 ? tmp20084 : tmp20086;
  assign tmp20089 = s1 ? tmp19637 : tmp20072;
  assign tmp20088 = s2 ? tmp19635 : tmp20089;
  assign tmp20087 = s3 ? tmp20088 : tmp19945;
  assign tmp20082 = s4 ? tmp20083 : tmp20087;
  assign tmp20064 = s5 ? tmp20065 : tmp20082;
  assign tmp20056 = s6 ? tmp20057 : tmp20064;
  assign tmp20094 = s1 ? tmp19896 : tmp19720;
  assign tmp20093 = s2 ? tmp20061 : tmp20094;
  assign tmp20092 = s3 ? tmp20093 : tmp19953;
  assign tmp20091 = s4 ? tmp20058 : tmp20092;
  assign tmp20099 = s1 ? tmp19635 : tmp19896;
  assign tmp20098 = s2 ? tmp19895 : tmp20099;
  assign tmp20100 = s2 ? tmp19635 : tmp20071;
  assign tmp20097 = s3 ? tmp20098 : tmp20100;
  assign tmp20102 = s2 ? tmp20076 : tmp19635;
  assign tmp20104 = s1 ? tmp20072 : tmp19635;
  assign tmp20103 = s2 ? tmp20104 : 1;
  assign tmp20101 = s3 ? tmp20102 : tmp20103;
  assign tmp20096 = s4 ? tmp20097 : tmp20101;
  assign tmp20108 = s1 ? tmp19635 : tmp20085;
  assign tmp20107 = s2 ? tmp19938 : tmp20108;
  assign tmp20111 = s0 ? tmp20073 : 1;
  assign tmp20110 = s1 ? tmp20111 : 1;
  assign tmp20109 = s2 ? tmp20110 : tmp19888;
  assign tmp20106 = s3 ? tmp20107 : tmp20109;
  assign tmp20114 = s1 ? tmp19635 : tmp20072;
  assign tmp20113 = s2 ? 1 : tmp20114;
  assign tmp20112 = s3 ? tmp20113 : tmp19635;
  assign tmp20105 = s4 ? tmp20106 : tmp20112;
  assign tmp20095 = s5 ? tmp20096 : tmp20105;
  assign tmp20090 = s6 ? tmp20091 : tmp20095;
  assign tmp20055 = s7 ? tmp20056 : tmp20090;
  assign tmp20120 = l1 ? tmp19635 : 1;
  assign tmp20122 = ~(l1 ? tmp19635 : 1);
  assign tmp20121 = ~(s0 ? tmp19614 : tmp20122);
  assign tmp20119 = s1 ? tmp20120 : tmp20121;
  assign tmp20125 = s0 ? tmp20120 : 1;
  assign tmp20124 = s1 ? tmp20125 : tmp20120;
  assign tmp20123 = s2 ? tmp20120 : tmp20124;
  assign tmp20118 = s3 ? tmp20119 : tmp20123;
  assign tmp20129 = s0 ? tmp20120 : tmp19720;
  assign tmp20128 = s1 ? tmp20129 : tmp20120;
  assign tmp20130 = s1 ? tmp20125 : tmp19789;
  assign tmp20127 = s2 ? tmp20128 : tmp20130;
  assign tmp20133 = s0 ? 1 : tmp20120;
  assign tmp20132 = ~(s1 ? tmp20120 : tmp20133);
  assign tmp20131 = ~(s2 ? tmp19954 : tmp20132);
  assign tmp20126 = s3 ? tmp20127 : tmp20131;
  assign tmp20117 = s4 ? tmp20118 : tmp20126;
  assign tmp20138 = s1 ? tmp20125 : tmp20133;
  assign tmp20139 = s1 ? tmp20133 : tmp20125;
  assign tmp20137 = s2 ? tmp20138 : tmp20139;
  assign tmp20141 = s1 ? 1 : tmp20120;
  assign tmp20140 = s2 ? tmp20133 : tmp20141;
  assign tmp20136 = s3 ? tmp20137 : tmp20140;
  assign tmp20144 = s1 ? tmp20133 : tmp19720;
  assign tmp20146 = ~(s0 ? tmp20120 : tmp19720);
  assign tmp20145 = ~(s1 ? tmp19614 : tmp20146);
  assign tmp20143 = s2 ? tmp20144 : tmp20145;
  assign tmp20148 = s1 ? tmp20120 : tmp19917;
  assign tmp20147 = s2 ? tmp20148 : 1;
  assign tmp20142 = s3 ? tmp20143 : tmp20147;
  assign tmp20135 = s4 ? tmp20136 : tmp20142;
  assign tmp20152 = s1 ? tmp20125 : 1;
  assign tmp20154 = s0 ? tmp19635 : tmp20120;
  assign tmp20153 = s1 ? tmp20133 : tmp20154;
  assign tmp20151 = s2 ? tmp20152 : tmp20153;
  assign tmp20150 = s3 ? tmp20151 : tmp20086;
  assign tmp20158 = s0 ? tmp20120 : tmp19635;
  assign tmp20157 = s1 ? tmp20133 : tmp20158;
  assign tmp20156 = s2 ? tmp19846 : tmp20157;
  assign tmp20155 = s3 ? tmp20156 : tmp19945;
  assign tmp20149 = s4 ? tmp20150 : tmp20155;
  assign tmp20134 = s5 ? tmp20135 : tmp20149;
  assign tmp20116 = s6 ? tmp20117 : tmp20134;
  assign tmp20163 = s1 ? tmp20125 : tmp19720;
  assign tmp20162 = s2 ? tmp20128 : tmp20163;
  assign tmp20161 = s3 ? tmp20162 : tmp20131;
  assign tmp20160 = s4 ? tmp20118 : tmp20161;
  assign tmp20168 = s1 ? tmp20120 : tmp20125;
  assign tmp20167 = s2 ? tmp20124 : tmp20168;
  assign tmp20169 = s2 ? tmp20120 : tmp20141;
  assign tmp20166 = s3 ? tmp20167 : tmp20169;
  assign tmp20171 = s2 ? tmp20144 : tmp20120;
  assign tmp20173 = s1 ? tmp20120 : tmp19635;
  assign tmp20172 = s2 ? tmp20173 : 1;
  assign tmp20170 = s3 ? tmp20171 : tmp20172;
  assign tmp20165 = s4 ? tmp20166 : tmp20170;
  assign tmp20176 = s2 ? tmp20152 : tmp20173;
  assign tmp20175 = s3 ? tmp20176 : tmp20109;
  assign tmp20179 = s1 ? tmp20120 : tmp20073;
  assign tmp20178 = s2 ? 1 : tmp20179;
  assign tmp20177 = s3 ? tmp20178 : tmp19635;
  assign tmp20174 = s4 ? tmp20175 : tmp20177;
  assign tmp20164 = s5 ? tmp20165 : tmp20174;
  assign tmp20159 = s6 ? tmp20160 : tmp20164;
  assign tmp20115 = s7 ? tmp20116 : tmp20159;
  assign tmp20054 = s8 ? tmp20055 : tmp20115;
  assign tmp20187 = s1 ? 1 : tmp20158;
  assign tmp20186 = s2 ? tmp20133 : tmp20187;
  assign tmp20185 = s3 ? tmp20137 : tmp20186;
  assign tmp20190 = s1 ? tmp20133 : tmp19806;
  assign tmp20191 = ~(s1 ? tmp19622 : tmp20146);
  assign tmp20189 = s2 ? tmp20190 : tmp20191;
  assign tmp20193 = s1 ? tmp20158 : tmp20081;
  assign tmp20192 = s2 ? tmp20193 : 1;
  assign tmp20188 = s3 ? tmp20189 : tmp20192;
  assign tmp20184 = s4 ? tmp20185 : tmp20188;
  assign tmp20196 = s2 ? tmp20152 : tmp20154;
  assign tmp20195 = s3 ? tmp20196 : tmp20086;
  assign tmp20198 = s2 ? tmp19635 : tmp20157;
  assign tmp20197 = s3 ? tmp20198 : tmp19945;
  assign tmp20194 = s4 ? tmp20195 : tmp20197;
  assign tmp20183 = s5 ? tmp20184 : tmp20194;
  assign tmp20182 = s6 ? tmp20117 : tmp20183;
  assign tmp20203 = s2 ? tmp20120 : tmp20187;
  assign tmp20202 = s3 ? tmp20167 : tmp20203;
  assign tmp20205 = s2 ? tmp20190 : tmp20120;
  assign tmp20207 = s1 ? tmp20158 : tmp19635;
  assign tmp20206 = s2 ? tmp20207 : 1;
  assign tmp20204 = s3 ? tmp20205 : tmp20206;
  assign tmp20201 = s4 ? tmp20202 : tmp20204;
  assign tmp20210 = s2 ? tmp19938 : tmp19888;
  assign tmp20209 = s3 ? tmp20176 : tmp20210;
  assign tmp20212 = s2 ? 1 : tmp20173;
  assign tmp20211 = s3 ? tmp20212 : tmp19635;
  assign tmp20208 = s4 ? tmp20209 : tmp20211;
  assign tmp20200 = s5 ? tmp20201 : tmp20208;
  assign tmp20199 = s6 ? tmp20160 : tmp20200;
  assign tmp20181 = s7 ? tmp20182 : tmp20199;
  assign tmp20180 = s8 ? tmp20115 : tmp20181;
  assign tmp20053 = s9 ? tmp20054 : tmp20180;
  assign tmp20220 = s2 ? tmp19938 : tmp19635;
  assign tmp20219 = s3 ? tmp20220 : tmp20109;
  assign tmp20223 = s1 ? tmp19635 : tmp20073;
  assign tmp20222 = s2 ? 1 : tmp20223;
  assign tmp20221 = s3 ? tmp20222 : tmp19635;
  assign tmp20218 = s4 ? tmp20219 : tmp20221;
  assign tmp20217 = s5 ? tmp20096 : tmp20218;
  assign tmp20216 = s6 ? tmp20091 : tmp20217;
  assign tmp20215 = s7 ? tmp20056 : tmp20216;
  assign tmp20214 = s8 ? tmp20215 : tmp20056;
  assign tmp20229 = s3 ? tmp19967 : tmp19635;
  assign tmp20228 = s4 ? tmp20106 : tmp20229;
  assign tmp20227 = s5 ? tmp20096 : tmp20228;
  assign tmp20226 = s6 ? tmp20091 : tmp20227;
  assign tmp20234 = s2 ? 1 : tmp20120;
  assign tmp20233 = s3 ? tmp20234 : tmp19635;
  assign tmp20232 = s4 ? tmp20209 : tmp20233;
  assign tmp20231 = s5 ? tmp20201 : tmp20232;
  assign tmp20230 = s6 ? tmp20160 : tmp20231;
  assign tmp20225 = s7 ? tmp20226 : tmp20230;
  assign tmp20238 = s4 ? tmp20175 : tmp20233;
  assign tmp20237 = s5 ? tmp20165 : tmp20238;
  assign tmp20236 = s6 ? tmp20160 : tmp20237;
  assign tmp20241 = s4 ? tmp20219 : tmp20229;
  assign tmp20240 = s5 ? tmp20096 : tmp20241;
  assign tmp20239 = s6 ? tmp20091 : tmp20240;
  assign tmp20235 = s7 ? tmp20236 : tmp20239;
  assign tmp20224 = s8 ? tmp20225 : tmp20235;
  assign tmp20213 = s9 ? tmp20214 : tmp20224;
  assign tmp20052 = s10 ? tmp20053 : tmp20213;
  assign tmp20245 = s7 ? tmp20090 : tmp20199;
  assign tmp20246 = s7 ? tmp20159 : tmp20216;
  assign tmp20244 = s8 ? tmp20245 : tmp20246;
  assign tmp20243 = s9 ? tmp20214 : tmp20244;
  assign tmp20242 = s10 ? tmp20053 : tmp20243;
  assign tmp20051 = s11 ? tmp20052 : tmp20242;
  assign tmp20255 = ~(s2 ? tmp19635 : tmp19919);
  assign tmp20254 = s3 ? tmp19651 : tmp20255;
  assign tmp20257 = s2 ? tmp19919 : tmp19648;
  assign tmp20259 = s1 ? 1 : tmp19780;
  assign tmp20258 = ~(s2 ? tmp20259 : tmp19612);
  assign tmp20256 = ~(s3 ? tmp20257 : tmp20258);
  assign tmp20253 = s4 ? tmp20254 : tmp20256;
  assign tmp20264 = s1 ? tmp19649 : tmp20081;
  assign tmp20263 = s2 ? tmp20264 : tmp19974;
  assign tmp20262 = s3 ? tmp20263 : tmp19975;
  assign tmp20267 = ~(s1 ? 1 : tmp19933);
  assign tmp20266 = s2 ? tmp19944 : tmp20267;
  assign tmp20269 = s1 ? tmp19635 : tmp20081;
  assign tmp20268 = s2 ? tmp20269 : 1;
  assign tmp20265 = s3 ? tmp20266 : tmp20268;
  assign tmp20261 = s4 ? tmp20262 : tmp20265;
  assign tmp20271 = s3 ? tmp20220 : tmp20086;
  assign tmp20274 = s1 ? tmp19637 : tmp19635;
  assign tmp20273 = s2 ? tmp19635 : tmp20274;
  assign tmp20272 = s3 ? tmp20273 : tmp19945;
  assign tmp20270 = s4 ? tmp20271 : tmp20272;
  assign tmp20260 = ~(s5 ? tmp20261 : tmp20270);
  assign tmp20252 = s6 ? tmp20253 : tmp20260;
  assign tmp20279 = s1 ? 1 : 0;
  assign tmp20278 = ~(s2 ? tmp20279 : tmp19612);
  assign tmp20277 = ~(s3 ? tmp20257 : tmp20278);
  assign tmp20276 = s4 ? tmp20254 : tmp20277;
  assign tmp20283 = s2 ? tmp19919 : tmp19982;
  assign tmp20282 = s3 ? tmp20283 : tmp19887;
  assign tmp20285 = s2 ? tmp19944 : tmp19635;
  assign tmp20284 = s3 ? tmp20285 : tmp19879;
  assign tmp20281 = s4 ? tmp20282 : tmp20284;
  assign tmp20287 = s3 ? tmp20073 : tmp19635;
  assign tmp20286 = s4 ? tmp20219 : tmp20287;
  assign tmp20280 = ~(s5 ? tmp20281 : tmp20286);
  assign tmp20275 = s6 ? tmp20276 : tmp20280;
  assign tmp20251 = s7 ? tmp20252 : tmp20275;
  assign tmp20294 = s0 ? tmp20120 : 0;
  assign tmp20293 = s1 ? tmp20294 : tmp20120;
  assign tmp20295 = s1 ? tmp20294 : tmp19806;
  assign tmp20292 = s2 ? tmp20293 : tmp20295;
  assign tmp20296 = ~(s2 ? tmp19924 : tmp20122);
  assign tmp20291 = s3 ? tmp20292 : tmp20296;
  assign tmp20290 = s4 ? tmp20118 : tmp20291;
  assign tmp20302 = ~(s0 ? 1 : tmp20122);
  assign tmp20301 = s1 ? tmp20294 : tmp20302;
  assign tmp20304 = s0 ? 1 : tmp20122;
  assign tmp20305 = ~(s0 ? tmp20120 : 1);
  assign tmp20303 = ~(s1 ? tmp20304 : tmp20305);
  assign tmp20300 = s2 ? tmp20301 : tmp20303;
  assign tmp20299 = s3 ? tmp20300 : tmp20140;
  assign tmp20309 = ~(s0 ? 1 : tmp19614);
  assign tmp20308 = s1 ? tmp20133 : tmp20309;
  assign tmp20311 = ~(s0 ? tmp20120 : 0);
  assign tmp20310 = ~(s1 ? tmp19711 : tmp20311);
  assign tmp20307 = s2 ? tmp20308 : tmp20310;
  assign tmp20306 = s3 ? tmp20307 : tmp20147;
  assign tmp20298 = s4 ? tmp20299 : tmp20306;
  assign tmp20315 = s1 ? tmp20120 : tmp20154;
  assign tmp20314 = s2 ? tmp20152 : tmp20315;
  assign tmp20313 = s3 ? tmp20314 : tmp20086;
  assign tmp20312 = s4 ? tmp20313 : tmp20155;
  assign tmp20297 = s5 ? tmp20298 : tmp20312;
  assign tmp20289 = s6 ? tmp20290 : tmp20297;
  assign tmp20320 = s1 ? tmp20294 : tmp19720;
  assign tmp20319 = s2 ? tmp20293 : tmp20320;
  assign tmp20321 = ~(s2 ? tmp19954 : tmp20122);
  assign tmp20318 = s3 ? tmp20319 : tmp20321;
  assign tmp20317 = s4 ? tmp20118 : tmp20318;
  assign tmp20325 = s2 ? tmp20293 : tmp20168;
  assign tmp20324 = s3 ? tmp20325 : tmp20169;
  assign tmp20327 = s2 ? tmp20308 : tmp20120;
  assign tmp20326 = s3 ? tmp20327 : tmp20172;
  assign tmp20323 = s4 ? tmp20324 : tmp20326;
  assign tmp20322 = s5 ? tmp20323 : tmp20174;
  assign tmp20316 = s6 ? tmp20317 : tmp20322;
  assign tmp20288 = ~(s7 ? tmp20289 : tmp20316);
  assign tmp20250 = s8 ? tmp20251 : tmp20288;
  assign tmp20329 = s7 ? tmp20289 : tmp20316;
  assign tmp20335 = s2 ? tmp20264 : tmp19650;
  assign tmp20334 = s3 ? tmp20335 : tmp19887;
  assign tmp20333 = s4 ? tmp20334 : tmp20265;
  assign tmp20332 = ~(s5 ? tmp20333 : tmp20270);
  assign tmp20331 = s6 ? tmp20253 : tmp20332;
  assign tmp20340 = s2 ? tmp19919 : tmp19635;
  assign tmp20339 = s3 ? tmp20340 : tmp19887;
  assign tmp20338 = s4 ? tmp20339 : tmp20284;
  assign tmp20342 = s3 ? tmp20220 : tmp20210;
  assign tmp20341 = s4 ? tmp20342 : tmp19635;
  assign tmp20337 = ~(s5 ? tmp20338 : tmp20341);
  assign tmp20336 = s6 ? tmp20276 : tmp20337;
  assign tmp20330 = ~(s7 ? tmp20331 : tmp20336);
  assign tmp20328 = ~(s8 ? tmp20329 : tmp20330);
  assign tmp20249 = s9 ? tmp20250 : tmp20328;
  assign tmp20347 = ~(s5 ? tmp20338 : tmp20286);
  assign tmp20346 = s6 ? tmp20276 : tmp20347;
  assign tmp20345 = s7 ? tmp20331 : tmp20346;
  assign tmp20344 = s8 ? tmp20345 : tmp20331;
  assign tmp20350 = ~(s5 ? tmp20281 : tmp20241);
  assign tmp20349 = s6 ? tmp20276 : tmp20350;
  assign tmp20353 = s5 ? tmp20323 : tmp20238;
  assign tmp20352 = s6 ? tmp20317 : tmp20353;
  assign tmp20355 = ~(s5 ? tmp20338 : tmp20241);
  assign tmp20354 = ~(s6 ? tmp20276 : tmp20355);
  assign tmp20351 = ~(s7 ? tmp20352 : tmp20354);
  assign tmp20348 = s8 ? tmp20349 : tmp20351;
  assign tmp20343 = s9 ? tmp20344 : tmp20348;
  assign tmp20248 = s10 ? tmp20249 : tmp20343;
  assign tmp20360 = ~(s6 ? tmp20276 : tmp20347);
  assign tmp20359 = ~(s7 ? tmp20316 : tmp20360);
  assign tmp20358 = s8 ? tmp20275 : tmp20359;
  assign tmp20357 = s9 ? tmp20344 : tmp20358;
  assign tmp20356 = s10 ? tmp20249 : tmp20357;
  assign tmp20247 = ~(s11 ? tmp20248 : tmp20356);
  assign tmp20050 = s12 ? tmp20051 : tmp20247;
  assign tmp19862 = ~(s13 ? tmp19863 : tmp20050);
  assign tmp19600 = s14 ? tmp19601 : tmp19862;
  assign tmp20371 = s1 ? 1 : tmp20122;
  assign tmp20370 = ~(s2 ? tmp20304 : tmp20371);
  assign tmp20369 = s3 ? tmp19644 : tmp20370;
  assign tmp20374 = ~(s1 ? tmp19649 : 0);
  assign tmp20373 = s2 ? tmp20371 : tmp20374;
  assign tmp20376 = s1 ? 1 : tmp20304;
  assign tmp20375 = s2 ? tmp20376 : tmp20122;
  assign tmp20372 = ~(s3 ? tmp20373 : tmp20375);
  assign tmp20368 = s4 ? tmp20369 : tmp20372;
  assign tmp20381 = s1 ? 1 : tmp20311;
  assign tmp20380 = s2 ? 1 : tmp20381;
  assign tmp20379 = s3 ? tmp20380 : tmp20375;
  assign tmp20384 = s1 ? tmp20120 : 0;
  assign tmp20383 = s2 ? tmp20384 : 0;
  assign tmp20386 = s1 ? tmp19651 : tmp20304;
  assign tmp20385 = ~(s2 ? tmp20386 : tmp20122);
  assign tmp20382 = ~(s3 ? tmp20383 : tmp20385);
  assign tmp20378 = s4 ? tmp20379 : tmp20382;
  assign tmp20390 = s1 ? tmp20120 : tmp20294;
  assign tmp20389 = s2 ? tmp20390 : 0;
  assign tmp20392 = s1 ? 1 : tmp19711;
  assign tmp20393 = s1 ? tmp19687 : tmp19933;
  assign tmp20391 = ~(s2 ? tmp20392 : tmp20393);
  assign tmp20388 = s3 ? tmp20389 : tmp20391;
  assign tmp20396 = ~(s1 ? tmp20294 : 0);
  assign tmp20395 = s2 ? tmp20376 : tmp20396;
  assign tmp20398 = s1 ? tmp19614 : tmp19687;
  assign tmp20397 = s2 ? tmp20398 : tmp20374;
  assign tmp20394 = ~(s3 ? tmp20395 : tmp20397);
  assign tmp20387 = ~(s4 ? tmp20388 : tmp20394);
  assign tmp20377 = ~(s5 ? tmp20378 : tmp20387);
  assign tmp20367 = s6 ? tmp20368 : tmp20377;
  assign tmp20402 = s2 ? tmp20371 : tmp20122;
  assign tmp20401 = ~(s3 ? tmp20373 : tmp20402);
  assign tmp20400 = s4 ? tmp20369 : tmp20401;
  assign tmp20405 = s3 ? tmp20380 : tmp20402;
  assign tmp20408 = s1 ? tmp19651 : tmp20122;
  assign tmp20407 = ~(s2 ? tmp20408 : tmp20122);
  assign tmp20406 = ~(s3 ? tmp20383 : tmp20407);
  assign tmp20404 = s4 ? tmp20405 : tmp20406;
  assign tmp20412 = s1 ? 1 : tmp19614;
  assign tmp20413 = ~(s1 ? tmp19635 : 0);
  assign tmp20411 = ~(s2 ? tmp20412 : tmp20413);
  assign tmp20410 = s3 ? tmp20389 : tmp20411;
  assign tmp20415 = s2 ? tmp20371 : tmp20311;
  assign tmp20414 = ~(s3 ? tmp20415 : tmp19844);
  assign tmp20409 = ~(s4 ? tmp20410 : tmp20414);
  assign tmp20403 = ~(s5 ? tmp20404 : tmp20409);
  assign tmp20399 = s6 ? tmp20400 : tmp20403;
  assign tmp20366 = s7 ? tmp20367 : tmp20399;
  assign tmp20417 = s8 ? tmp20366 : tmp20367;
  assign tmp20422 = s2 ? tmp20371 : 1;
  assign tmp20421 = ~(s3 ? tmp20422 : tmp19844);
  assign tmp20420 = ~(s4 ? tmp20410 : tmp20421);
  assign tmp20419 = ~(s5 ? tmp20404 : tmp20420);
  assign tmp20418 = s6 ? tmp20400 : tmp20419;
  assign tmp20416 = s9 ? tmp20417 : tmp20418;
  assign tmp20365 = s10 ? tmp20366 : tmp20416;
  assign tmp20424 = s9 ? tmp20417 : tmp20399;
  assign tmp20423 = s10 ? tmp20366 : tmp20424;
  assign tmp20364 = s11 ? tmp20365 : tmp20423;
  assign tmp20432 = l1 ? 1 : tmp19635;
  assign tmp20431 = s0 ? tmp19614 : tmp20432;
  assign tmp20434 = s0 ? tmp20432 : tmp19614;
  assign tmp20433 = s1 ? tmp19614 : tmp20434;
  assign tmp20430 = s2 ? tmp20431 : tmp20433;
  assign tmp20429 = s3 ? tmp19954 : tmp20430;
  assign tmp20437 = s1 ? tmp19614 : tmp20431;
  assign tmp20436 = s2 ? tmp20437 : tmp19614;
  assign tmp20438 = s2 ? tmp20437 : tmp20432;
  assign tmp20435 = s3 ? tmp20436 : tmp20438;
  assign tmp20428 = s4 ? tmp20429 : tmp20435;
  assign tmp20444 = ~(s0 ? tmp20432 : 1);
  assign tmp20443 = s1 ? 1 : tmp20444;
  assign tmp20442 = s2 ? 1 : tmp20443;
  assign tmp20447 = s0 ? 1 : tmp20432;
  assign tmp20446 = s1 ? tmp19614 : tmp20447;
  assign tmp20445 = ~(s2 ? tmp20446 : tmp20432);
  assign tmp20441 = s3 ? tmp20442 : tmp20445;
  assign tmp20450 = s1 ? tmp20434 : tmp19614;
  assign tmp20449 = s2 ? tmp20450 : tmp19614;
  assign tmp20448 = ~(s3 ? tmp20449 : tmp20438);
  assign tmp20440 = s4 ? tmp20441 : tmp20448;
  assign tmp20454 = s1 ? tmp20432 : tmp19711;
  assign tmp20453 = s2 ? tmp20454 : tmp19614;
  assign tmp20456 = s1 ? 1 : tmp19651;
  assign tmp20458 = s0 ? tmp19635 : tmp19614;
  assign tmp20457 = ~(s1 ? tmp20458 : tmp19614);
  assign tmp20455 = ~(s2 ? tmp20456 : tmp20457);
  assign tmp20452 = s3 ? tmp20453 : tmp20455;
  assign tmp20463 = ~(l1 ? 1 : tmp19635);
  assign tmp20462 = s0 ? 1 : tmp20463;
  assign tmp20461 = s1 ? 1 : tmp20462;
  assign tmp20460 = s2 ? tmp20461 : tmp20008;
  assign tmp20466 = ~(s0 ? tmp19635 : tmp19614);
  assign tmp20465 = s1 ? tmp19651 : tmp20466;
  assign tmp20467 = ~(s1 ? tmp19717 : 0);
  assign tmp20464 = s2 ? tmp20465 : tmp20467;
  assign tmp20459 = ~(s3 ? tmp20460 : tmp20464);
  assign tmp20451 = ~(s4 ? tmp20452 : tmp20459);
  assign tmp20439 = ~(s5 ? tmp20440 : tmp20451);
  assign tmp20427 = s6 ? tmp20428 : tmp20439;
  assign tmp20472 = s1 ? tmp19614 : tmp20432;
  assign tmp20471 = s2 ? tmp20472 : tmp20432;
  assign tmp20470 = s3 ? tmp20436 : tmp20471;
  assign tmp20469 = s4 ? tmp20429 : tmp20470;
  assign tmp20476 = ~(s2 ? tmp20472 : tmp20432);
  assign tmp20475 = s3 ? tmp20442 : tmp20476;
  assign tmp20477 = ~(s3 ? tmp20449 : tmp20471);
  assign tmp20474 = s4 ? tmp20475 : tmp20477;
  assign tmp20481 = s1 ? tmp20432 : tmp19614;
  assign tmp20480 = s2 ? tmp20481 : tmp19614;
  assign tmp20483 = s1 ? 1 : tmp19612;
  assign tmp20482 = ~(s2 ? tmp20483 : tmp19720);
  assign tmp20479 = s3 ? tmp20480 : tmp20482;
  assign tmp20486 = s1 ? 1 : tmp20463;
  assign tmp20485 = s2 ? tmp20486 : 1;
  assign tmp20487 = ~(s1 ? tmp19635 : tmp19614);
  assign tmp20484 = ~(s3 ? tmp20485 : tmp20487);
  assign tmp20478 = ~(s4 ? tmp20479 : tmp20484);
  assign tmp20473 = ~(s5 ? tmp20474 : tmp20478);
  assign tmp20468 = s6 ? tmp20469 : tmp20473;
  assign tmp20426 = s7 ? tmp20427 : tmp20468;
  assign tmp20489 = s8 ? tmp20426 : tmp20427;
  assign tmp20488 = s9 ? tmp20489 : tmp20468;
  assign tmp20425 = s10 ? tmp20426 : tmp20488;
  assign tmp20363 = s12 ? tmp20364 : tmp20425;
  assign tmp20499 = s1 ? tmp19635 : tmp19783;
  assign tmp20501 = s1 ? tmp19637 : tmp19917;
  assign tmp20502 = ~(s1 ? tmp19717 : tmp19612);
  assign tmp20500 = s2 ? tmp20501 : tmp20502;
  assign tmp20498 = s3 ? tmp20499 : tmp20500;
  assign tmp20504 = s2 ? tmp19895 : tmp19938;
  assign tmp20505 = s2 ? tmp19946 : tmp19635;
  assign tmp20503 = s3 ? tmp20504 : tmp20505;
  assign tmp20497 = s4 ? tmp20498 : tmp20503;
  assign tmp20509 = s2 ? tmp19818 : tmp19664;
  assign tmp20511 = s1 ? tmp19719 : tmp19637;
  assign tmp20510 = ~(s2 ? tmp20511 : tmp20104);
  assign tmp20508 = s3 ? tmp20509 : tmp20510;
  assign tmp20514 = s1 ? 1 : tmp19896;
  assign tmp20513 = s2 ? tmp19846 : tmp20514;
  assign tmp20516 = s1 ? tmp19614 : tmp20458;
  assign tmp20515 = s2 ? tmp19635 : tmp20516;
  assign tmp20512 = ~(s3 ? tmp20513 : tmp20515);
  assign tmp20507 = s4 ? tmp20508 : tmp20512;
  assign tmp20520 = s1 ? tmp19635 : tmp20062;
  assign tmp20519 = s2 ? tmp20520 : tmp20467;
  assign tmp20521 = ~(s2 ? 1 : tmp19654);
  assign tmp20518 = s3 ? tmp20519 : tmp20521;
  assign tmp20525 = s0 ? tmp19635 : tmp19783;
  assign tmp20524 = s1 ? tmp20525 : 1;
  assign tmp20523 = s2 ? tmp20264 : tmp20524;
  assign tmp20527 = s1 ? tmp19622 : tmp19651;
  assign tmp20526 = ~(s2 ? tmp20527 : tmp20413);
  assign tmp20522 = s3 ? tmp20523 : tmp20526;
  assign tmp20517 = ~(s4 ? tmp20518 : tmp20522);
  assign tmp20506 = ~(s5 ? tmp20507 : tmp20517);
  assign tmp20496 = s6 ? tmp20497 : tmp20506;
  assign tmp20531 = s2 ? tmp19888 : tmp19635;
  assign tmp20530 = s3 ? tmp20504 : tmp20531;
  assign tmp20529 = s4 ? tmp20498 : tmp20530;
  assign tmp20536 = ~(s1 ? tmp20072 : tmp19635);
  assign tmp20535 = s2 ? tmp19844 : tmp20536;
  assign tmp20534 = s3 ? tmp20509 : tmp20535;
  assign tmp20538 = s2 ? tmp19846 : tmp19635;
  assign tmp20540 = s1 ? tmp19614 : tmp19635;
  assign tmp20539 = s2 ? tmp19635 : tmp20540;
  assign tmp20537 = ~(s3 ? tmp20538 : tmp20539);
  assign tmp20533 = s4 ? tmp20534 : tmp20537;
  assign tmp20544 = s1 ? tmp19635 : tmp19720;
  assign tmp20543 = s2 ? tmp20544 : 1;
  assign tmp20545 = ~(s2 ? 1 : tmp19612);
  assign tmp20542 = s3 ? tmp20543 : tmp20545;
  assign tmp20547 = s2 ? tmp20483 : tmp19611;
  assign tmp20548 = s2 ? tmp20483 : tmp19612;
  assign tmp20546 = ~(s3 ? tmp20547 : tmp20548);
  assign tmp20541 = ~(s4 ? tmp20542 : tmp20546);
  assign tmp20532 = ~(s5 ? tmp20533 : tmp20541);
  assign tmp20528 = s6 ? tmp20529 : tmp20532;
  assign tmp20495 = s7 ? tmp20496 : tmp20528;
  assign tmp20553 = s2 ? tmp19635 : tmp19938;
  assign tmp20552 = s3 ? tmp20553 : tmp20505;
  assign tmp20551 = s4 ? tmp20498 : tmp20552;
  assign tmp20557 = s2 ? tmp19846 : tmp19888;
  assign tmp20556 = ~(s3 ? tmp20557 : tmp20515);
  assign tmp20555 = s4 ? tmp20508 : tmp20556;
  assign tmp20554 = ~(s5 ? tmp20555 : tmp20517);
  assign tmp20550 = s6 ? tmp20551 : tmp20554;
  assign tmp20560 = s3 ? tmp20553 : tmp20531;
  assign tmp20559 = s4 ? tmp20498 : tmp20560;
  assign tmp20558 = s6 ? tmp20559 : tmp20532;
  assign tmp20549 = s7 ? tmp20550 : tmp20558;
  assign tmp20494 = s8 ? tmp20495 : tmp20549;
  assign tmp20567 = s2 ? tmp20520 : tmp19720;
  assign tmp20566 = s3 ? tmp20567 : tmp20521;
  assign tmp20569 = s2 ? tmp20264 : tmp20525;
  assign tmp20568 = s3 ? tmp20569 : tmp20526;
  assign tmp20565 = ~(s4 ? tmp20566 : tmp20568);
  assign tmp20564 = ~(s5 ? tmp20555 : tmp20565);
  assign tmp20563 = s6 ? tmp20551 : tmp20564;
  assign tmp20573 = s3 ? tmp20544 : tmp20545;
  assign tmp20572 = ~(s4 ? tmp20573 : tmp20546);
  assign tmp20571 = ~(s5 ? tmp20533 : tmp20572);
  assign tmp20570 = s6 ? tmp20559 : tmp20571;
  assign tmp20562 = s7 ? tmp20563 : tmp20570;
  assign tmp20561 = s8 ? tmp20549 : tmp20562;
  assign tmp20493 = s9 ? tmp20494 : tmp20561;
  assign tmp20575 = s8 ? tmp20562 : tmp20563;
  assign tmp20581 = ~(s3 ? tmp20547 : tmp20483);
  assign tmp20580 = ~(s4 ? tmp20542 : tmp20581);
  assign tmp20579 = ~(s5 ? tmp20533 : tmp20580);
  assign tmp20578 = s6 ? tmp20529 : tmp20579;
  assign tmp20584 = ~(s4 ? tmp20573 : tmp20581);
  assign tmp20583 = ~(s5 ? tmp20533 : tmp20584);
  assign tmp20582 = s6 ? tmp20559 : tmp20583;
  assign tmp20577 = s7 ? tmp20578 : tmp20582;
  assign tmp20586 = s6 ? tmp20559 : tmp20579;
  assign tmp20585 = s7 ? tmp20586 : tmp20582;
  assign tmp20576 = s8 ? tmp20577 : tmp20585;
  assign tmp20574 = s9 ? tmp20575 : tmp20576;
  assign tmp20492 = s10 ? tmp20493 : tmp20574;
  assign tmp20590 = s7 ? tmp20528 : tmp20570;
  assign tmp20591 = s7 ? tmp20558 : tmp20570;
  assign tmp20589 = s8 ? tmp20590 : tmp20591;
  assign tmp20588 = s9 ? tmp20575 : tmp20589;
  assign tmp20587 = s10 ? tmp20493 : tmp20588;
  assign tmp20491 = s11 ? tmp20492 : tmp20587;
  assign tmp20598 = s2 ? tmp19627 : tmp19688;
  assign tmp20597 = s3 ? 1 : tmp20598;
  assign tmp20601 = s1 ? 1 : tmp19627;
  assign tmp20600 = s2 ? tmp20601 : 1;
  assign tmp20602 = s2 ? tmp20601 : tmp19611;
  assign tmp20599 = s3 ? tmp20600 : tmp20602;
  assign tmp20596 = s4 ? tmp20597 : tmp20599;
  assign tmp20606 = s2 ? 1 : tmp19688;
  assign tmp20605 = s3 ? tmp20606 : tmp20602;
  assign tmp20609 = s1 ? tmp19621 : 1;
  assign tmp20608 = s2 ? tmp20609 : 1;
  assign tmp20607 = s3 ? tmp20608 : tmp20602;
  assign tmp20604 = s4 ? tmp20605 : tmp20607;
  assign tmp20613 = s1 ? tmp19611 : tmp19622;
  assign tmp20612 = s2 ? tmp20613 : 1;
  assign tmp20614 = s2 ? tmp20601 : tmp20609;
  assign tmp20611 = s3 ? tmp20612 : tmp20614;
  assign tmp20616 = s2 ? tmp20601 : tmp19730;
  assign tmp20618 = s1 ? tmp19627 : tmp19621;
  assign tmp20617 = s2 ? tmp20618 : 1;
  assign tmp20615 = s3 ? tmp20616 : tmp20617;
  assign tmp20610 = s4 ? tmp20611 : tmp20615;
  assign tmp20603 = s5 ? tmp20604 : tmp20610;
  assign tmp20595 = s6 ? tmp20596 : tmp20603;
  assign tmp20623 = s1 ? 1 : tmp19611;
  assign tmp20622 = s2 ? tmp20623 : tmp19611;
  assign tmp20621 = s3 ? tmp20600 : tmp20622;
  assign tmp20620 = s4 ? tmp20597 : tmp20621;
  assign tmp20626 = s3 ? tmp20606 : tmp20622;
  assign tmp20627 = s3 ? tmp20608 : tmp20622;
  assign tmp20625 = s4 ? tmp20626 : tmp20627;
  assign tmp20631 = s1 ? tmp19611 : 1;
  assign tmp20630 = s2 ? tmp20631 : 1;
  assign tmp20632 = s2 ? tmp20623 : tmp20609;
  assign tmp20629 = s3 ? tmp20630 : tmp20632;
  assign tmp20634 = s2 ? tmp20623 : 1;
  assign tmp20635 = s1 ? tmp19611 : tmp19621;
  assign tmp20633 = s3 ? tmp20634 : tmp20635;
  assign tmp20628 = s4 ? tmp20629 : tmp20633;
  assign tmp20624 = s5 ? tmp20625 : tmp20628;
  assign tmp20619 = s6 ? tmp20620 : tmp20624;
  assign tmp20594 = s7 ? tmp20595 : tmp20619;
  assign tmp20637 = s8 ? tmp20594 : tmp20595;
  assign tmp20641 = s3 ? tmp20634 : tmp20631;
  assign tmp20640 = s4 ? tmp20629 : tmp20641;
  assign tmp20639 = s5 ? tmp20625 : tmp20640;
  assign tmp20638 = s6 ? tmp20620 : tmp20639;
  assign tmp20636 = s9 ? tmp20637 : tmp20638;
  assign tmp20593 = s10 ? tmp20594 : tmp20636;
  assign tmp20643 = s9 ? tmp20637 : tmp20619;
  assign tmp20642 = s10 ? tmp20594 : tmp20643;
  assign tmp20592 = ~(s11 ? tmp20593 : tmp20642);
  assign tmp20490 = s12 ? tmp20491 : tmp20592;
  assign tmp20362 = s13 ? tmp20363 : tmp20490;
  assign tmp20655 = s1 ? tmp20085 : tmp19635;
  assign tmp20654 = s2 ? tmp20655 : tmp19919;
  assign tmp20653 = s3 ? tmp19916 : tmp20654;
  assign tmp20658 = s1 ? tmp19614 : tmp19651;
  assign tmp20657 = ~(s2 ? tmp20658 : tmp19612);
  assign tmp20656 = s3 ? tmp19921 : tmp20657;
  assign tmp20652 = s4 ? tmp20653 : tmp20656;
  assign tmp20663 = ~(s1 ? tmp19649 : tmp19635);
  assign tmp20662 = ~(s2 ? tmp19651 : tmp20663);
  assign tmp20661 = s3 ? tmp20263 : tmp20662;
  assign tmp20666 = s1 ? tmp19635 : tmp20309;
  assign tmp20667 = ~(s1 ? tmp19711 : tmp19933);
  assign tmp20665 = s2 ? tmp20666 : tmp20667;
  assign tmp20668 = s2 ? tmp19916 : tmp19635;
  assign tmp20664 = s3 ? tmp20665 : tmp20668;
  assign tmp20660 = s4 ? tmp20661 : tmp20664;
  assign tmp20671 = s2 ? tmp19846 : tmp20274;
  assign tmp20670 = s3 ? tmp20671 : tmp19647;
  assign tmp20675 = s0 ? tmp19614 : tmp19635;
  assign tmp20674 = s1 ? tmp20458 : tmp20675;
  assign tmp20673 = s2 ? tmp20674 : tmp19635;
  assign tmp20677 = s1 ? tmp19711 : tmp20081;
  assign tmp20678 = s1 ? tmp19635 : tmp19994;
  assign tmp20676 = s2 ? tmp20677 : tmp20678;
  assign tmp20672 = s3 ? tmp20673 : tmp20676;
  assign tmp20669 = s4 ? tmp20670 : tmp20672;
  assign tmp20659 = s5 ? tmp20660 : tmp20669;
  assign tmp20651 = s6 ? tmp20652 : tmp20659;
  assign tmp20682 = ~(s2 ? tmp19611 : tmp19612);
  assign tmp20681 = s3 ? tmp19951 : tmp20682;
  assign tmp20680 = s4 ? tmp20653 : tmp20681;
  assign tmp20685 = s3 ? tmp20283 : tmp19918;
  assign tmp20687 = s2 ? tmp20666 : tmp19961;
  assign tmp20686 = s3 ? tmp20687 : tmp20668;
  assign tmp20684 = s4 ? tmp20685 : tmp20686;
  assign tmp20692 = s0 ? tmp20073 : 0;
  assign tmp20691 = s1 ? tmp20692 : 0;
  assign tmp20690 = s2 ? tmp20691 : tmp19635;
  assign tmp20689 = s3 ? tmp20538 : tmp20690;
  assign tmp20695 = s1 ? tmp20458 : tmp19635;
  assign tmp20694 = s2 ? tmp20695 : tmp20223;
  assign tmp20696 = s2 ? tmp20540 : tmp19635;
  assign tmp20693 = s3 ? tmp20694 : tmp20696;
  assign tmp20688 = s4 ? tmp20689 : tmp20693;
  assign tmp20683 = s5 ? tmp20684 : tmp20688;
  assign tmp20679 = s6 ? tmp20680 : tmp20683;
  assign tmp20650 = s7 ? tmp20651 : tmp20679;
  assign tmp20702 = s1 ? tmp20125 : tmp19635;
  assign tmp20701 = s2 ? tmp19635 : tmp20702;
  assign tmp20700 = s3 ? tmp19916 : tmp20701;
  assign tmp20699 = s4 ? tmp20700 : tmp20656;
  assign tmp20707 = s1 ? tmp19649 : tmp20302;
  assign tmp20708 = ~(s1 ? tmp19651 : tmp19634);
  assign tmp20706 = s2 ? tmp20707 : tmp20708;
  assign tmp20711 = s0 ? tmp20432 : 0;
  assign tmp20710 = s1 ? tmp20711 : tmp19635;
  assign tmp20709 = s2 ? tmp19637 : tmp20710;
  assign tmp20705 = s3 ? tmp20706 : tmp20709;
  assign tmp20704 = s4 ? tmp20705 : tmp20664;
  assign tmp20714 = s2 ? tmp19846 : tmp20153;
  assign tmp20713 = s3 ? tmp20714 : tmp19647;
  assign tmp20717 = s1 ? tmp20458 : tmp20431;
  assign tmp20718 = s1 ? tmp19635 : tmp20158;
  assign tmp20716 = s2 ? tmp20717 : tmp20718;
  assign tmp20715 = s3 ? tmp20716 : tmp20676;
  assign tmp20712 = s4 ? tmp20713 : tmp20715;
  assign tmp20703 = s5 ? tmp20704 : tmp20712;
  assign tmp20698 = s6 ? tmp20699 : tmp20703;
  assign tmp20722 = ~(s2 ? tmp19844 : tmp19612);
  assign tmp20721 = s3 ? tmp19951 : tmp20722;
  assign tmp20720 = s4 ? tmp20700 : tmp20721;
  assign tmp20727 = s1 ? tmp19649 : tmp20120;
  assign tmp20726 = s2 ? tmp20727 : tmp20099;
  assign tmp20728 = s2 ? tmp19635 : tmp20710;
  assign tmp20725 = s3 ? tmp20726 : tmp20728;
  assign tmp20730 = s2 ? tmp20666 : tmp19635;
  assign tmp20729 = s3 ? tmp20730 : tmp19635;
  assign tmp20724 = s4 ? tmp20725 : tmp20729;
  assign tmp20733 = s2 ? tmp19846 : tmp20173;
  assign tmp20732 = s3 ? tmp20733 : tmp20690;
  assign tmp20736 = s1 ? tmp20458 : tmp20432;
  assign tmp20735 = s2 ? tmp20736 : tmp20223;
  assign tmp20734 = s3 ? tmp20735 : tmp20696;
  assign tmp20731 = s4 ? tmp20732 : tmp20734;
  assign tmp20723 = s5 ? tmp20724 : tmp20731;
  assign tmp20719 = s6 ? tmp20720 : tmp20723;
  assign tmp20697 = s7 ? tmp20698 : tmp20719;
  assign tmp20649 = s8 ? tmp20650 : tmp20697;
  assign tmp20740 = s4 ? tmp19915 : tmp20656;
  assign tmp20743 = s3 ? tmp20335 : tmp19918;
  assign tmp20742 = s4 ? tmp20743 : tmp20664;
  assign tmp20741 = s5 ? tmp20742 : tmp20669;
  assign tmp20739 = s6 ? tmp20740 : tmp20741;
  assign tmp20745 = s4 ? tmp19915 : tmp20681;
  assign tmp20748 = s3 ? tmp20340 : tmp19918;
  assign tmp20747 = s4 ? tmp20748 : tmp20729;
  assign tmp20750 = s3 ? tmp20538 : tmp19958;
  assign tmp20752 = s2 ? tmp20695 : tmp19635;
  assign tmp20751 = s3 ? tmp20752 : tmp20696;
  assign tmp20749 = s4 ? tmp20750 : tmp20751;
  assign tmp20746 = s5 ? tmp20747 : tmp20749;
  assign tmp20744 = s6 ? tmp20745 : tmp20746;
  assign tmp20738 = s7 ? tmp20739 : tmp20744;
  assign tmp20737 = s8 ? tmp20697 : tmp20738;
  assign tmp20648 = s9 ? tmp20649 : tmp20737;
  assign tmp20756 = s6 ? tmp20652 : tmp20741;
  assign tmp20758 = s5 ? tmp20747 : tmp20688;
  assign tmp20757 = s6 ? tmp20680 : tmp20758;
  assign tmp20755 = s7 ? tmp20756 : tmp20757;
  assign tmp20754 = s8 ? tmp20755 : tmp20756;
  assign tmp20764 = s3 ? tmp20687 : tmp19635;
  assign tmp20763 = s4 ? tmp20685 : tmp20764;
  assign tmp20766 = s3 ? tmp20752 : tmp20540;
  assign tmp20765 = s4 ? tmp20689 : tmp20766;
  assign tmp20762 = s5 ? tmp20763 : tmp20765;
  assign tmp20761 = s6 ? tmp20680 : tmp20762;
  assign tmp20769 = s4 ? tmp20750 : tmp20766;
  assign tmp20768 = s5 ? tmp20747 : tmp20769;
  assign tmp20767 = s6 ? tmp20745 : tmp20768;
  assign tmp20760 = s7 ? tmp20761 : tmp20767;
  assign tmp20775 = s2 ? tmp20736 : tmp19635;
  assign tmp20774 = s3 ? tmp20775 : tmp20540;
  assign tmp20773 = s4 ? tmp20732 : tmp20774;
  assign tmp20772 = s5 ? tmp20724 : tmp20773;
  assign tmp20771 = s6 ? tmp20720 : tmp20772;
  assign tmp20777 = s5 ? tmp20747 : tmp20765;
  assign tmp20776 = s6 ? tmp20680 : tmp20777;
  assign tmp20770 = s7 ? tmp20771 : tmp20776;
  assign tmp20759 = s8 ? tmp20760 : tmp20770;
  assign tmp20753 = s9 ? tmp20754 : tmp20759;
  assign tmp20647 = s10 ? tmp20648 : tmp20753;
  assign tmp20781 = s7 ? tmp20679 : tmp20744;
  assign tmp20782 = s7 ? tmp20719 : tmp20757;
  assign tmp20780 = s8 ? tmp20781 : tmp20782;
  assign tmp20779 = s9 ? tmp20754 : tmp20780;
  assign tmp20778 = s10 ? tmp20648 : tmp20779;
  assign tmp20646 = s11 ? tmp20647 : tmp20778;
  assign tmp20791 = s1 ? tmp20120 : tmp20133;
  assign tmp20793 = s1 ? tmp20133 : tmp20120;
  assign tmp20792 = s2 ? tmp20793 : tmp20124;
  assign tmp20790 = s3 ? tmp20791 : tmp20792;
  assign tmp20795 = s2 ? tmp20141 : tmp20152;
  assign tmp20796 = s2 ? tmp20015 : tmp20120;
  assign tmp20794 = s3 ? tmp20795 : tmp20796;
  assign tmp20789 = s4 ? tmp20790 : tmp20794;
  assign tmp20800 = s2 ? tmp20152 : tmp20139;
  assign tmp20801 = s2 ? tmp20133 : tmp20293;
  assign tmp20799 = s3 ? tmp20800 : tmp20801;
  assign tmp20805 = s0 ? tmp19614 : tmp20122;
  assign tmp20804 = s1 ? tmp20805 : 0;
  assign tmp20803 = s2 ? tmp20804 : 0;
  assign tmp20806 = ~(s2 ? tmp20791 : tmp19721);
  assign tmp20802 = ~(s3 ? tmp20803 : tmp20806);
  assign tmp20798 = s4 ? tmp20799 : tmp20802;
  assign tmp20809 = s2 ? tmp20301 : tmp20152;
  assign tmp20811 = ~(s1 ? tmp19614 : tmp19717);
  assign tmp20810 = s2 ? tmp19939 : tmp20811;
  assign tmp20808 = s3 ? tmp20809 : tmp20810;
  assign tmp20814 = s1 ? tmp19637 : tmp20120;
  assign tmp20815 = ~(s1 ? tmp20304 : 0);
  assign tmp20813 = s2 ? tmp20814 : tmp20815;
  assign tmp20817 = s1 ? tmp20120 : tmp20302;
  assign tmp20818 = ~(s1 ? tmp19717 : tmp19651);
  assign tmp20816 = s2 ? tmp20817 : tmp20818;
  assign tmp20812 = s3 ? tmp20813 : tmp20816;
  assign tmp20807 = s4 ? tmp20808 : tmp20812;
  assign tmp20797 = s5 ? tmp20798 : tmp20807;
  assign tmp20788 = s6 ? tmp20789 : tmp20797;
  assign tmp20822 = s2 ? tmp20029 : tmp20120;
  assign tmp20821 = s3 ? tmp20795 : tmp20822;
  assign tmp20820 = s4 ? tmp20790 : tmp20821;
  assign tmp20826 = s2 ? tmp20152 : tmp20168;
  assign tmp20827 = s2 ? tmp20120 : tmp20293;
  assign tmp20825 = s3 ? tmp20826 : tmp20827;
  assign tmp20830 = ~(s1 ? 1 : tmp19614);
  assign tmp20829 = ~(s2 ? tmp20120 : tmp20830);
  assign tmp20828 = ~(s3 ? tmp20803 : tmp20829);
  assign tmp20824 = s4 ? tmp20825 : tmp20828;
  assign tmp20833 = s2 ? tmp20293 : tmp20152;
  assign tmp20834 = ~(s2 ? 1 : tmp19954);
  assign tmp20832 = s3 ? tmp20833 : tmp20834;
  assign tmp20831 = s4 ? tmp20832 : tmp20120;
  assign tmp20823 = s5 ? tmp20824 : tmp20831;
  assign tmp20819 = s6 ? tmp20820 : tmp20823;
  assign tmp20787 = s7 ? tmp20788 : tmp20819;
  assign tmp20841 = s1 ? tmp19637 : tmp20154;
  assign tmp20840 = s2 ? tmp20841 : tmp20815;
  assign tmp20843 = s1 ? tmp20158 : tmp20302;
  assign tmp20842 = s2 ? tmp20843 : tmp20818;
  assign tmp20839 = s3 ? tmp20840 : tmp20842;
  assign tmp20838 = s4 ? tmp20808 : tmp20839;
  assign tmp20837 = s5 ? tmp20798 : tmp20838;
  assign tmp20836 = s6 ? tmp20789 : tmp20837;
  assign tmp20848 = s2 ? tmp20293 : 1;
  assign tmp20847 = s3 ? tmp20848 : tmp20834;
  assign tmp20851 = s1 ? tmp19635 : tmp20120;
  assign tmp20850 = s2 ? tmp20851 : tmp20120;
  assign tmp20849 = s3 ? tmp20850 : tmp20851;
  assign tmp20846 = s4 ? tmp20847 : tmp20849;
  assign tmp20845 = s5 ? tmp20824 : tmp20846;
  assign tmp20844 = s6 ? tmp20820 : tmp20845;
  assign tmp20835 = s7 ? tmp20836 : tmp20844;
  assign tmp20786 = s8 ? tmp20787 : tmp20835;
  assign tmp20856 = s4 ? tmp20847 : tmp20120;
  assign tmp20855 = s5 ? tmp20824 : tmp20856;
  assign tmp20854 = s6 ? tmp20820 : tmp20855;
  assign tmp20853 = s7 ? tmp20788 : tmp20854;
  assign tmp20852 = s8 ? tmp20835 : tmp20853;
  assign tmp20785 = s9 ? tmp20786 : tmp20852;
  assign tmp20863 = s3 ? tmp20120 : tmp20851;
  assign tmp20862 = s4 ? tmp20847 : tmp20863;
  assign tmp20861 = s5 ? tmp20824 : tmp20862;
  assign tmp20860 = s6 ? tmp20820 : tmp20861;
  assign tmp20859 = s7 ? tmp20788 : tmp20860;
  assign tmp20858 = s8 ? tmp20859 : tmp20788;
  assign tmp20868 = s4 ? tmp20832 : tmp20863;
  assign tmp20867 = s5 ? tmp20824 : tmp20868;
  assign tmp20866 = s6 ? tmp20820 : tmp20867;
  assign tmp20865 = s7 ? tmp20866 : tmp20854;
  assign tmp20869 = s7 ? tmp20844 : tmp20860;
  assign tmp20864 = s8 ? tmp20865 : tmp20869;
  assign tmp20857 = s9 ? tmp20858 : tmp20864;
  assign tmp20784 = s10 ? tmp20785 : tmp20857;
  assign tmp20873 = s7 ? tmp20819 : tmp20854;
  assign tmp20872 = s8 ? tmp20873 : tmp20869;
  assign tmp20871 = s9 ? tmp20858 : tmp20872;
  assign tmp20870 = s10 ? tmp20785 : tmp20871;
  assign tmp20783 = s11 ? tmp20784 : tmp20870;
  assign tmp20645 = s12 ? tmp20646 : tmp20783;
  assign tmp20887 = ~(l4 ? 1 : 0);
  assign tmp20886 = l3 ? 1 : tmp20887;
  assign tmp20885 = ~(l2 ? 1 : tmp20886);
  assign tmp20884 = l1 ? tmp19635 : tmp20885;
  assign tmp20888 = s0 ? 1 : tmp20884;
  assign tmp20883 = s1 ? tmp20884 : tmp20888;
  assign tmp20890 = s1 ? tmp20120 : tmp20884;
  assign tmp20889 = s2 ? tmp20884 : tmp20890;
  assign tmp20882 = s3 ? tmp20883 : tmp20889;
  assign tmp20895 = l1 ? 1 : tmp20885;
  assign tmp20894 = s0 ? tmp20895 : 1;
  assign tmp20893 = s1 ? tmp20894 : tmp20884;
  assign tmp20897 = s0 ? tmp20884 : tmp19614;
  assign tmp20896 = s1 ? tmp20897 : 1;
  assign tmp20892 = s2 ? tmp20893 : tmp20896;
  assign tmp20899 = s1 ? 1 : tmp19717;
  assign tmp20901 = s0 ? tmp20073 : tmp20884;
  assign tmp20900 = s1 ? tmp20884 : tmp20901;
  assign tmp20898 = s2 ? tmp20899 : tmp20900;
  assign tmp20891 = s3 ? tmp20892 : tmp20898;
  assign tmp20881 = s4 ? tmp20882 : tmp20891;
  assign tmp20907 = s0 ? tmp20884 : 1;
  assign tmp20906 = s1 ? tmp20907 : 1;
  assign tmp20908 = s1 ? tmp20888 : tmp20884;
  assign tmp20905 = s2 ? tmp20906 : tmp20908;
  assign tmp20910 = s1 ? tmp20692 : tmp20884;
  assign tmp20909 = s2 ? tmp20884 : tmp20910;
  assign tmp20904 = s3 ? tmp20905 : tmp20909;
  assign tmp20915 = ~(l1 ? tmp19635 : tmp20885);
  assign tmp20914 = s0 ? 1 : tmp20915;
  assign tmp20913 = s1 ? tmp20914 : 0;
  assign tmp20916 = ~(s1 ? 1 : tmp20894);
  assign tmp20912 = s2 ? tmp20913 : tmp20916;
  assign tmp20917 = ~(s2 ? tmp20883 : 0);
  assign tmp20911 = ~(s3 ? tmp20912 : tmp20917);
  assign tmp20903 = s4 ? tmp20904 : tmp20911;
  assign tmp20922 = s0 ? tmp20884 : 0;
  assign tmp20921 = s1 ? tmp20922 : tmp20081;
  assign tmp20920 = s2 ? tmp20921 : tmp19938;
  assign tmp20926 = ~(l1 ? 1 : tmp20885);
  assign tmp20925 = s0 ? 1 : tmp20926;
  assign tmp20924 = ~(s1 ? 1 : tmp20925);
  assign tmp20923 = s2 ? tmp19939 : tmp20924;
  assign tmp20919 = s3 ? tmp20920 : tmp20923;
  assign tmp20930 = s0 ? tmp20895 : tmp20073;
  assign tmp20929 = s1 ? tmp20930 : tmp20073;
  assign tmp20931 = ~(s1 ? tmp20914 : 0);
  assign tmp20928 = s2 ? tmp20929 : tmp20931;
  assign tmp20934 = ~(s0 ? 1 : tmp20915);
  assign tmp20933 = s1 ? tmp20073 : tmp20934;
  assign tmp20937 = ~(l1 ? tmp19635 : 0);
  assign tmp20936 = s0 ? 1 : tmp20937;
  assign tmp20935 = ~(s1 ? tmp20925 : tmp20936);
  assign tmp20932 = s2 ? tmp20933 : tmp20935;
  assign tmp20927 = s3 ? tmp20928 : tmp20932;
  assign tmp20918 = s4 ? tmp20919 : tmp20927;
  assign tmp20902 = s5 ? tmp20903 : tmp20918;
  assign tmp20880 = s6 ? tmp20881 : tmp20902;
  assign tmp20941 = s2 ? tmp20279 : tmp20900;
  assign tmp20940 = s3 ? tmp20892 : tmp20941;
  assign tmp20939 = s4 ? tmp20882 : tmp20940;
  assign tmp20945 = s2 ? tmp20906 : tmp20884;
  assign tmp20944 = s3 ? tmp20945 : tmp20909;
  assign tmp20947 = s2 ? tmp20913 : tmp20926;
  assign tmp20948 = ~(s2 ? tmp20884 : 0);
  assign tmp20946 = ~(s3 ? tmp20947 : tmp20948);
  assign tmp20943 = s4 ? tmp20944 : tmp20946;
  assign tmp20952 = s1 ? tmp20922 : tmp19635;
  assign tmp20951 = s2 ? tmp20952 : 1;
  assign tmp20954 = s1 ? 1 : tmp20926;
  assign tmp20953 = ~(s2 ? 1 : tmp20954);
  assign tmp20950 = s3 ? tmp20951 : tmp20953;
  assign tmp20956 = s2 ? tmp20073 : tmp20884;
  assign tmp20958 = s1 ? tmp20073 : tmp20884;
  assign tmp20957 = s2 ? tmp20958 : tmp20073;
  assign tmp20955 = s3 ? tmp20956 : tmp20957;
  assign tmp20949 = s4 ? tmp20950 : tmp20955;
  assign tmp20942 = s5 ? tmp20943 : tmp20949;
  assign tmp20938 = s6 ? tmp20939 : tmp20942;
  assign tmp20879 = s7 ? tmp20880 : tmp20938;
  assign tmp20965 = ~(l3 ? 1 : tmp20887);
  assign tmp20964 = l1 ? tmp19635 : tmp20965;
  assign tmp20966 = s0 ? 1 : tmp20964;
  assign tmp20963 = s1 ? tmp20964 : tmp20966;
  assign tmp20968 = s1 ? tmp20125 : tmp20964;
  assign tmp20967 = s2 ? tmp20964 : tmp20968;
  assign tmp20962 = s3 ? tmp20963 : tmp20967;
  assign tmp20973 = l1 ? 1 : tmp20965;
  assign tmp20972 = s0 ? tmp20973 : 1;
  assign tmp20971 = s1 ? tmp20972 : tmp20964;
  assign tmp20975 = s0 ? tmp20964 : tmp19614;
  assign tmp20974 = s1 ? tmp20975 : 1;
  assign tmp20970 = s2 ? tmp20971 : tmp20974;
  assign tmp20978 = s0 ? tmp19635 : tmp20964;
  assign tmp20977 = s1 ? tmp20964 : tmp20978;
  assign tmp20976 = s2 ? tmp20899 : tmp20977;
  assign tmp20969 = s3 ? tmp20970 : tmp20976;
  assign tmp20961 = s4 ? tmp20962 : tmp20969;
  assign tmp20984 = s0 ? tmp20964 : 1;
  assign tmp20983 = s1 ? tmp20984 : 1;
  assign tmp20985 = s1 ? tmp20966 : tmp20984;
  assign tmp20982 = s2 ? tmp20983 : tmp20985;
  assign tmp20987 = s1 ? tmp19649 : tmp20964;
  assign tmp20986 = s2 ? tmp20966 : tmp20987;
  assign tmp20981 = s3 ? tmp20982 : tmp20986;
  assign tmp20992 = ~(l1 ? tmp19635 : tmp20965);
  assign tmp20991 = s0 ? 1 : tmp20992;
  assign tmp20990 = s1 ? tmp20991 : 0;
  assign tmp20993 = ~(s1 ? 1 : tmp20972);
  assign tmp20989 = s2 ? tmp20990 : tmp20993;
  assign tmp20995 = s1 ? tmp20964 : tmp20888;
  assign tmp20994 = ~(s2 ? tmp20995 : 0);
  assign tmp20988 = ~(s3 ? tmp20989 : tmp20994);
  assign tmp20980 = s4 ? tmp20981 : tmp20988;
  assign tmp21000 = s0 ? tmp20964 : 0;
  assign tmp20999 = s1 ? tmp21000 : tmp20302;
  assign tmp20998 = s2 ? tmp20999 : tmp20152;
  assign tmp20997 = s3 ? tmp20998 : tmp20923;
  assign tmp21003 = s1 ? tmp20930 : tmp20085;
  assign tmp21004 = ~(s1 ? tmp20991 : 0);
  assign tmp21002 = s2 ? tmp21003 : tmp21004;
  assign tmp21007 = s0 ? tmp20120 : tmp20073;
  assign tmp21006 = s1 ? tmp21007 : tmp20934;
  assign tmp21005 = s2 ? tmp21006 : tmp20935;
  assign tmp21001 = s3 ? tmp21002 : tmp21005;
  assign tmp20996 = s4 ? tmp20997 : tmp21001;
  assign tmp20979 = s5 ? tmp20980 : tmp20996;
  assign tmp20960 = s6 ? tmp20961 : tmp20979;
  assign tmp21011 = s2 ? tmp20279 : tmp20977;
  assign tmp21010 = s3 ? tmp20970 : tmp21011;
  assign tmp21009 = s4 ? tmp20962 : tmp21010;
  assign tmp21016 = s1 ? tmp20964 : tmp20984;
  assign tmp21015 = s2 ? tmp20983 : tmp21016;
  assign tmp21017 = s2 ? tmp20964 : tmp20987;
  assign tmp21014 = s3 ? tmp21015 : tmp21017;
  assign tmp21020 = ~(l1 ? 1 : tmp20965);
  assign tmp21019 = s2 ? tmp20990 : tmp21020;
  assign tmp21022 = s1 ? tmp20964 : tmp20884;
  assign tmp21021 = ~(s2 ? tmp21022 : 0);
  assign tmp21018 = ~(s3 ? tmp21019 : tmp21021);
  assign tmp21013 = s4 ? tmp21014 : tmp21018;
  assign tmp21026 = s1 ? tmp21000 : tmp20120;
  assign tmp21025 = s2 ? tmp21026 : 1;
  assign tmp21024 = s3 ? tmp21025 : tmp20953;
  assign tmp21029 = s1 ? tmp20073 : tmp20085;
  assign tmp21028 = s2 ? tmp21029 : tmp20964;
  assign tmp21027 = s3 ? tmp21028 : tmp20957;
  assign tmp21023 = s4 ? tmp21024 : tmp21027;
  assign tmp21012 = s5 ? tmp21013 : tmp21023;
  assign tmp21008 = s6 ? tmp21009 : tmp21012;
  assign tmp20959 = s7 ? tmp20960 : tmp21008;
  assign tmp20878 = s8 ? tmp20879 : tmp20959;
  assign tmp21036 = s0 ? 1 : tmp20073;
  assign tmp21035 = s1 ? tmp20073 : tmp21036;
  assign tmp21038 = s1 ? tmp19896 : tmp20073;
  assign tmp21037 = s2 ? tmp20073 : tmp21038;
  assign tmp21034 = s3 ? tmp21035 : tmp21037;
  assign tmp21041 = s1 ? tmp19622 : tmp20073;
  assign tmp21043 = s0 ? tmp20073 : tmp19614;
  assign tmp21042 = s1 ? tmp21043 : 1;
  assign tmp21040 = s2 ? tmp21041 : tmp21042;
  assign tmp21044 = s2 ? tmp20899 : tmp20073;
  assign tmp21039 = s3 ? tmp21040 : tmp21044;
  assign tmp21033 = s4 ? tmp21034 : tmp21039;
  assign tmp21049 = s1 ? tmp21036 : tmp20111;
  assign tmp21048 = s2 ? tmp20110 : tmp21049;
  assign tmp21051 = s1 ? tmp20692 : tmp20073;
  assign tmp21050 = s2 ? tmp21036 : tmp21051;
  assign tmp21047 = s3 ? tmp21048 : tmp21050;
  assign tmp21054 = s1 ? tmp20936 : 0;
  assign tmp21053 = s2 ? tmp21054 : tmp19721;
  assign tmp21057 = s0 ? tmp19614 : tmp20073;
  assign tmp21056 = s1 ? tmp20073 : tmp21057;
  assign tmp21055 = ~(s2 ? tmp21056 : 0);
  assign tmp21052 = ~(s3 ? tmp21053 : tmp21055);
  assign tmp21046 = s4 ? tmp21047 : tmp21052;
  assign tmp21061 = s1 ? tmp20692 : tmp20081;
  assign tmp21060 = s2 ? tmp21061 : tmp19635;
  assign tmp21059 = s3 ? tmp21060 : tmp20009;
  assign tmp21064 = ~(s1 ? tmp20936 : 0);
  assign tmp21063 = s2 ? tmp20073 : tmp21064;
  assign tmp21067 = ~(s0 ? 1 : tmp20937);
  assign tmp21066 = s1 ? tmp20073 : tmp21067;
  assign tmp21065 = s2 ? tmp21066 : tmp21067;
  assign tmp21062 = s3 ? tmp21063 : tmp21065;
  assign tmp21058 = s4 ? tmp21059 : tmp21062;
  assign tmp21045 = s5 ? tmp21046 : tmp21058;
  assign tmp21032 = s6 ? tmp21033 : tmp21045;
  assign tmp21071 = s2 ? tmp20279 : tmp20073;
  assign tmp21070 = s3 ? tmp21040 : tmp21071;
  assign tmp21069 = s4 ? tmp21034 : tmp21070;
  assign tmp21076 = s1 ? tmp20073 : tmp20111;
  assign tmp21075 = s2 ? tmp20110 : tmp21076;
  assign tmp21077 = s2 ? tmp20073 : tmp21051;
  assign tmp21074 = s3 ? tmp21075 : tmp21077;
  assign tmp21079 = s2 ? tmp21054 : tmp19720;
  assign tmp21080 = ~(s2 ? tmp20073 : 0);
  assign tmp21078 = ~(s3 ? tmp21079 : tmp21080);
  assign tmp21073 = s4 ? tmp21074 : tmp21078;
  assign tmp21084 = s1 ? tmp20692 : tmp19635;
  assign tmp21083 = s2 ? tmp21084 : 1;
  assign tmp21082 = s3 ? tmp21083 : tmp20028;
  assign tmp21081 = s4 ? tmp21082 : tmp20073;
  assign tmp21072 = s5 ? tmp21073 : tmp21081;
  assign tmp21068 = s6 ? tmp21069 : tmp21072;
  assign tmp21031 = s7 ? tmp21032 : tmp21068;
  assign tmp21030 = s8 ? tmp20959 : tmp21031;
  assign tmp20877 = s9 ? tmp20878 : tmp21030;
  assign tmp21092 = s1 ? tmp20125 : tmp20884;
  assign tmp21091 = s2 ? tmp20884 : tmp21092;
  assign tmp21090 = s3 ? tmp20883 : tmp21091;
  assign tmp21097 = ~(l2 ? tmp20886 : 1);
  assign tmp21096 = s0 ? tmp20884 : tmp21097;
  assign tmp21095 = s1 ? tmp21096 : 1;
  assign tmp21094 = s2 ? tmp20893 : tmp21095;
  assign tmp21093 = s3 ? tmp21094 : tmp20898;
  assign tmp21089 = s4 ? tmp21090 : tmp21093;
  assign tmp21102 = s1 ? tmp20888 : tmp20907;
  assign tmp21101 = s2 ? tmp20906 : tmp21102;
  assign tmp21103 = s2 ? tmp20888 : tmp20910;
  assign tmp21100 = s3 ? tmp21101 : tmp21103;
  assign tmp21107 = s0 ? tmp19614 : tmp20884;
  assign tmp21106 = s1 ? tmp20884 : tmp21107;
  assign tmp21105 = ~(s2 ? tmp21106 : 0);
  assign tmp21104 = ~(s3 ? tmp20912 : tmp21105);
  assign tmp21099 = s4 ? tmp21100 : tmp21104;
  assign tmp21098 = s5 ? tmp21099 : tmp20918;
  assign tmp21088 = s6 ? tmp21089 : tmp21098;
  assign tmp21110 = s3 ? tmp21094 : tmp20941;
  assign tmp21109 = s4 ? tmp21090 : tmp21110;
  assign tmp21115 = s1 ? tmp20884 : tmp20907;
  assign tmp21114 = s2 ? tmp20906 : tmp21115;
  assign tmp21113 = s3 ? tmp21114 : tmp20909;
  assign tmp21112 = s4 ? tmp21113 : tmp20946;
  assign tmp21111 = s5 ? tmp21112 : tmp20949;
  assign tmp21108 = s6 ? tmp21109 : tmp21111;
  assign tmp21087 = s7 ? tmp21088 : tmp21108;
  assign tmp21086 = s8 ? tmp21087 : tmp21088;
  assign tmp21121 = s3 ? tmp20956 : tmp20958;
  assign tmp21120 = s4 ? tmp20950 : tmp21121;
  assign tmp21119 = s5 ? tmp20943 : tmp21120;
  assign tmp21118 = s6 ? tmp20939 : tmp21119;
  assign tmp21117 = s7 ? tmp21118 : tmp21068;
  assign tmp21126 = s3 ? tmp21028 : tmp20958;
  assign tmp21125 = s4 ? tmp21024 : tmp21126;
  assign tmp21124 = s5 ? tmp21013 : tmp21125;
  assign tmp21123 = s6 ? tmp21009 : tmp21124;
  assign tmp21128 = s5 ? tmp21112 : tmp21120;
  assign tmp21127 = s6 ? tmp21109 : tmp21128;
  assign tmp21122 = s7 ? tmp21123 : tmp21127;
  assign tmp21116 = s8 ? tmp21117 : tmp21122;
  assign tmp21085 = s9 ? tmp21086 : tmp21116;
  assign tmp20876 = s10 ? tmp20877 : tmp21085;
  assign tmp21132 = s7 ? tmp20938 : tmp21068;
  assign tmp21133 = s7 ? tmp21008 : tmp21108;
  assign tmp21131 = s8 ? tmp21132 : tmp21133;
  assign tmp21130 = s9 ? tmp21086 : tmp21131;
  assign tmp21129 = s10 ? tmp20877 : tmp21130;
  assign tmp20875 = ~(s11 ? tmp20876 : tmp21129);
  assign tmp20874 = ~(s12 ? 1 : tmp20875);
  assign tmp20644 = s13 ? tmp20645 : tmp20874;
  assign tmp20361 = ~(s14 ? tmp20362 : tmp20644);
  assign tmp19599 = s15 ? tmp19600 : tmp20361;
  assign tmp21146 = s2 ? tmp19644 : tmp19650;
  assign tmp21145 = s3 ? tmp21146 : 0;
  assign tmp21144 = ~(s4 ? tmp21145 : tmp19672);
  assign tmp21143 = s5 ? tmp19629 : tmp21144;
  assign tmp21142 = s6 ? tmp19608 : tmp21143;
  assign tmp21150 = s3 ? tmp19644 : 0;
  assign tmp21149 = ~(s4 ? tmp21150 : tmp19672);
  assign tmp21148 = s5 ? tmp19661 : tmp21149;
  assign tmp21147 = s6 ? tmp19656 : tmp21148;
  assign tmp21141 = s7 ? tmp21142 : tmp21147;
  assign tmp21158 = s0 ? tmp19611 : 0;
  assign tmp21157 = s1 ? tmp19613 : tmp21158;
  assign tmp21156 = s2 ? tmp19632 : tmp21157;
  assign tmp21161 = s0 ? 1 : tmp19783;
  assign tmp21160 = s1 ? tmp21161 : tmp19637;
  assign tmp21159 = ~(s2 ? tmp21160 : tmp19638);
  assign tmp21155 = s3 ? tmp21156 : tmp21159;
  assign tmp21154 = s4 ? tmp21155 : tmp19689;
  assign tmp21153 = s5 ? tmp21154 : tmp21144;
  assign tmp21152 = s6 ? tmp19676 : tmp21153;
  assign tmp21167 = s1 ? tmp19611 : tmp21158;
  assign tmp21166 = s2 ? tmp19616 : tmp21167;
  assign tmp21165 = s3 ? tmp21166 : tmp19699;
  assign tmp21171 = ~(s0 ? tmp19611 : tmp20122);
  assign tmp21170 = ~(s1 ? tmp20120 : tmp21171);
  assign tmp21169 = s2 ? tmp19641 : tmp21170;
  assign tmp21168 = s3 ? tmp21169 : tmp19690;
  assign tmp21164 = s4 ? tmp21165 : tmp21168;
  assign tmp21163 = s5 ? tmp21164 : tmp21149;
  assign tmp21162 = s6 ? tmp19692 : tmp21163;
  assign tmp21151 = s7 ? tmp21152 : tmp21162;
  assign tmp21140 = s8 ? tmp21141 : tmp21151;
  assign tmp21177 = s2 ? tmp20120 : tmp20158;
  assign tmp21179 = s1 ? tmp20120 : tmp19649;
  assign tmp21178 = s2 ? tmp21179 : tmp20817;
  assign tmp21176 = s3 ? tmp21177 : tmp21178;
  assign tmp21175 = s4 ? tmp20120 : tmp21176;
  assign tmp21184 = s1 ? tmp20129 : tmp20121;
  assign tmp21185 = ~(s1 ? tmp20805 : tmp20122);
  assign tmp21183 = s2 ? tmp21184 : tmp21185;
  assign tmp21187 = s1 ? tmp20120 : tmp19719;
  assign tmp21189 = ~(s0 ? tmp20120 : tmp19635);
  assign tmp21188 = ~(s1 ? 1 : tmp21189);
  assign tmp21186 = s2 ? tmp21187 : tmp21188;
  assign tmp21182 = s3 ? tmp21183 : tmp21186;
  assign tmp21192 = s1 ? tmp20304 : tmp21189;
  assign tmp21193 = ~(s1 ? tmp20158 : tmp20120);
  assign tmp21191 = s2 ? tmp21192 : tmp21193;
  assign tmp21194 = s2 ? tmp20393 : 1;
  assign tmp21190 = ~(s3 ? tmp21191 : tmp21194);
  assign tmp21181 = s4 ? tmp21182 : tmp21190;
  assign tmp21197 = s2 ? tmp19624 : tmp19731;
  assign tmp21196 = s3 ? tmp21197 : 1;
  assign tmp21195 = ~(s4 ? tmp21196 : tmp19746);
  assign tmp21180 = s5 ? tmp21181 : tmp21195;
  assign tmp21174 = s6 ? tmp21175 : tmp21180;
  assign tmp21202 = s1 ? tmp20158 : tmp20120;
  assign tmp21201 = s2 ? tmp20120 : tmp21202;
  assign tmp21203 = s2 ? tmp20384 : tmp20817;
  assign tmp21200 = s3 ? tmp21201 : tmp21203;
  assign tmp21199 = s4 ? tmp20120 : tmp21200;
  assign tmp21207 = s2 ? tmp20128 : tmp20120;
  assign tmp21209 = s1 ? tmp20120 : tmp19720;
  assign tmp21208 = s2 ? tmp21209 : tmp21188;
  assign tmp21206 = s3 ? tmp21207 : tmp21208;
  assign tmp21211 = s2 ? tmp21192 : tmp20122;
  assign tmp21213 = s1 ? tmp19687 : 1;
  assign tmp21212 = s2 ? tmp21213 : 1;
  assign tmp21210 = ~(s3 ? tmp21211 : tmp21212);
  assign tmp21205 = s4 ? tmp21206 : tmp21210;
  assign tmp21215 = s3 ? tmp19624 : 1;
  assign tmp21214 = ~(s4 ? tmp21215 : tmp19746);
  assign tmp21204 = s5 ? tmp21205 : tmp21214;
  assign tmp21198 = s6 ? tmp21199 : tmp21204;
  assign tmp21173 = ~(s7 ? tmp21174 : tmp21198);
  assign tmp21172 = s8 ? tmp21151 : tmp21173;
  assign tmp21139 = s9 ? tmp21140 : tmp21172;
  assign tmp21223 = s1 ? tmp20154 : tmp19635;
  assign tmp21222 = s2 ? tmp19635 : tmp21223;
  assign tmp21221 = s3 ? tmp20718 : tmp21222;
  assign tmp21225 = s2 ? tmp21223 : tmp20718;
  assign tmp21226 = s2 ? tmp21179 : tmp20269;
  assign tmp21224 = s3 ? tmp21225 : tmp21226;
  assign tmp21220 = s4 ? tmp21221 : tmp21224;
  assign tmp21231 = s1 ? tmp20062 : tmp19917;
  assign tmp21232 = ~(s1 ? tmp19687 : tmp19634);
  assign tmp21230 = s2 ? tmp21231 : tmp21232;
  assign tmp21235 = ~(s0 ? tmp19635 : tmp20073);
  assign tmp21234 = ~(s1 ? 1 : tmp21235);
  assign tmp21233 = s2 ? tmp19637 : tmp21234;
  assign tmp21229 = s3 ? tmp21230 : tmp21233;
  assign tmp21238 = s1 ? tmp19651 : tmp21189;
  assign tmp21239 = ~(s1 ? tmp20158 : tmp20154);
  assign tmp21237 = s2 ? tmp21238 : tmp21239;
  assign tmp21241 = s1 ? tmp20072 : tmp19649;
  assign tmp21240 = ~(s2 ? tmp21241 : 0);
  assign tmp21236 = ~(s3 ? tmp21237 : tmp21240);
  assign tmp21228 = s4 ? tmp21229 : tmp21236;
  assign tmp21242 = s4 ? tmp21145 : tmp19672;
  assign tmp21227 = s5 ? tmp21228 : tmp21242;
  assign tmp21219 = s6 ? tmp21220 : tmp21227;
  assign tmp21246 = s2 ? tmp21223 : tmp20851;
  assign tmp21247 = s2 ? tmp20384 : tmp20269;
  assign tmp21245 = s3 ? tmp21246 : tmp21247;
  assign tmp21244 = s4 ? tmp21221 : tmp21245;
  assign tmp21251 = s2 ? tmp20061 : tmp20099;
  assign tmp21252 = s2 ? tmp19635 : tmp21234;
  assign tmp21250 = s3 ? tmp21251 : tmp21252;
  assign tmp21255 = ~(s1 ? tmp20120 : tmp20154);
  assign tmp21254 = s2 ? tmp21238 : tmp21255;
  assign tmp21257 = s1 ? tmp20072 : 0;
  assign tmp21256 = ~(s2 ? tmp21257 : 0);
  assign tmp21253 = ~(s3 ? tmp21254 : tmp21256);
  assign tmp21249 = s4 ? tmp21250 : tmp21253;
  assign tmp21258 = s4 ? tmp21150 : tmp19672;
  assign tmp21248 = s5 ? tmp21249 : tmp21258;
  assign tmp21243 = s6 ? tmp21244 : tmp21248;
  assign tmp21218 = s7 ? tmp21219 : tmp21243;
  assign tmp21217 = s8 ? tmp21218 : tmp21219;
  assign tmp21262 = s5 ? tmp19759 : tmp21149;
  assign tmp21261 = s6 ? tmp19656 : tmp21262;
  assign tmp21263 = ~(s6 ? tmp21199 : tmp21204);
  assign tmp21260 = s7 ? tmp21261 : tmp21263;
  assign tmp21270 = ~(s1 ? tmp20120 : tmp19783);
  assign tmp21269 = s2 ? tmp19641 : tmp21270;
  assign tmp21268 = s3 ? tmp21269 : tmp19690;
  assign tmp21267 = s4 ? tmp21165 : tmp21268;
  assign tmp21266 = s5 ? tmp21267 : tmp21149;
  assign tmp21265 = s6 ? tmp19692 : tmp21266;
  assign tmp21276 = ~(s1 ? tmp20120 : tmp19635);
  assign tmp21275 = s2 ? tmp21238 : tmp21276;
  assign tmp21274 = ~(s3 ? tmp21275 : tmp21256);
  assign tmp21273 = s4 ? tmp21250 : tmp21274;
  assign tmp21272 = s5 ? tmp21273 : tmp21258;
  assign tmp21271 = ~(s6 ? tmp21244 : tmp21272);
  assign tmp21264 = s7 ? tmp21265 : tmp21271;
  assign tmp21259 = ~(s8 ? tmp21260 : tmp21264);
  assign tmp21216 = ~(s9 ? tmp21217 : tmp21259);
  assign tmp21138 = s10 ? tmp21139 : tmp21216;
  assign tmp21280 = s7 ? tmp21147 : tmp21263;
  assign tmp21282 = ~(s6 ? tmp21244 : tmp21248);
  assign tmp21281 = s7 ? tmp21162 : tmp21282;
  assign tmp21279 = ~(s8 ? tmp21280 : tmp21281);
  assign tmp21278 = ~(s9 ? tmp21217 : tmp21279);
  assign tmp21277 = s10 ? tmp21139 : tmp21278;
  assign tmp21137 = s11 ? tmp21138 : tmp21277;
  assign tmp21293 = s1 ? 1 : tmp19813;
  assign tmp21292 = s2 ? tmp20259 : tmp21293;
  assign tmp21291 = s3 ? 1 : tmp21292;
  assign tmp21290 = s4 ? 1 : tmp21291;
  assign tmp21298 = ~(s1 ? 1 : tmp19813);
  assign tmp21297 = s2 ? tmp20259 : tmp21298;
  assign tmp21296 = s3 ? 1 : tmp21297;
  assign tmp21301 = ~(s1 ? tmp19780 : 1);
  assign tmp21300 = s2 ? tmp19812 : tmp21301;
  assign tmp21299 = ~(s3 ? tmp21300 : 1);
  assign tmp21295 = s4 ? tmp21296 : tmp21299;
  assign tmp21294 = s5 ? tmp21295 : 0;
  assign tmp21289 = s6 ? tmp21290 : tmp21294;
  assign tmp21306 = s2 ? tmp20279 : tmp21298;
  assign tmp21305 = s3 ? 1 : tmp21306;
  assign tmp21308 = s2 ? tmp19812 : 0;
  assign tmp21307 = ~(s3 ? tmp21308 : 1);
  assign tmp21304 = s4 ? tmp21305 : tmp21307;
  assign tmp21303 = s5 ? tmp21304 : 0;
  assign tmp21302 = s6 ? tmp21290 : tmp21303;
  assign tmp21288 = s7 ? tmp21289 : tmp21302;
  assign tmp21315 = ~(s1 ? 1 : 0);
  assign tmp21314 = s2 ? tmp20259 : tmp21315;
  assign tmp21313 = s3 ? 1 : tmp21314;
  assign tmp21317 = s2 ? tmp19939 : 0;
  assign tmp21316 = ~(s3 ? tmp21317 : 1);
  assign tmp21312 = s4 ? tmp21313 : tmp21316;
  assign tmp21311 = s5 ? tmp21312 : 0;
  assign tmp21310 = s6 ? tmp21290 : tmp21311;
  assign tmp21322 = s1 ? 1 : tmp20936;
  assign tmp21321 = s2 ? 1 : tmp21322;
  assign tmp21325 = ~(s0 ? tmp20073 : 1);
  assign tmp21324 = s1 ? 1 : tmp21325;
  assign tmp21323 = s2 ? tmp21324 : tmp21293;
  assign tmp21320 = s3 ? tmp21321 : tmp21323;
  assign tmp21319 = s4 ? 1 : tmp21320;
  assign tmp21329 = s2 ? tmp20279 : tmp21315;
  assign tmp21328 = s3 ? 1 : tmp21329;
  assign tmp21327 = s4 ? tmp21328 : tmp21316;
  assign tmp21326 = s5 ? tmp21327 : 0;
  assign tmp21318 = s6 ? tmp21319 : tmp21326;
  assign tmp21309 = s7 ? tmp21310 : tmp21318;
  assign tmp21287 = s8 ? tmp21288 : tmp21309;
  assign tmp21335 = s2 ? tmp21076 : tmp21035;
  assign tmp21334 = s3 ? tmp20073 : tmp21335;
  assign tmp21333 = s4 ? tmp20073 : tmp21334;
  assign tmp21340 = s1 ? tmp20692 : tmp21067;
  assign tmp21341 = ~(s1 ? tmp19651 : tmp19720);
  assign tmp21339 = s2 ? tmp21340 : tmp21341;
  assign tmp21343 = s1 ? tmp19614 : tmp19622;
  assign tmp21342 = s2 ? tmp21343 : tmp19888;
  assign tmp21338 = s3 ? tmp21339 : tmp21342;
  assign tmp21345 = s2 ? tmp20274 : tmp19635;
  assign tmp21344 = s3 ? tmp21345 : 1;
  assign tmp21337 = s4 ? tmp21338 : tmp21344;
  assign tmp21336 = s5 ? tmp21337 : 1;
  assign tmp21332 = s6 ? tmp21333 : tmp21336;
  assign tmp21351 = s1 ? tmp19635 : tmp19614;
  assign tmp21350 = s2 ? tmp21051 : tmp21351;
  assign tmp21352 = s2 ? tmp19624 : tmp19888;
  assign tmp21349 = s3 ? tmp21350 : tmp21352;
  assign tmp21348 = s4 ? tmp21349 : tmp21344;
  assign tmp21347 = s5 ? tmp21348 : 1;
  assign tmp21346 = s6 ? tmp21333 : tmp21347;
  assign tmp21331 = ~(s7 ? tmp21332 : tmp21346);
  assign tmp21330 = s8 ? tmp21309 : tmp21331;
  assign tmp21286 = s9 ? tmp21287 : tmp21330;
  assign tmp21355 = s7 ? tmp21332 : tmp21346;
  assign tmp21354 = s8 ? tmp21355 : tmp21332;
  assign tmp21361 = s2 ? tmp20279 : tmp21293;
  assign tmp21360 = s3 ? 1 : tmp21361;
  assign tmp21359 = s4 ? 1 : tmp21360;
  assign tmp21358 = s6 ? tmp21359 : tmp21303;
  assign tmp21366 = s1 ? tmp20073 : 1;
  assign tmp21365 = s2 ? tmp21366 : tmp21035;
  assign tmp21364 = s3 ? tmp20073 : tmp21365;
  assign tmp21363 = s4 ? tmp20073 : tmp21364;
  assign tmp21362 = ~(s6 ? tmp21363 : tmp21347);
  assign tmp21357 = s7 ? tmp21358 : tmp21362;
  assign tmp21370 = s3 ? tmp21321 : tmp21361;
  assign tmp21369 = s4 ? 1 : tmp21370;
  assign tmp21368 = s6 ? tmp21369 : tmp21326;
  assign tmp21367 = s7 ? tmp21368 : tmp21362;
  assign tmp21356 = ~(s8 ? tmp21357 : tmp21367);
  assign tmp21353 = ~(s9 ? tmp21354 : tmp21356);
  assign tmp21285 = s10 ? tmp21286 : tmp21353;
  assign tmp21375 = ~(s6 ? tmp21333 : tmp21347);
  assign tmp21374 = s7 ? tmp21302 : tmp21375;
  assign tmp21376 = s7 ? tmp21318 : tmp21375;
  assign tmp21373 = ~(s8 ? tmp21374 : tmp21376);
  assign tmp21372 = ~(s9 ? tmp21354 : tmp21373);
  assign tmp21371 = s10 ? tmp21286 : tmp21372;
  assign tmp21284 = s11 ? tmp21285 : tmp21371;
  assign tmp21283 = s12 ? tmp19769 : tmp21284;
  assign tmp21136 = s13 ? tmp21137 : tmp21283;
  assign tmp21387 = s2 ? tmp20432 : tmp20434;
  assign tmp21389 = s1 ? tmp20432 : tmp19622;
  assign tmp21390 = s1 ? tmp20432 : tmp20447;
  assign tmp21388 = s2 ? tmp21389 : tmp21390;
  assign tmp21386 = s3 ? tmp21387 : tmp21388;
  assign tmp21385 = s4 ? tmp20432 : tmp21386;
  assign tmp21396 = s0 ? tmp20432 : tmp19635;
  assign tmp21397 = s0 ? tmp19635 : tmp20432;
  assign tmp21395 = s1 ? tmp21396 : tmp21397;
  assign tmp21398 = s1 ? tmp19896 : tmp20432;
  assign tmp21394 = s2 ? tmp21395 : tmp21398;
  assign tmp21401 = s0 ? tmp20432 : 1;
  assign tmp21400 = s1 ? tmp20432 : tmp21401;
  assign tmp21399 = s2 ? tmp21400 : 1;
  assign tmp21393 = s3 ? tmp21394 : tmp21399;
  assign tmp21392 = s4 ? tmp21393 : 1;
  assign tmp21391 = s5 ? tmp21392 : 1;
  assign tmp21384 = s6 ? tmp21385 : tmp21391;
  assign tmp21406 = s1 ? tmp20434 : 1;
  assign tmp21405 = s2 ? tmp20432 : tmp21406;
  assign tmp21408 = s1 ? tmp20432 : 1;
  assign tmp21407 = s2 ? tmp21408 : tmp21390;
  assign tmp21404 = s3 ? tmp21405 : tmp21407;
  assign tmp21403 = s4 ? tmp20432 : tmp21404;
  assign tmp21413 = s1 ? tmp21396 : tmp20432;
  assign tmp21414 = s1 ? 1 : tmp20432;
  assign tmp21412 = s2 ? tmp21413 : tmp21414;
  assign tmp21411 = s3 ? tmp21412 : tmp21399;
  assign tmp21410 = s4 ? tmp21411 : 1;
  assign tmp21409 = s5 ? tmp21410 : 1;
  assign tmp21402 = s6 ? tmp21403 : tmp21409;
  assign tmp21383 = s7 ? tmp21384 : tmp21402;
  assign tmp21382 = s8 ? tmp19868 : tmp21383;
  assign tmp21381 = s9 ? tmp21382 : tmp21383;
  assign tmp21416 = s8 ? tmp21383 : tmp21384;
  assign tmp21423 = s2 ? tmp21408 : 1;
  assign tmp21422 = s3 ? tmp21412 : tmp21423;
  assign tmp21421 = s4 ? tmp21422 : 1;
  assign tmp21420 = s5 ? tmp21421 : 1;
  assign tmp21419 = s6 ? tmp21403 : tmp21420;
  assign tmp21418 = s7 ? tmp19901 : tmp21419;
  assign tmp21417 = s8 ? tmp21418 : tmp21419;
  assign tmp21415 = s9 ? tmp21416 : tmp21417;
  assign tmp21380 = s10 ? tmp21381 : tmp21415;
  assign tmp21427 = s7 ? tmp19880 : tmp21402;
  assign tmp21426 = s8 ? tmp21427 : tmp21402;
  assign tmp21425 = s9 ? tmp21416 : tmp21426;
  assign tmp21424 = s10 ? tmp21381 : tmp21425;
  assign tmp21379 = s11 ? tmp21380 : tmp21424;
  assign tmp21436 = s2 ? tmp19919 : tmp20063;
  assign tmp21435 = s3 ? tmp21436 : tmp19953;
  assign tmp21434 = s4 ? tmp20058 : tmp21435;
  assign tmp21441 = s1 ? tmp19896 : tmp19780;
  assign tmp21440 = s2 ? tmp21441 : tmp20069;
  assign tmp21442 = s2 ? tmp19637 : tmp19888;
  assign tmp21439 = s3 ? tmp21440 : tmp21442;
  assign tmp21438 = s4 ? tmp21439 : tmp19929;
  assign tmp21437 = s5 ? tmp21438 : tmp19935;
  assign tmp21433 = s6 ? tmp21434 : tmp21437;
  assign tmp21446 = s2 ? tmp19919 : tmp20094;
  assign tmp21445 = s3 ? tmp21446 : tmp19953;
  assign tmp21444 = s4 ? tmp20058 : tmp21445;
  assign tmp21451 = s1 ? tmp19896 : 0;
  assign tmp21450 = s2 ? tmp21451 : tmp20099;
  assign tmp21449 = s3 ? tmp21450 : tmp19887;
  assign tmp21448 = s4 ? tmp21449 : tmp19959;
  assign tmp21447 = s5 ? tmp21448 : tmp19962;
  assign tmp21443 = s6 ? tmp21444 : tmp21447;
  assign tmp21432 = s7 ? tmp21433 : tmp21443;
  assign tmp21455 = s3 ? tmp20718 : tmp19894;
  assign tmp21458 = s1 ? tmp19896 : tmp20125;
  assign tmp21457 = s2 ? tmp19635 : tmp21458;
  assign tmp21460 = s1 ? tmp20120 : 1;
  assign tmp21459 = s2 ? tmp21460 : tmp19875;
  assign tmp21456 = s3 ? tmp21457 : tmp21459;
  assign tmp21454 = s4 ? tmp21455 : tmp21456;
  assign tmp21463 = s3 ? tmp20067 : tmp21442;
  assign tmp21465 = s2 ? tmp20814 : tmp20173;
  assign tmp21466 = s2 ? tmp20718 : 1;
  assign tmp21464 = s3 ? tmp21465 : tmp21466;
  assign tmp21462 = s4 ? tmp21463 : tmp21464;
  assign tmp21469 = s2 ? tmp19938 : tmp20274;
  assign tmp21468 = s3 ? tmp21469 : tmp19940;
  assign tmp21470 = s3 ? tmp21469 : tmp19945;
  assign tmp21467 = s4 ? tmp21468 : tmp21470;
  assign tmp21461 = s5 ? tmp21462 : tmp21467;
  assign tmp21453 = s6 ? tmp21454 : tmp21461;
  assign tmp21475 = s1 ? tmp19896 : tmp20120;
  assign tmp21474 = s2 ? tmp19635 : tmp21475;
  assign tmp21473 = s3 ? tmp21474 : tmp21459;
  assign tmp21472 = s4 ? tmp21455 : tmp21473;
  assign tmp21478 = s3 ? tmp20098 : tmp19887;
  assign tmp21477 = s4 ? tmp21478 : tmp21464;
  assign tmp21481 = s2 ? tmp19938 : tmp19644;
  assign tmp21480 = s3 ? tmp21481 : tmp19965;
  assign tmp21479 = s4 ? tmp21480 : tmp19966;
  assign tmp21476 = s5 ? tmp21477 : tmp21479;
  assign tmp21471 = s6 ? tmp21472 : tmp21476;
  assign tmp21452 = s7 ? tmp21453 : tmp21471;
  assign tmp21431 = s8 ? tmp21432 : tmp21452;
  assign tmp21487 = s2 ? tmp20120 : tmp20125;
  assign tmp21488 = s2 ? tmp21460 : tmp20791;
  assign tmp21486 = s3 ? tmp21487 : tmp21488;
  assign tmp21485 = s4 ? tmp20120 : tmp21486;
  assign tmp21492 = s2 ? tmp20138 : tmp20793;
  assign tmp21493 = s2 ? tmp21187 : tmp20141;
  assign tmp21491 = s3 ? tmp21492 : tmp21493;
  assign tmp21495 = s2 ? tmp20793 : tmp20120;
  assign tmp21497 = s1 ? tmp20805 : tmp20146;
  assign tmp21496 = ~(s2 ? tmp21497 : 0);
  assign tmp21494 = s3 ? tmp21495 : tmp21496;
  assign tmp21490 = s4 ? tmp21491 : tmp21494;
  assign tmp21501 = ~(s1 ? tmp19719 : tmp19720);
  assign tmp21500 = s2 ? tmp20007 : tmp21501;
  assign tmp21499 = s3 ? tmp21500 : tmp20009;
  assign tmp21502 = s3 ? tmp21500 : tmp20014;
  assign tmp21498 = ~(s4 ? tmp21499 : tmp21502);
  assign tmp21489 = s5 ? tmp21490 : tmp21498;
  assign tmp21484 = s6 ? tmp21485 : tmp21489;
  assign tmp21505 = s3 ? tmp20123 : tmp21488;
  assign tmp21504 = s4 ? tmp20120 : tmp21505;
  assign tmp21509 = s2 ? tmp20124 : tmp20120;
  assign tmp21510 = s2 ? tmp21209 : tmp20141;
  assign tmp21508 = s3 ? tmp21509 : tmp21510;
  assign tmp21507 = s4 ? tmp21508 : tmp21494;
  assign tmp21513 = s2 ? tmp20007 : tmp19624;
  assign tmp21512 = s3 ? tmp21513 : tmp20028;
  assign tmp21511 = ~(s4 ? tmp21512 : tmp20030);
  assign tmp21506 = s5 ? tmp21507 : tmp21511;
  assign tmp21503 = s6 ? tmp21504 : tmp21506;
  assign tmp21483 = s7 ? tmp21484 : tmp21503;
  assign tmp21482 = s8 ? tmp21452 : tmp21483;
  assign tmp21430 = s9 ? tmp21431 : tmp21482;
  assign tmp21515 = s8 ? tmp21452 : tmp21453;
  assign tmp21520 = s4 ? tmp21449 : tmp20043;
  assign tmp21519 = s5 ? tmp21520 : tmp19962;
  assign tmp21518 = s6 ? tmp21444 : tmp21519;
  assign tmp21526 = s1 ? tmp20805 : tmp19614;
  assign tmp21525 = ~(s2 ? tmp21526 : 0);
  assign tmp21524 = s3 ? tmp21495 : tmp21525;
  assign tmp21523 = s4 ? tmp21508 : tmp21524;
  assign tmp21522 = s5 ? tmp21523 : tmp21511;
  assign tmp21521 = s6 ? tmp21504 : tmp21522;
  assign tmp21517 = s7 ? tmp21518 : tmp21521;
  assign tmp21530 = s3 ? tmp21465 : tmp19879;
  assign tmp21529 = s4 ? tmp21478 : tmp21530;
  assign tmp21528 = s5 ? tmp21529 : tmp21479;
  assign tmp21527 = s6 ? tmp21472 : tmp21528;
  assign tmp21516 = s8 ? tmp21517 : tmp21527;
  assign tmp21514 = s9 ? tmp21515 : tmp21516;
  assign tmp21429 = s10 ? tmp21430 : tmp21514;
  assign tmp21534 = s7 ? tmp21443 : tmp21503;
  assign tmp21533 = s8 ? tmp21534 : tmp21471;
  assign tmp21532 = s9 ? tmp21515 : tmp21533;
  assign tmp21531 = s10 ? tmp21430 : tmp21532;
  assign tmp21428 = s11 ? tmp21429 : tmp21531;
  assign tmp21378 = s12 ? tmp21379 : tmp21428;
  assign tmp21545 = s1 ? tmp20120 : tmp20081;
  assign tmp21544 = s2 ? tmp21545 : 1;
  assign tmp21543 = s3 ? tmp20143 : tmp21544;
  assign tmp21542 = s4 ? tmp20136 : tmp21543;
  assign tmp21548 = s2 ? tmp20152 : tmp20793;
  assign tmp21547 = s3 ? tmp21548 : tmp20086;
  assign tmp21550 = s2 ? tmp19635 : tmp20793;
  assign tmp21549 = s3 ? tmp21550 : tmp19945;
  assign tmp21546 = s4 ? tmp21547 : tmp21549;
  assign tmp21541 = s5 ? tmp21542 : tmp21546;
  assign tmp21540 = s6 ? tmp20117 : tmp21541;
  assign tmp21554 = s3 ? tmp20176 : tmp19965;
  assign tmp21553 = s4 ? tmp21554 : tmp20233;
  assign tmp21552 = s5 ? tmp20165 : tmp21553;
  assign tmp21551 = s6 ? tmp20160 : tmp21552;
  assign tmp21539 = s7 ? tmp21540 : tmp21551;
  assign tmp21560 = s2 ? tmp19846 : tmp20793;
  assign tmp21559 = s3 ? tmp21560 : tmp19945;
  assign tmp21558 = s4 ? tmp21547 : tmp21559;
  assign tmp21557 = s5 ? tmp20135 : tmp21558;
  assign tmp21556 = s6 ? tmp20117 : tmp21557;
  assign tmp21555 = s7 ? tmp21556 : tmp21551;
  assign tmp21538 = s8 ? tmp21539 : tmp21555;
  assign tmp21565 = s3 ? tmp20127 : tmp20321;
  assign tmp21564 = s4 ? tmp20118 : tmp21565;
  assign tmp21569 = s2 ? tmp20152 : tmp20120;
  assign tmp21568 = s3 ? tmp21569 : tmp20086;
  assign tmp21567 = s4 ? tmp21568 : tmp21559;
  assign tmp21566 = s5 ? tmp20135 : tmp21567;
  assign tmp21563 = s6 ? tmp21564 : tmp21566;
  assign tmp21572 = s3 ? tmp20162 : tmp20321;
  assign tmp21571 = s4 ? tmp20118 : tmp21572;
  assign tmp21575 = s3 ? tmp21569 : tmp20210;
  assign tmp21574 = s4 ? tmp21575 : tmp20233;
  assign tmp21573 = s5 ? tmp20165 : tmp21574;
  assign tmp21570 = s6 ? tmp21571 : tmp21573;
  assign tmp21562 = s7 ? tmp21563 : tmp21570;
  assign tmp21561 = s8 ? tmp21555 : tmp21562;
  assign tmp21537 = s9 ? tmp21538 : tmp21561;
  assign tmp21577 = s8 ? tmp21555 : tmp21556;
  assign tmp21579 = s7 ? tmp21551 : tmp21570;
  assign tmp21578 = s8 ? tmp21579 : tmp21551;
  assign tmp21576 = s9 ? tmp21577 : tmp21578;
  assign tmp21536 = s10 ? tmp21537 : tmp21576;
  assign tmp21588 = s3 ? tmp20220 : tmp19965;
  assign tmp21587 = s4 ? tmp21588 : tmp20229;
  assign tmp21586 = ~(s5 ? tmp20281 : tmp21587);
  assign tmp21585 = s6 ? tmp20276 : tmp21586;
  assign tmp21584 = s7 ? tmp20252 : tmp21585;
  assign tmp21591 = s5 ? tmp20323 : tmp21553;
  assign tmp21590 = s6 ? tmp20317 : tmp21591;
  assign tmp21589 = ~(s7 ? tmp20289 : tmp21590);
  assign tmp21583 = s8 ? tmp21584 : tmp21589;
  assign tmp21593 = s7 ? tmp20289 : tmp21590;
  assign tmp21592 = ~(s8 ? tmp21593 : tmp20330);
  assign tmp21582 = s9 ? tmp21583 : tmp21592;
  assign tmp21598 = ~(s5 ? tmp20338 : tmp21587);
  assign tmp21597 = s6 ? tmp20276 : tmp21598;
  assign tmp21596 = s7 ? tmp20331 : tmp21597;
  assign tmp21595 = s8 ? tmp21596 : tmp20331;
  assign tmp21603 = s4 ? tmp20342 : tmp20229;
  assign tmp21602 = ~(s5 ? tmp20338 : tmp21603);
  assign tmp21601 = s6 ? tmp20276 : tmp21602;
  assign tmp21600 = s7 ? tmp21585 : tmp21601;
  assign tmp21605 = ~(s6 ? tmp20276 : tmp21598);
  assign tmp21604 = ~(s7 ? tmp21590 : tmp21605);
  assign tmp21599 = s8 ? tmp21600 : tmp21604;
  assign tmp21594 = s9 ? tmp21595 : tmp21599;
  assign tmp21581 = s10 ? tmp21582 : tmp21594;
  assign tmp21609 = s7 ? tmp21585 : tmp20336;
  assign tmp21608 = s8 ? tmp21609 : tmp21604;
  assign tmp21607 = s9 ? tmp21595 : tmp21608;
  assign tmp21606 = s10 ? tmp21582 : tmp21607;
  assign tmp21580 = ~(s11 ? tmp21581 : tmp21606);
  assign tmp21535 = s12 ? tmp21536 : tmp21580;
  assign tmp21377 = ~(s13 ? tmp21378 : tmp21535);
  assign tmp21135 = s14 ? tmp21136 : tmp21377;
  assign tmp21623 = ~(s1 ? tmp19651 : tmp20078);
  assign tmp21622 = s2 ? tmp20264 : tmp21623;
  assign tmp21624 = ~(s2 ? tmp19687 : tmp20663);
  assign tmp21621 = s3 ? tmp21622 : tmp21624;
  assign tmp21620 = s4 ? tmp21621 : tmp20664;
  assign tmp21619 = s5 ? tmp21620 : tmp20669;
  assign tmp21618 = s6 ? tmp20740 : tmp21619;
  assign tmp21629 = s2 ? tmp19919 : tmp20520;
  assign tmp21628 = s3 ? tmp21629 : tmp19918;
  assign tmp21627 = s4 ? tmp21628 : tmp20686;
  assign tmp21631 = s3 ? tmp20538 : tmp20545;
  assign tmp21632 = s3 ? tmp20696 : tmp20540;
  assign tmp21630 = s4 ? tmp21631 : tmp21632;
  assign tmp21626 = s5 ? tmp21627 : tmp21630;
  assign tmp21625 = s6 ? tmp20745 : tmp21626;
  assign tmp21617 = s7 ? tmp21618 : tmp21625;
  assign tmp21637 = s2 ? tmp20207 : tmp20702;
  assign tmp21636 = s3 ? tmp19916 : tmp21637;
  assign tmp21635 = s4 ? tmp21636 : tmp20656;
  assign tmp21634 = s6 ? tmp21635 : tmp20703;
  assign tmp21639 = s4 ? tmp21636 : tmp20721;
  assign tmp21642 = s3 ? tmp20733 : tmp20545;
  assign tmp21644 = s2 ? tmp20472 : tmp19635;
  assign tmp21643 = s3 ? tmp21644 : tmp20540;
  assign tmp21641 = s4 ? tmp21642 : tmp21643;
  assign tmp21640 = s5 ? tmp20724 : tmp21641;
  assign tmp21638 = s6 ? tmp21639 : tmp21640;
  assign tmp21633 = s7 ? tmp21634 : tmp21638;
  assign tmp21616 = s8 ? tmp21617 : tmp21633;
  assign tmp21651 = s2 ? tmp20264 : tmp20708;
  assign tmp21652 = s2 ? tmp19637 : tmp19919;
  assign tmp21650 = s3 ? tmp21651 : tmp21652;
  assign tmp21649 = s4 ? tmp21650 : tmp20664;
  assign tmp21648 = s5 ? tmp21649 : tmp20669;
  assign tmp21647 = s6 ? tmp20740 : tmp21648;
  assign tmp21657 = s2 ? tmp19919 : tmp20099;
  assign tmp21656 = s3 ? tmp21657 : tmp19918;
  assign tmp21655 = s4 ? tmp21656 : tmp20729;
  assign tmp21654 = s5 ? tmp21655 : tmp20749;
  assign tmp21653 = s6 ? tmp20745 : tmp21654;
  assign tmp21646 = s7 ? tmp21647 : tmp21653;
  assign tmp21645 = s8 ? tmp21633 : tmp21646;
  assign tmp21615 = s9 ? tmp21616 : tmp21645;
  assign tmp21662 = s5 ? tmp21655 : tmp21630;
  assign tmp21661 = s6 ? tmp20745 : tmp21662;
  assign tmp21660 = s7 ? tmp21647 : tmp21661;
  assign tmp21659 = s8 ? tmp21660 : tmp21647;
  assign tmp21667 = s4 ? tmp21628 : tmp20764;
  assign tmp21666 = s5 ? tmp21667 : tmp21630;
  assign tmp21665 = s6 ? tmp20745 : tmp21666;
  assign tmp21669 = s5 ? tmp21655 : tmp20769;
  assign tmp21668 = s6 ? tmp20745 : tmp21669;
  assign tmp21664 = s7 ? tmp21665 : tmp21668;
  assign tmp21670 = s7 ? tmp21638 : tmp21661;
  assign tmp21663 = s8 ? tmp21664 : tmp21670;
  assign tmp21658 = s9 ? tmp21659 : tmp21663;
  assign tmp21614 = s10 ? tmp21615 : tmp21658;
  assign tmp21674 = s7 ? tmp21625 : tmp21653;
  assign tmp21673 = s8 ? tmp21674 : tmp21670;
  assign tmp21672 = s9 ? tmp21659 : tmp21673;
  assign tmp21671 = s10 ? tmp21615 : tmp21672;
  assign tmp21613 = s11 ? tmp21614 : tmp21671;
  assign tmp21682 = s3 ? tmp20791 : tmp20123;
  assign tmp21681 = s4 ? tmp21682 : tmp20794;
  assign tmp21686 = s2 ? tmp20301 : tmp20120;
  assign tmp21685 = s3 ? tmp21686 : tmp20810;
  assign tmp21684 = s4 ? tmp21685 : tmp20812;
  assign tmp21683 = s5 ? tmp20798 : tmp21684;
  assign tmp21680 = s6 ? tmp21681 : tmp21683;
  assign tmp21688 = s4 ? tmp21682 : tmp20821;
  assign tmp21692 = s2 ? tmp20293 : tmp21460;
  assign tmp21691 = s3 ? tmp21692 : tmp20834;
  assign tmp21690 = s4 ? tmp21691 : tmp20120;
  assign tmp21689 = s5 ? tmp20824 : tmp21690;
  assign tmp21687 = s6 ? tmp21688 : tmp21689;
  assign tmp21679 = s7 ? tmp21680 : tmp21687;
  assign tmp21678 = s8 ? tmp20787 : tmp21679;
  assign tmp21677 = s9 ? tmp20787 : tmp21678;
  assign tmp21696 = s6 ? tmp21681 : tmp20797;
  assign tmp21697 = s6 ? tmp21688 : tmp20823;
  assign tmp21695 = s7 ? tmp21696 : tmp21697;
  assign tmp21694 = s8 ? tmp21695 : tmp21696;
  assign tmp21699 = s7 ? tmp20866 : tmp21687;
  assign tmp21700 = s6 ? tmp21688 : tmp20867;
  assign tmp21698 = s8 ? tmp21699 : tmp21700;
  assign tmp21693 = s9 ? tmp21694 : tmp21698;
  assign tmp21676 = s10 ? tmp21677 : tmp21693;
  assign tmp21704 = s7 ? tmp20819 : tmp21687;
  assign tmp21703 = s8 ? tmp21704 : tmp21697;
  assign tmp21702 = s9 ? tmp21694 : tmp21703;
  assign tmp21701 = s10 ? tmp21677 : tmp21702;
  assign tmp21675 = s11 ? tmp21676 : tmp21701;
  assign tmp21612 = s12 ? tmp21613 : tmp21675;
  assign tmp21611 = s13 ? tmp21612 : tmp20874;
  assign tmp21610 = ~(s14 ? tmp20362 : tmp21611);
  assign tmp21134 = s15 ? tmp21135 : tmp21610;
  assign tmp19598 = s16 ? tmp19599 : tmp21134;
  assign tmp21716 = s4 ? tmp21196 : tmp19746;
  assign tmp21715 = s5 ? tmp19713 : tmp21716;
  assign tmp21714 = s6 ? tmp19706 : tmp21715;
  assign tmp21719 = s4 ? tmp21215 : tmp19746;
  assign tmp21718 = s5 ? tmp19736 : tmp21719;
  assign tmp21717 = s6 ? tmp19706 : tmp21718;
  assign tmp21713 = s7 ? tmp21714 : tmp21717;
  assign tmp21712 = s8 ? tmp21151 : tmp21713;
  assign tmp21711 = s9 ? tmp21140 : tmp21712;
  assign tmp21724 = s5 ? tmp19753 : tmp21149;
  assign tmp21723 = s6 ? tmp19656 : tmp21724;
  assign tmp21722 = s7 ? tmp21142 : tmp21723;
  assign tmp21721 = s8 ? tmp21722 : tmp21142;
  assign tmp21726 = s7 ? tmp21261 : tmp21717;
  assign tmp21727 = s7 ? tmp21265 : tmp21723;
  assign tmp21725 = s8 ? tmp21726 : tmp21727;
  assign tmp21720 = s9 ? tmp21721 : tmp21725;
  assign tmp21710 = s10 ? tmp21711 : tmp21720;
  assign tmp21731 = s7 ? tmp21147 : tmp21717;
  assign tmp21732 = s7 ? tmp21162 : tmp21723;
  assign tmp21730 = s8 ? tmp21731 : tmp21732;
  assign tmp21729 = s9 ? tmp21721 : tmp21730;
  assign tmp21728 = s10 ? tmp21711 : tmp21729;
  assign tmp21709 = s11 ? tmp21710 : tmp21728;
  assign tmp21738 = s7 ? tmp21289 : tmp21358;
  assign tmp21737 = s8 ? tmp21309 : tmp21738;
  assign tmp21736 = s9 ? tmp21287 : tmp21737;
  assign tmp21740 = s8 ? tmp21738 : tmp21289;
  assign tmp21742 = s7 ? tmp21368 : tmp21358;
  assign tmp21741 = s8 ? tmp21358 : tmp21742;
  assign tmp21739 = s9 ? tmp21740 : tmp21741;
  assign tmp21735 = s10 ? tmp21736 : tmp21739;
  assign tmp21746 = s7 ? tmp21318 : tmp21358;
  assign tmp21745 = s8 ? tmp21302 : tmp21746;
  assign tmp21744 = s9 ? tmp21740 : tmp21745;
  assign tmp21743 = s10 ? tmp21736 : tmp21744;
  assign tmp21734 = s11 ? tmp21735 : tmp21743;
  assign tmp21733 = s12 ? tmp19769 : tmp21734;
  assign tmp21708 = s13 ? tmp21709 : tmp21733;
  assign tmp21752 = s8 ? tmp21383 : tmp19889;
  assign tmp21751 = s9 ? tmp21382 : tmp21752;
  assign tmp21755 = s7 ? tmp21419 : tmp19880;
  assign tmp21754 = s8 ? tmp19900 : tmp21755;
  assign tmp21753 = s9 ? tmp19898 : tmp21754;
  assign tmp21750 = s10 ? tmp21751 : tmp21753;
  assign tmp21759 = s7 ? tmp21402 : tmp19880;
  assign tmp21758 = s8 ? tmp19880 : tmp21759;
  assign tmp21757 = s9 ? tmp19898 : tmp21758;
  assign tmp21756 = s10 ? tmp21751 : tmp21757;
  assign tmp21749 = s11 ? tmp21750 : tmp21756;
  assign tmp21769 = s1 ? tmp19717 : tmp19614;
  assign tmp21768 = s2 ? tmp19614 : tmp21769;
  assign tmp21767 = s3 ? tmp19614 : tmp21768;
  assign tmp21771 = s2 ? tmp19614 : tmp19717;
  assign tmp21770 = s3 ? tmp21771 : tmp20020;
  assign tmp21766 = s4 ? tmp21767 : tmp21770;
  assign tmp21776 = s1 ? tmp19717 : tmp19813;
  assign tmp21777 = ~(s1 ? tmp19719 : tmp19789);
  assign tmp21775 = s2 ? tmp21776 : tmp21777;
  assign tmp21778 = ~(s2 ? tmp19719 : tmp20029);
  assign tmp21774 = s3 ? tmp21775 : tmp21778;
  assign tmp21773 = s4 ? tmp21774 : tmp20000;
  assign tmp21772 = s5 ? tmp21773 : tmp20004;
  assign tmp21765 = s6 ? tmp21766 : tmp21772;
  assign tmp21781 = s3 ? tmp21768 : tmp20020;
  assign tmp21780 = s4 ? tmp21767 : tmp21781;
  assign tmp21786 = s1 ? tmp19717 : 1;
  assign tmp21785 = s2 ? tmp21786 : tmp19716;
  assign tmp21784 = s3 ? tmp21785 : tmp19998;
  assign tmp21783 = s4 ? tmp21784 : tmp20000;
  assign tmp21782 = s5 ? tmp21783 : tmp20025;
  assign tmp21779 = s6 ? tmp21780 : tmp21782;
  assign tmp21764 = ~(s7 ? tmp21765 : tmp21779);
  assign tmp21763 = s8 ? tmp21452 : tmp21764;
  assign tmp21762 = s9 ? tmp21431 : tmp21763;
  assign tmp21792 = s4 ? tmp21449 : tmp19983;
  assign tmp21791 = s5 ? tmp21792 : tmp19962;
  assign tmp21790 = s6 ? tmp21444 : tmp21791;
  assign tmp21789 = s7 ? tmp21433 : tmp21790;
  assign tmp21788 = s8 ? tmp21789 : tmp21433;
  assign tmp21795 = ~(s6 ? tmp21780 : tmp21782);
  assign tmp21794 = s7 ? tmp21518 : tmp21795;
  assign tmp21796 = s7 ? tmp21527 : tmp21790;
  assign tmp21793 = s8 ? tmp21794 : tmp21796;
  assign tmp21787 = s9 ? tmp21788 : tmp21793;
  assign tmp21761 = s10 ? tmp21762 : tmp21787;
  assign tmp21800 = s7 ? tmp21443 : tmp21795;
  assign tmp21801 = s7 ? tmp21471 : tmp21790;
  assign tmp21799 = s8 ? tmp21800 : tmp21801;
  assign tmp21798 = s9 ? tmp21788 : tmp21799;
  assign tmp21797 = s10 ? tmp21762 : tmp21798;
  assign tmp21760 = s11 ? tmp21761 : tmp21797;
  assign tmp21748 = s12 ? tmp21749 : tmp21760;
  assign tmp21813 = s1 ? tmp20675 : tmp19806;
  assign tmp21812 = s2 ? tmp21813 : tmp20077;
  assign tmp21811 = s3 ? tmp21812 : tmp20079;
  assign tmp21810 = s4 ? tmp20066 : tmp21811;
  assign tmp21809 = s5 ? tmp21810 : tmp20082;
  assign tmp21808 = s6 ? tmp20057 : tmp21809;
  assign tmp21818 = s2 ? tmp21813 : tmp19635;
  assign tmp21817 = s3 ? tmp21818 : tmp20103;
  assign tmp21816 = s4 ? tmp20097 : tmp21817;
  assign tmp21815 = s5 ? tmp21816 : tmp20105;
  assign tmp21814 = s6 ? tmp20091 : tmp21815;
  assign tmp21807 = s7 ? tmp21808 : tmp21814;
  assign tmp21825 = s1 ? tmp20675 : tmp19720;
  assign tmp21826 = ~(s1 ? tmp19614 : tmp20078);
  assign tmp21824 = s2 ? tmp21825 : tmp21826;
  assign tmp21823 = s3 ? tmp21824 : tmp19934;
  assign tmp21822 = s4 ? tmp21463 : tmp21823;
  assign tmp21830 = s1 ? tmp19637 : tmp20085;
  assign tmp21829 = s2 ? tmp19938 : tmp21830;
  assign tmp21828 = s3 ? tmp21829 : tmp20086;
  assign tmp21832 = s2 ? tmp19846 : tmp20089;
  assign tmp21831 = s3 ? tmp21832 : tmp19945;
  assign tmp21827 = s4 ? tmp21828 : tmp21831;
  assign tmp21821 = s5 ? tmp21822 : tmp21827;
  assign tmp21820 = s6 ? tmp20057 : tmp21821;
  assign tmp21837 = s2 ? tmp21825 : tmp19635;
  assign tmp21836 = s3 ? tmp21837 : tmp19879;
  assign tmp21835 = s4 ? tmp21478 : tmp21836;
  assign tmp21834 = s5 ? tmp21835 : tmp20105;
  assign tmp21833 = s6 ? tmp20091 : tmp21834;
  assign tmp21819 = s7 ? tmp21820 : tmp21833;
  assign tmp21806 = s8 ? tmp21807 : tmp21819;
  assign tmp21846 = s0 ? tmp19614 : tmp20120;
  assign tmp21845 = s1 ? tmp21846 : tmp19806;
  assign tmp21844 = s2 ? tmp21845 : tmp20191;
  assign tmp21843 = s3 ? tmp21844 : tmp20192;
  assign tmp21842 = s4 ? tmp20185 : tmp21843;
  assign tmp21841 = s5 ? tmp21842 : tmp20194;
  assign tmp21840 = s6 ? tmp20117 : tmp21841;
  assign tmp21851 = s2 ? tmp21845 : tmp20120;
  assign tmp21850 = s3 ? tmp21851 : tmp20206;
  assign tmp21849 = s4 ? tmp20202 : tmp21850;
  assign tmp21848 = s5 ? tmp21849 : tmp20208;
  assign tmp21847 = s6 ? tmp20160 : tmp21848;
  assign tmp21839 = s7 ? tmp21840 : tmp21847;
  assign tmp21838 = s8 ? tmp21819 : tmp21839;
  assign tmp21805 = s9 ? tmp21806 : tmp21838;
  assign tmp21856 = s5 ? tmp21816 : tmp20218;
  assign tmp21855 = s6 ? tmp20091 : tmp21856;
  assign tmp21854 = s7 ? tmp21808 : tmp21855;
  assign tmp21853 = s8 ? tmp21854 : tmp21808;
  assign tmp21860 = s5 ? tmp21816 : tmp20228;
  assign tmp21859 = s6 ? tmp20091 : tmp21860;
  assign tmp21862 = s5 ? tmp21849 : tmp20232;
  assign tmp21861 = s6 ? tmp20160 : tmp21862;
  assign tmp21858 = s7 ? tmp21859 : tmp21861;
  assign tmp21865 = s5 ? tmp21835 : tmp20228;
  assign tmp21864 = s6 ? tmp20091 : tmp21865;
  assign tmp21867 = s5 ? tmp21816 : tmp20241;
  assign tmp21866 = s6 ? tmp20091 : tmp21867;
  assign tmp21863 = s7 ? tmp21864 : tmp21866;
  assign tmp21857 = s8 ? tmp21858 : tmp21863;
  assign tmp21852 = s9 ? tmp21853 : tmp21857;
  assign tmp21804 = s10 ? tmp21805 : tmp21852;
  assign tmp21871 = s7 ? tmp21814 : tmp21847;
  assign tmp21872 = s7 ? tmp21833 : tmp21855;
  assign tmp21870 = s8 ? tmp21871 : tmp21872;
  assign tmp21869 = s9 ? tmp21853 : tmp21870;
  assign tmp21868 = s10 ? tmp21805 : tmp21869;
  assign tmp21803 = s11 ? tmp21804 : tmp21868;
  assign tmp21802 = s12 ? tmp21803 : tmp20247;
  assign tmp21747 = ~(s13 ? tmp21748 : tmp21802);
  assign tmp21707 = s14 ? tmp21708 : tmp21747;
  assign tmp21879 = s8 ? tmp20787 : tmp20853;
  assign tmp21878 = s9 ? tmp20787 : tmp21879;
  assign tmp21882 = s7 ? tmp20866 : tmp20860;
  assign tmp21881 = s8 ? tmp20865 : tmp21882;
  assign tmp21880 = s9 ? tmp20858 : tmp21881;
  assign tmp21877 = s10 ? tmp21878 : tmp21880;
  assign tmp21886 = s7 ? tmp20819 : tmp20860;
  assign tmp21885 = s8 ? tmp20873 : tmp21886;
  assign tmp21884 = s9 ? tmp20858 : tmp21885;
  assign tmp21883 = s10 ? tmp21878 : tmp21884;
  assign tmp21876 = s11 ? tmp21877 : tmp21883;
  assign tmp21875 = s12 ? tmp20646 : tmp21876;
  assign tmp21874 = s13 ? tmp21875 : tmp20874;
  assign tmp21873 = ~(s14 ? tmp20362 : tmp21874);
  assign tmp21706 = s15 ? tmp21707 : tmp21873;
  assign tmp21901 = s1 ? tmp21846 : tmp19720;
  assign tmp21900 = s2 ? tmp21901 : tmp20145;
  assign tmp21899 = s3 ? tmp21900 : tmp20147;
  assign tmp21898 = s4 ? tmp20136 : tmp21899;
  assign tmp21897 = s5 ? tmp21898 : tmp20149;
  assign tmp21896 = s6 ? tmp20117 : tmp21897;
  assign tmp21906 = s2 ? tmp21901 : tmp20120;
  assign tmp21905 = s3 ? tmp21906 : tmp20172;
  assign tmp21904 = s4 ? tmp20166 : tmp21905;
  assign tmp21908 = s3 ? tmp20314 : tmp20210;
  assign tmp21911 = s1 ? tmp20120 : tmp20158;
  assign tmp21910 = s2 ? 1 : tmp21911;
  assign tmp21909 = s3 ? tmp21910 : tmp19635;
  assign tmp21907 = s4 ? tmp21908 : tmp21909;
  assign tmp21903 = s5 ? tmp21904 : tmp21907;
  assign tmp21902 = s6 ? tmp20160 : tmp21903;
  assign tmp21895 = s7 ? tmp21896 : tmp21902;
  assign tmp21894 = s8 ? tmp21819 : tmp21895;
  assign tmp21893 = s9 ? tmp21806 : tmp21894;
  assign tmp21913 = s8 ? tmp21819 : tmp21820;
  assign tmp21918 = s4 ? tmp21908 : tmp20233;
  assign tmp21917 = s5 ? tmp21904 : tmp21918;
  assign tmp21916 = s6 ? tmp20160 : tmp21917;
  assign tmp21915 = s7 ? tmp21859 : tmp21916;
  assign tmp21914 = s8 ? tmp21915 : tmp21864;
  assign tmp21912 = s9 ? tmp21913 : tmp21914;
  assign tmp21892 = s10 ? tmp21893 : tmp21912;
  assign tmp21922 = s7 ? tmp21814 : tmp21902;
  assign tmp21921 = s8 ? tmp21922 : tmp21833;
  assign tmp21920 = s9 ? tmp21913 : tmp21921;
  assign tmp21919 = s10 ? tmp21893 : tmp21920;
  assign tmp21891 = s11 ? tmp21892 : tmp21919;
  assign tmp21890 = s12 ? tmp21891 : tmp20247;
  assign tmp21889 = ~(s13 ? tmp21378 : tmp21890);
  assign tmp21888 = s14 ? tmp21136 : tmp21889;
  assign tmp21925 = s12 ? tmp20646 : tmp21675;
  assign tmp21924 = s13 ? tmp21925 : tmp20874;
  assign tmp21923 = ~(s14 ? tmp20362 : tmp21924);
  assign tmp21887 = s15 ? tmp21888 : tmp21923;
  assign tmp21705 = s16 ? tmp21706 : tmp21887;
  assign tmp19597 = ~(s17 ? tmp19598 : tmp21705);
  assign s13n = tmp19597;

  assign tmp21941 = ~(l2 ? 1 : 0);
  assign tmp21940 = l1 ? 1 : tmp21941;
  assign tmp21943 = l1 ? 1 : 0;
  assign tmp21942 = s0 ? tmp21943 : tmp21940;
  assign tmp21939 = s1 ? tmp21940 : tmp21942;
  assign tmp21946 = s0 ? tmp21940 : tmp21943;
  assign tmp21945 = s1 ? tmp21946 : tmp21940;
  assign tmp21944 = s2 ? tmp21940 : tmp21945;
  assign tmp21938 = s3 ? tmp21939 : tmp21944;
  assign tmp21950 = s0 ? tmp21940 : 1;
  assign tmp21951 = s0 ? tmp21943 : 1;
  assign tmp21949 = s1 ? tmp21950 : tmp21951;
  assign tmp21948 = s2 ? tmp21945 : tmp21949;
  assign tmp21953 = s1 ? tmp21943 : 1;
  assign tmp21955 = s0 ? tmp21940 : tmp21941;
  assign tmp21956 = s0 ? 1 : tmp21940;
  assign tmp21954 = s1 ? tmp21955 : tmp21956;
  assign tmp21952 = s2 ? tmp21953 : tmp21954;
  assign tmp21947 = s3 ? tmp21948 : tmp21952;
  assign tmp21937 = s4 ? tmp21938 : tmp21947;
  assign tmp21961 = s1 ? tmp21946 : tmp21942;
  assign tmp21964 = l2 ? 1 : 0;
  assign tmp21963 = ~(s0 ? tmp21964 : 1);
  assign tmp21962 = s1 ? tmp21942 : tmp21963;
  assign tmp21960 = s2 ? tmp21961 : tmp21962;
  assign tmp21966 = s0 ? 1 : tmp21964;
  assign tmp21967 = ~(s1 ? 1 : tmp21950);
  assign tmp21965 = ~(s2 ? tmp21966 : tmp21967);
  assign tmp21959 = s3 ? tmp21960 : tmp21965;
  assign tmp21970 = s1 ? tmp21956 : tmp21951;
  assign tmp21971 = s1 ? tmp21951 : tmp21946;
  assign tmp21969 = s2 ? tmp21970 : tmp21971;
  assign tmp21973 = s1 ? tmp21964 : 0;
  assign tmp21972 = ~(s2 ? tmp21973 : 0);
  assign tmp21968 = s3 ? tmp21969 : tmp21972;
  assign tmp21958 = s4 ? tmp21959 : tmp21968;
  assign tmp21978 = s0 ? tmp21964 : 0;
  assign tmp21977 = s1 ? tmp21978 : 0;
  assign tmp21980 = s0 ? 1 : tmp21941;
  assign tmp21979 = ~(s1 ? tmp21980 : tmp21941);
  assign tmp21976 = s2 ? tmp21977 : tmp21979;
  assign tmp21975 = s3 ? tmp21976 : 0;
  assign tmp21983 = s1 ? tmp21980 : tmp21941;
  assign tmp21982 = s2 ? 1 : tmp21983;
  assign tmp21981 = ~(s3 ? tmp21982 : 1);
  assign tmp21974 = ~(s4 ? tmp21975 : tmp21981);
  assign tmp21957 = s5 ? tmp21958 : tmp21974;
  assign tmp21936 = s6 ? tmp21937 : tmp21957;
  assign tmp21988 = s1 ? tmp21950 : tmp21943;
  assign tmp21987 = s2 ? tmp21945 : tmp21988;
  assign tmp21986 = s3 ? tmp21987 : tmp21952;
  assign tmp21985 = s4 ? tmp21938 : tmp21986;
  assign tmp21993 = s1 ? tmp21940 : tmp21963;
  assign tmp21992 = s2 ? tmp21945 : tmp21993;
  assign tmp21994 = ~(s2 ? tmp21964 : tmp21967);
  assign tmp21991 = s3 ? tmp21992 : tmp21994;
  assign tmp21997 = s1 ? tmp21943 : tmp21946;
  assign tmp21996 = s2 ? tmp21970 : tmp21997;
  assign tmp21995 = s3 ? tmp21996 : tmp21972;
  assign tmp21990 = s4 ? tmp21991 : tmp21995;
  assign tmp22000 = s2 ? tmp21977 : tmp21973;
  assign tmp21999 = s3 ? tmp22000 : 0;
  assign tmp22002 = s2 ? 1 : tmp21941;
  assign tmp22001 = ~(s3 ? tmp22002 : 1);
  assign tmp21998 = ~(s4 ? tmp21999 : tmp22001);
  assign tmp21989 = s5 ? tmp21990 : tmp21998;
  assign tmp21984 = s6 ? tmp21985 : tmp21989;
  assign tmp21935 = s7 ? tmp21936 : tmp21984;
  assign tmp22008 = s1 ? tmp21940 : tmp21956;
  assign tmp22007 = s2 ? tmp21953 : tmp22008;
  assign tmp22006 = s3 ? tmp21948 : tmp22007;
  assign tmp22005 = s4 ? tmp21938 : tmp22006;
  assign tmp22013 = s1 ? tmp21942 : tmp21946;
  assign tmp22012 = s2 ? tmp21961 : tmp22013;
  assign tmp22016 = s0 ? tmp21943 : tmp21941;
  assign tmp22015 = s1 ? tmp21942 : tmp22016;
  assign tmp22017 = s1 ? 1 : tmp21950;
  assign tmp22014 = s2 ? tmp22015 : tmp22017;
  assign tmp22011 = s3 ? tmp22012 : tmp22014;
  assign tmp22019 = ~(s2 ? tmp21977 : 0);
  assign tmp22018 = s3 ? tmp21969 : tmp22019;
  assign tmp22010 = s4 ? tmp22011 : tmp22018;
  assign tmp22009 = s5 ? tmp22010 : tmp21974;
  assign tmp22004 = s6 ? tmp22005 : tmp22009;
  assign tmp22022 = s3 ? tmp21987 : tmp22007;
  assign tmp22021 = s4 ? tmp21938 : tmp22022;
  assign tmp22027 = s1 ? tmp21940 : tmp21946;
  assign tmp22026 = s2 ? tmp21945 : tmp22027;
  assign tmp22029 = s1 ? tmp21940 : tmp21941;
  assign tmp22028 = s2 ? tmp22029 : tmp22017;
  assign tmp22025 = s3 ? tmp22026 : tmp22028;
  assign tmp22031 = s2 ? tmp21970 : tmp21940;
  assign tmp22030 = s3 ? tmp22031 : tmp22019;
  assign tmp22024 = s4 ? tmp22025 : tmp22030;
  assign tmp22023 = s5 ? tmp22024 : tmp21998;
  assign tmp22020 = s6 ? tmp22021 : tmp22023;
  assign tmp22003 = s7 ? tmp22004 : tmp22020;
  assign tmp21934 = s8 ? tmp21935 : tmp22003;
  assign tmp22037 = s2 ? tmp21943 : tmp21951;
  assign tmp22040 = s0 ? 1 : tmp21943;
  assign tmp22039 = s1 ? tmp21943 : tmp22040;
  assign tmp22038 = s2 ? tmp21953 : tmp22039;
  assign tmp22036 = s3 ? tmp22037 : tmp22038;
  assign tmp22035 = s4 ? tmp21943 : tmp22036;
  assign tmp22046 = s0 ? tmp21943 : 0;
  assign tmp22045 = s1 ? tmp21943 : tmp22046;
  assign tmp22044 = s2 ? tmp21943 : tmp22045;
  assign tmp22049 = ~(l1 ? 1 : 0);
  assign tmp22048 = s0 ? 1 : tmp22049;
  assign tmp22050 = ~(s1 ? 1 : tmp21951);
  assign tmp22047 = ~(s2 ? tmp22048 : tmp22050);
  assign tmp22043 = s3 ? tmp22044 : tmp22047;
  assign tmp22053 = s1 ? tmp22040 : tmp21951;
  assign tmp22054 = s1 ? tmp21951 : tmp21943;
  assign tmp22052 = s2 ? tmp22053 : tmp22054;
  assign tmp22055 = s2 ? tmp21943 : 1;
  assign tmp22051 = s3 ? tmp22052 : tmp22055;
  assign tmp22042 = s4 ? tmp22043 : tmp22051;
  assign tmp22059 = s1 ? tmp21951 : 1;
  assign tmp22060 = s1 ? tmp22040 : tmp21943;
  assign tmp22058 = s2 ? tmp22059 : tmp22060;
  assign tmp22057 = s3 ? tmp22058 : 1;
  assign tmp22062 = s2 ? 1 : tmp22060;
  assign tmp22061 = s3 ? tmp22062 : 1;
  assign tmp22056 = s4 ? tmp22057 : tmp22061;
  assign tmp22041 = s5 ? tmp22042 : tmp22056;
  assign tmp22034 = s6 ? tmp22035 : tmp22041;
  assign tmp22066 = s2 ? tmp21943 : tmp22054;
  assign tmp22065 = s3 ? tmp22066 : tmp22038;
  assign tmp22064 = s4 ? tmp21943 : tmp22065;
  assign tmp22071 = s1 ? 1 : tmp21951;
  assign tmp22070 = s2 ? tmp21943 : tmp22071;
  assign tmp22069 = s3 ? tmp22044 : tmp22070;
  assign tmp22073 = s2 ? tmp22053 : tmp21943;
  assign tmp22074 = s2 ? tmp21953 : 1;
  assign tmp22072 = s3 ? tmp22073 : tmp22074;
  assign tmp22068 = s4 ? tmp22069 : tmp22072;
  assign tmp22077 = s2 ? tmp22059 : tmp21953;
  assign tmp22076 = s3 ? tmp22077 : 1;
  assign tmp22079 = s2 ? 1 : tmp21943;
  assign tmp22078 = s3 ? tmp22079 : 1;
  assign tmp22075 = s4 ? tmp22076 : tmp22078;
  assign tmp22067 = s5 ? tmp22068 : tmp22075;
  assign tmp22063 = s6 ? tmp22064 : tmp22067;
  assign tmp22033 = s7 ? tmp22034 : tmp22063;
  assign tmp22032 = s8 ? tmp22003 : tmp22033;
  assign tmp21933 = s9 ? tmp21934 : tmp22032;
  assign tmp22086 = s3 ? tmp22031 : tmp21972;
  assign tmp22085 = s4 ? tmp21991 : tmp22086;
  assign tmp22084 = s5 ? tmp22085 : tmp21998;
  assign tmp22083 = s6 ? tmp21985 : tmp22084;
  assign tmp22082 = s7 ? tmp21936 : tmp22083;
  assign tmp22081 = s8 ? tmp22082 : tmp21936;
  assign tmp22094 = s1 ? tmp21943 : tmp21940;
  assign tmp22093 = s2 ? tmp21970 : tmp22094;
  assign tmp22092 = s3 ? tmp22093 : tmp21972;
  assign tmp22091 = s4 ? tmp21991 : tmp22092;
  assign tmp22090 = s5 ? tmp22091 : tmp21998;
  assign tmp22089 = s6 ? tmp21985 : tmp22090;
  assign tmp22088 = s7 ? tmp22089 : tmp22063;
  assign tmp22095 = s7 ? tmp22020 : tmp22083;
  assign tmp22087 = s8 ? tmp22088 : tmp22095;
  assign tmp22080 = s9 ? tmp22081 : tmp22087;
  assign tmp21932 = s10 ? tmp21933 : tmp22080;
  assign tmp22099 = s7 ? tmp21984 : tmp22063;
  assign tmp22098 = s8 ? tmp22099 : tmp22095;
  assign tmp22097 = s9 ? tmp22081 : tmp22098;
  assign tmp22096 = s10 ? tmp21933 : tmp22097;
  assign tmp21931 = s11 ? tmp21932 : tmp22096;
  assign tmp22111 = ~(s0 ? 1 : tmp22049);
  assign tmp22110 = s1 ? tmp22046 : tmp22111;
  assign tmp22109 = s2 ? tmp22045 : tmp22110;
  assign tmp22108 = s3 ? tmp21943 : tmp22109;
  assign tmp22107 = s4 ? tmp21943 : tmp22108;
  assign tmp22116 = s1 ? tmp21943 : 0;
  assign tmp22115 = s2 ? tmp21943 : tmp22116;
  assign tmp22119 = ~(s0 ? tmp21943 : 0);
  assign tmp22118 = s1 ? 1 : tmp22119;
  assign tmp22117 = ~(s2 ? 1 : tmp22118);
  assign tmp22114 = s3 ? tmp22115 : tmp22117;
  assign tmp22122 = s1 ? tmp22048 : tmp22119;
  assign tmp22123 = ~(s1 ? tmp22046 : tmp21943);
  assign tmp22121 = s2 ? tmp22122 : tmp22123;
  assign tmp22120 = ~(s3 ? tmp22121 : 1);
  assign tmp22113 = s4 ? tmp22114 : tmp22120;
  assign tmp22112 = s5 ? tmp22113 : 0;
  assign tmp22106 = s6 ? tmp22107 : tmp22112;
  assign tmp22128 = s2 ? tmp22122 : tmp22049;
  assign tmp22127 = ~(s3 ? tmp22128 : 1);
  assign tmp22126 = s4 ? tmp22114 : tmp22127;
  assign tmp22125 = s5 ? tmp22126 : 0;
  assign tmp22124 = s6 ? tmp22107 : tmp22125;
  assign tmp22105 = s7 ? tmp22106 : tmp22124;
  assign tmp22134 = s1 ? tmp21943 : tmp22111;
  assign tmp22133 = s2 ? tmp22045 : tmp22134;
  assign tmp22132 = s3 ? tmp21943 : tmp22133;
  assign tmp22131 = s4 ? tmp21943 : tmp22132;
  assign tmp22140 = ~(s0 ? tmp21943 : 1);
  assign tmp22139 = ~(s1 ? 1 : tmp22140);
  assign tmp22138 = s2 ? tmp22045 : tmp22139;
  assign tmp22137 = s3 ? tmp21943 : tmp22138;
  assign tmp22143 = s1 ? tmp22048 : tmp22140;
  assign tmp22144 = ~(s1 ? tmp21951 : tmp21943);
  assign tmp22142 = s2 ? tmp22143 : tmp22144;
  assign tmp22147 = s0 ? 1 : 0;
  assign tmp22148 = ~(s0 ? 1 : 0);
  assign tmp22146 = s1 ? tmp22147 : tmp22148;
  assign tmp22145 = s2 ? tmp22146 : 1;
  assign tmp22141 = ~(s3 ? tmp22142 : tmp22145);
  assign tmp22136 = s4 ? tmp22137 : tmp22141;
  assign tmp22135 = s5 ? tmp22136 : 0;
  assign tmp22130 = s6 ? tmp22131 : tmp22135;
  assign tmp22152 = s2 ? tmp22116 : tmp22134;
  assign tmp22151 = s3 ? tmp21943 : tmp22152;
  assign tmp22150 = s4 ? tmp21943 : tmp22151;
  assign tmp22156 = s2 ? tmp22116 : tmp22139;
  assign tmp22155 = s3 ? tmp21943 : tmp22156;
  assign tmp22158 = s2 ? tmp22143 : tmp22049;
  assign tmp22160 = s1 ? tmp22147 : 1;
  assign tmp22159 = s2 ? tmp22160 : 1;
  assign tmp22157 = ~(s3 ? tmp22158 : tmp22159);
  assign tmp22154 = s4 ? tmp22155 : tmp22157;
  assign tmp22153 = s5 ? tmp22154 : 0;
  assign tmp22149 = s6 ? tmp22150 : tmp22153;
  assign tmp22129 = s7 ? tmp22130 : tmp22149;
  assign tmp22104 = s8 ? tmp22105 : tmp22129;
  assign tmp22168 = s1 ? tmp22048 : tmp22049;
  assign tmp22167 = s2 ? tmp22168 : tmp22049;
  assign tmp22166 = ~(s3 ? tmp22167 : 1);
  assign tmp22165 = s4 ? tmp22114 : tmp22166;
  assign tmp22164 = s5 ? tmp22165 : 0;
  assign tmp22163 = s6 ? tmp22107 : tmp22164;
  assign tmp22172 = s2 ? tmp22116 : tmp22110;
  assign tmp22171 = s3 ? tmp21943 : tmp22172;
  assign tmp22170 = s4 ? tmp21943 : tmp22171;
  assign tmp22169 = s6 ? tmp22170 : tmp22164;
  assign tmp22162 = s7 ? tmp22163 : tmp22169;
  assign tmp22161 = s8 ? tmp22129 : tmp22162;
  assign tmp22103 = s9 ? tmp22104 : tmp22161;
  assign tmp22174 = s8 ? tmp22162 : tmp22163;
  assign tmp22177 = s6 ? tmp22170 : tmp22125;
  assign tmp22176 = s7 ? tmp22177 : tmp22169;
  assign tmp22178 = s7 ? tmp22149 : tmp22169;
  assign tmp22175 = s8 ? tmp22176 : tmp22178;
  assign tmp22173 = s9 ? tmp22174 : tmp22175;
  assign tmp22102 = s10 ? tmp22103 : tmp22173;
  assign tmp22182 = s7 ? tmp22124 : tmp22169;
  assign tmp22181 = s8 ? tmp22182 : tmp22178;
  assign tmp22180 = s9 ? tmp22174 : tmp22181;
  assign tmp22179 = s10 ? tmp22103 : tmp22180;
  assign tmp22101 = s11 ? tmp22102 : tmp22179;
  assign tmp22193 = s0 ? tmp21943 : tmp22049;
  assign tmp22192 = s1 ? tmp21943 : tmp22193;
  assign tmp22191 = s2 ? tmp22192 : tmp22110;
  assign tmp22190 = s3 ? tmp21943 : tmp22191;
  assign tmp22189 = s4 ? tmp21943 : tmp22190;
  assign tmp22198 = s1 ? 1 : tmp22048;
  assign tmp22200 = ~(s0 ? 1 : tmp21943);
  assign tmp22199 = s1 ? 1 : tmp22200;
  assign tmp22197 = ~(s2 ? tmp22198 : tmp22199);
  assign tmp22196 = s3 ? tmp22115 : tmp22197;
  assign tmp22203 = s1 ? tmp22046 : tmp22200;
  assign tmp22204 = ~(s1 ? tmp22040 : 1);
  assign tmp22202 = s2 ? tmp22203 : tmp22204;
  assign tmp22206 = s1 ? tmp21943 : tmp21951;
  assign tmp22205 = ~(s2 ? tmp22206 : tmp22050);
  assign tmp22201 = ~(s3 ? tmp22202 : tmp22205);
  assign tmp22195 = s4 ? tmp22196 : tmp22201;
  assign tmp22210 = s1 ? tmp22046 : 0;
  assign tmp22211 = ~(s1 ? tmp22048 : tmp22200);
  assign tmp22209 = s2 ? tmp22210 : tmp22211;
  assign tmp22213 = s1 ? 1 : tmp22147;
  assign tmp22214 = ~(s1 ? tmp22040 : tmp22046);
  assign tmp22212 = s2 ? tmp22213 : tmp22214;
  assign tmp22208 = s3 ? tmp22209 : tmp22212;
  assign tmp22217 = ~(s1 ? tmp22048 : tmp22140);
  assign tmp22216 = s2 ? tmp22143 : tmp22217;
  assign tmp22219 = s1 ? tmp22040 : tmp22147;
  assign tmp22218 = ~(s2 ? tmp22219 : tmp22110);
  assign tmp22215 = s3 ? tmp22216 : tmp22218;
  assign tmp22207 = s4 ? tmp22208 : tmp22215;
  assign tmp22194 = s5 ? tmp22195 : tmp22207;
  assign tmp22188 = s6 ? tmp22189 : tmp22194;
  assign tmp22225 = s1 ? 1 : 0;
  assign tmp22224 = s2 ? tmp21943 : tmp22225;
  assign tmp22227 = s1 ? 1 : tmp22049;
  assign tmp22226 = ~(s2 ? tmp22227 : tmp22199);
  assign tmp22223 = s3 ? tmp22224 : tmp22226;
  assign tmp22229 = s2 ? tmp22203 : 0;
  assign tmp22231 = ~(s1 ? 1 : tmp21943);
  assign tmp22230 = ~(s2 ? tmp21953 : tmp22231);
  assign tmp22228 = ~(s3 ? tmp22229 : tmp22230);
  assign tmp22222 = s4 ? tmp22223 : tmp22228;
  assign tmp22234 = s2 ? tmp22210 : tmp21953;
  assign tmp22236 = ~(s1 ? tmp21943 : 0);
  assign tmp22235 = s2 ? tmp22225 : tmp22236;
  assign tmp22233 = s3 ? tmp22234 : tmp22235;
  assign tmp22238 = s2 ? tmp21953 : tmp22049;
  assign tmp22237 = ~(s3 ? tmp22238 : tmp22116);
  assign tmp22232 = s4 ? tmp22233 : tmp22237;
  assign tmp22221 = s5 ? tmp22222 : tmp22232;
  assign tmp22220 = s6 ? tmp22189 : tmp22221;
  assign tmp22187 = s7 ? tmp22188 : tmp22220;
  assign tmp22243 = s2 ? tmp22192 : tmp22134;
  assign tmp22242 = s3 ? tmp21943 : tmp22243;
  assign tmp22241 = s4 ? tmp21943 : tmp22242;
  assign tmp22248 = ~(s1 ? 1 : 0);
  assign tmp22247 = s2 ? tmp22206 : tmp22248;
  assign tmp22246 = s3 ? tmp22066 : tmp22247;
  assign tmp22250 = s2 ? tmp22210 : 0;
  assign tmp22251 = ~(s2 ? 1 : tmp22050);
  assign tmp22249 = ~(s3 ? tmp22250 : tmp22251);
  assign tmp22245 = s4 ? tmp22246 : tmp22249;
  assign tmp22255 = s1 ? tmp22147 : 0;
  assign tmp22256 = ~(s1 ? tmp22147 : 0);
  assign tmp22254 = s2 ? tmp22255 : tmp22256;
  assign tmp22253 = s3 ? tmp22254 : tmp22212;
  assign tmp22258 = s2 ? tmp22143 : tmp22256;
  assign tmp22257 = s3 ? tmp22258 : tmp22218;
  assign tmp22252 = s4 ? tmp22253 : tmp22257;
  assign tmp22244 = s5 ? tmp22245 : tmp22252;
  assign tmp22240 = s6 ? tmp22241 : tmp22244;
  assign tmp22262 = s2 ? tmp21943 : tmp21953;
  assign tmp22264 = s1 ? tmp21943 : tmp22049;
  assign tmp22263 = s2 ? tmp22264 : tmp22134;
  assign tmp22261 = s3 ? tmp22262 : tmp22263;
  assign tmp22260 = s4 ? tmp21943 : tmp22261;
  assign tmp22269 = s1 ? 1 : tmp21943;
  assign tmp22268 = s2 ? tmp21943 : tmp22269;
  assign tmp22270 = s2 ? tmp21953 : tmp22248;
  assign tmp22267 = s3 ? tmp22268 : tmp22270;
  assign tmp22272 = ~(s2 ? 1 : tmp22231);
  assign tmp22271 = ~(s3 ? tmp22250 : tmp22272);
  assign tmp22266 = s4 ? tmp22267 : tmp22271;
  assign tmp22275 = s2 ? tmp22255 : 1;
  assign tmp22274 = s3 ? tmp22275 : tmp22235;
  assign tmp22277 = s2 ? tmp21953 : 0;
  assign tmp22276 = ~(s3 ? tmp22277 : tmp22116);
  assign tmp22273 = s4 ? tmp22274 : tmp22276;
  assign tmp22265 = s5 ? tmp22266 : tmp22273;
  assign tmp22259 = s6 ? tmp22260 : tmp22265;
  assign tmp22239 = s7 ? tmp22240 : tmp22259;
  assign tmp22186 = s8 ? tmp22187 : tmp22239;
  assign tmp22284 = ~(s2 ? tmp22213 : tmp22225);
  assign tmp22283 = s3 ? tmp22115 : tmp22284;
  assign tmp22282 = s4 ? tmp22283 : tmp22249;
  assign tmp22281 = s5 ? tmp22282 : tmp22252;
  assign tmp22280 = s6 ? tmp22189 : tmp22281;
  assign tmp22288 = s2 ? tmp22264 : tmp22110;
  assign tmp22287 = s3 ? tmp22262 : tmp22288;
  assign tmp22286 = s4 ? tmp21943 : tmp22287;
  assign tmp22291 = s3 ? tmp22224 : tmp22248;
  assign tmp22290 = s4 ? tmp22291 : tmp22271;
  assign tmp22289 = s5 ? tmp22290 : tmp22273;
  assign tmp22285 = s6 ? tmp22286 : tmp22289;
  assign tmp22279 = s7 ? tmp22280 : tmp22285;
  assign tmp22278 = s8 ? tmp22239 : tmp22279;
  assign tmp22185 = s9 ? tmp22186 : tmp22278;
  assign tmp22293 = s8 ? tmp22279 : tmp22280;
  assign tmp22298 = s3 ? tmp21943 : tmp22288;
  assign tmp22297 = s4 ? tmp21943 : tmp22298;
  assign tmp22296 = s6 ? tmp22297 : tmp22221;
  assign tmp22295 = s7 ? tmp22296 : tmp22285;
  assign tmp22299 = s7 ? tmp22259 : tmp22285;
  assign tmp22294 = s8 ? tmp22295 : tmp22299;
  assign tmp22292 = s9 ? tmp22293 : tmp22294;
  assign tmp22184 = s10 ? tmp22185 : tmp22292;
  assign tmp22303 = s7 ? tmp22220 : tmp22285;
  assign tmp22302 = s8 ? tmp22303 : tmp22299;
  assign tmp22301 = s9 ? tmp22293 : tmp22302;
  assign tmp22300 = s10 ? tmp22185 : tmp22301;
  assign tmp22183 = s11 ? tmp22184 : tmp22300;
  assign tmp22100 = s12 ? tmp22101 : tmp22183;
  assign tmp21930 = s13 ? tmp21931 : tmp22100;
  assign tmp22315 = ~(s0 ? tmp21943 : tmp21941);
  assign tmp22314 = s1 ? tmp21964 : tmp22315;
  assign tmp22317 = s1 ? tmp21978 : tmp21964;
  assign tmp22316 = s2 ? tmp21964 : tmp22317;
  assign tmp22313 = s3 ? tmp22314 : tmp22316;
  assign tmp22320 = s1 ? tmp21978 : tmp22140;
  assign tmp22319 = s2 ? tmp22317 : tmp22320;
  assign tmp22322 = s1 ? tmp21943 : tmp22147;
  assign tmp22323 = ~(s1 ? tmp21964 : tmp21966);
  assign tmp22321 = ~(s2 ? tmp22322 : tmp22323);
  assign tmp22318 = s3 ? tmp22319 : tmp22321;
  assign tmp22312 = s4 ? tmp22313 : tmp22318;
  assign tmp22328 = s1 ? 1 : tmp21964;
  assign tmp22327 = s2 ? tmp21964 : tmp22328;
  assign tmp22326 = s3 ? tmp21976 : tmp22327;
  assign tmp22331 = s1 ? tmp21966 : tmp22049;
  assign tmp22333 = ~(s0 ? tmp21964 : 0);
  assign tmp22332 = ~(s1 ? tmp21943 : tmp22333);
  assign tmp22330 = s2 ? tmp22331 : tmp22332;
  assign tmp22334 = s2 ? tmp22314 : 1;
  assign tmp22329 = s3 ? tmp22330 : tmp22334;
  assign tmp22325 = s4 ? tmp22326 : tmp22329;
  assign tmp22339 = s0 ? tmp21964 : 1;
  assign tmp22338 = s1 ? tmp22339 : 1;
  assign tmp22337 = s2 ? tmp22338 : tmp22255;
  assign tmp22341 = ~(s1 ? 1 : tmp21966);
  assign tmp22340 = ~(s2 ? tmp22255 : tmp22341);
  assign tmp22336 = s3 ? tmp22337 : tmp22340;
  assign tmp22344 = s1 ? tmp21966 : 0;
  assign tmp22343 = s2 ? tmp22338 : tmp22344;
  assign tmp22346 = s1 ? 1 : tmp21966;
  assign tmp22347 = s1 ? tmp21966 : 1;
  assign tmp22345 = s2 ? tmp22346 : tmp22347;
  assign tmp22342 = s3 ? tmp22343 : tmp22345;
  assign tmp22335 = s4 ? tmp22336 : tmp22342;
  assign tmp22324 = s5 ? tmp22325 : tmp22335;
  assign tmp22311 = s6 ? tmp22312 : tmp22324;
  assign tmp22352 = s1 ? tmp21978 : tmp22049;
  assign tmp22351 = s2 ? tmp22317 : tmp22352;
  assign tmp22353 = ~(s2 ? tmp22116 : tmp22323);
  assign tmp22350 = s3 ? tmp22351 : tmp22353;
  assign tmp22349 = s4 ? tmp22313 : tmp22350;
  assign tmp22357 = s2 ? tmp21977 : tmp21964;
  assign tmp22356 = s3 ? tmp22357 : tmp22327;
  assign tmp22360 = ~(s1 ? tmp21943 : tmp21941);
  assign tmp22359 = s2 ? tmp22331 : tmp22360;
  assign tmp22358 = s3 ? tmp22359 : tmp22334;
  assign tmp22355 = s4 ? tmp22356 : tmp22358;
  assign tmp22363 = s2 ? tmp22338 : 0;
  assign tmp22364 = s2 ? 1 : tmp22328;
  assign tmp22362 = s3 ? tmp22363 : tmp22364;
  assign tmp22366 = s2 ? 1 : tmp21964;
  assign tmp22365 = s3 ? tmp22366 : tmp22328;
  assign tmp22361 = s4 ? tmp22362 : tmp22365;
  assign tmp22354 = s5 ? tmp22355 : tmp22361;
  assign tmp22348 = s6 ? tmp22349 : tmp22354;
  assign tmp22310 = s7 ? tmp22311 : tmp22348;
  assign tmp22373 = ~(s1 ? tmp21980 : tmp22333);
  assign tmp22372 = s2 ? tmp21977 : tmp22373;
  assign tmp22375 = ~(s1 ? 1 : tmp21964);
  assign tmp22374 = ~(s2 ? tmp21980 : tmp22375);
  assign tmp22371 = s3 ? tmp22372 : tmp22374;
  assign tmp22370 = s4 ? tmp22371 : tmp22329;
  assign tmp22369 = s5 ? tmp22370 : tmp22335;
  assign tmp22368 = s6 ? tmp22312 : tmp22369;
  assign tmp22381 = s1 ? tmp21964 : tmp21978;
  assign tmp22380 = s2 ? tmp21977 : tmp22381;
  assign tmp22379 = s3 ? tmp22380 : tmp22327;
  assign tmp22383 = s2 ? tmp22331 : tmp21964;
  assign tmp22384 = s2 ? tmp21964 : 1;
  assign tmp22382 = s3 ? tmp22383 : tmp22384;
  assign tmp22378 = s4 ? tmp22379 : tmp22382;
  assign tmp22377 = s5 ? tmp22378 : tmp22361;
  assign tmp22376 = s6 ? tmp22349 : tmp22377;
  assign tmp22367 = s7 ? tmp22368 : tmp22376;
  assign tmp22309 = s8 ? tmp22310 : tmp22367;
  assign tmp22389 = s3 ? tmp21943 : tmp22066;
  assign tmp22391 = s2 ? tmp22322 : tmp22134;
  assign tmp22390 = s3 ? tmp22037 : tmp22391;
  assign tmp22388 = s4 ? tmp22389 : tmp22390;
  assign tmp22396 = ~(s1 ? 1 : tmp22049);
  assign tmp22395 = s2 ? tmp21943 : tmp22396;
  assign tmp22394 = s3 ? tmp22058 : tmp22395;
  assign tmp22398 = ~(s2 ? tmp21943 : 0);
  assign tmp22397 = ~(s3 ? tmp22167 : tmp22398);
  assign tmp22393 = s4 ? tmp22394 : tmp22397;
  assign tmp22401 = s2 ? tmp22210 : tmp22256;
  assign tmp22403 = ~(s1 ? 1 : tmp22048);
  assign tmp22402 = s2 ? tmp22255 : tmp22403;
  assign tmp22400 = s3 ? tmp22401 : tmp22402;
  assign tmp22406 = ~(s1 ? tmp22048 : 0);
  assign tmp22405 = s2 ? tmp22210 : tmp22406;
  assign tmp22408 = s1 ? tmp22048 : 1;
  assign tmp22407 = ~(s2 ? tmp22198 : tmp22408);
  assign tmp22404 = s3 ? tmp22405 : tmp22407;
  assign tmp22399 = s4 ? tmp22400 : tmp22404;
  assign tmp22392 = s5 ? tmp22393 : tmp22399;
  assign tmp22387 = s6 ? tmp22388 : tmp22392;
  assign tmp22411 = s3 ? tmp22066 : tmp22152;
  assign tmp22410 = s4 ? tmp22389 : tmp22411;
  assign tmp22415 = s2 ? tmp22059 : tmp21943;
  assign tmp22414 = s3 ? tmp22415 : tmp22395;
  assign tmp22413 = s4 ? tmp22414 : tmp22397;
  assign tmp22418 = s2 ? tmp22210 : 1;
  assign tmp22419 = ~(s2 ? 1 : tmp22227);
  assign tmp22417 = s3 ? tmp22418 : tmp22419;
  assign tmp22421 = s2 ? 1 : tmp22049;
  assign tmp22420 = ~(s3 ? tmp22421 : tmp22227);
  assign tmp22416 = s4 ? tmp22417 : tmp22420;
  assign tmp22412 = s5 ? tmp22413 : tmp22416;
  assign tmp22409 = s6 ? tmp22410 : tmp22412;
  assign tmp22386 = ~(s7 ? tmp22387 : tmp22409);
  assign tmp22385 = s8 ? tmp22367 : tmp22386;
  assign tmp22308 = s9 ? tmp22309 : tmp22385;
  assign tmp22427 = s4 ? tmp22356 : tmp22382;
  assign tmp22426 = s5 ? tmp22427 : tmp22361;
  assign tmp22425 = s6 ? tmp22349 : tmp22426;
  assign tmp22424 = s7 ? tmp22311 : tmp22425;
  assign tmp22423 = s8 ? tmp22424 : tmp22311;
  assign tmp22433 = s3 ? tmp22359 : tmp22384;
  assign tmp22432 = s4 ? tmp22356 : tmp22433;
  assign tmp22431 = s5 ? tmp22432 : tmp22361;
  assign tmp22430 = s6 ? tmp22349 : tmp22431;
  assign tmp22434 = ~(s6 ? tmp22410 : tmp22412);
  assign tmp22429 = s7 ? tmp22430 : tmp22434;
  assign tmp22435 = s7 ? tmp22376 : tmp22425;
  assign tmp22428 = s8 ? tmp22429 : tmp22435;
  assign tmp22422 = s9 ? tmp22423 : tmp22428;
  assign tmp22307 = s10 ? tmp22308 : tmp22422;
  assign tmp22439 = s7 ? tmp22348 : tmp22434;
  assign tmp22438 = s8 ? tmp22439 : tmp22435;
  assign tmp22437 = s9 ? tmp22423 : tmp22438;
  assign tmp22436 = s10 ? tmp22308 : tmp22437;
  assign tmp22306 = s11 ? tmp22307 : tmp22436;
  assign tmp22305 = s12 ? 1 : tmp22306;
  assign tmp22450 = s1 ? tmp22046 : tmp21943;
  assign tmp22449 = s2 ? tmp21943 : tmp22450;
  assign tmp22448 = s3 ? tmp21943 : tmp22449;
  assign tmp22452 = s2 ? tmp21943 : tmp22046;
  assign tmp22454 = s1 ? tmp21943 : tmp22148;
  assign tmp22453 = s2 ? tmp22454 : tmp22039;
  assign tmp22451 = s3 ? tmp22452 : tmp22453;
  assign tmp22447 = s4 ? tmp22448 : tmp22451;
  assign tmp22459 = ~(s1 ? tmp22048 : tmp22119);
  assign tmp22458 = s2 ? tmp22110 : tmp22459;
  assign tmp22460 = ~(s2 ? tmp22048 : tmp22231);
  assign tmp22457 = s3 ? tmp22458 : tmp22460;
  assign tmp22462 = s2 ? tmp22060 : tmp21943;
  assign tmp22461 = s3 ? tmp22462 : tmp22074;
  assign tmp22456 = s4 ? tmp22457 : tmp22461;
  assign tmp22455 = s5 ? tmp22456 : tmp22056;
  assign tmp22446 = s6 ? tmp22447 : tmp22455;
  assign tmp22465 = s3 ? tmp22452 : tmp22038;
  assign tmp22464 = s4 ? tmp22448 : tmp22465;
  assign tmp22469 = s2 ? tmp22450 : tmp22045;
  assign tmp22468 = s3 ? tmp22469 : tmp22268;
  assign tmp22467 = s4 ? tmp22468 : tmp22461;
  assign tmp22472 = s2 ? tmp22059 : 1;
  assign tmp22471 = s3 ? tmp22415 : tmp22472;
  assign tmp22470 = s4 ? tmp22471 : tmp22078;
  assign tmp22466 = s5 ? tmp22467 : tmp22470;
  assign tmp22463 = s6 ? tmp22464 : tmp22466;
  assign tmp22445 = s7 ? tmp22446 : tmp22463;
  assign tmp22478 = ~(l3 ? 1 : 0);
  assign tmp22477 = l1 ? 1 : tmp22478;
  assign tmp22481 = s0 ? tmp22477 : tmp22478;
  assign tmp22480 = s1 ? tmp22481 : tmp22477;
  assign tmp22479 = s2 ? tmp22477 : tmp22480;
  assign tmp22476 = s3 ? tmp22477 : tmp22479;
  assign tmp22485 = s0 ? tmp22477 : tmp21943;
  assign tmp22484 = s1 ? tmp22485 : tmp22477;
  assign tmp22486 = s0 ? tmp22477 : 0;
  assign tmp22483 = s2 ? tmp22484 : tmp22486;
  assign tmp22488 = s1 ? tmp22477 : tmp22148;
  assign tmp22490 = s0 ? 1 : tmp22477;
  assign tmp22489 = s1 ? tmp22477 : tmp22490;
  assign tmp22487 = s2 ? tmp22488 : tmp22489;
  assign tmp22482 = s3 ? tmp22483 : tmp22487;
  assign tmp22475 = s4 ? tmp22476 : tmp22482;
  assign tmp22497 = ~(l1 ? 1 : tmp22478);
  assign tmp22496 = ~(s0 ? 1 : tmp22497);
  assign tmp22495 = s1 ? tmp22486 : tmp22496;
  assign tmp22499 = s0 ? 1 : tmp22497;
  assign tmp22500 = ~(s0 ? tmp22477 : tmp22478);
  assign tmp22498 = ~(s1 ? tmp22499 : tmp22500);
  assign tmp22494 = s2 ? tmp22495 : tmp22498;
  assign tmp22503 = l3 ? 1 : 0;
  assign tmp22502 = s0 ? tmp22503 : tmp22497;
  assign tmp22504 = ~(s1 ? 1 : tmp22477);
  assign tmp22501 = ~(s2 ? tmp22502 : tmp22504);
  assign tmp22493 = s3 ? tmp22494 : tmp22501;
  assign tmp22507 = s1 ? tmp22490 : tmp21951;
  assign tmp22508 = s1 ? tmp21951 : tmp22485;
  assign tmp22506 = s2 ? tmp22507 : tmp22508;
  assign tmp22510 = s1 ? tmp22477 : 1;
  assign tmp22509 = s2 ? tmp22510 : 1;
  assign tmp22505 = s3 ? tmp22506 : tmp22509;
  assign tmp22492 = s4 ? tmp22493 : tmp22505;
  assign tmp22515 = s0 ? tmp22477 : 1;
  assign tmp22514 = s1 ? tmp22515 : 1;
  assign tmp22513 = s2 ? tmp22514 : tmp22490;
  assign tmp22512 = s3 ? tmp22513 : 1;
  assign tmp22518 = s1 ? tmp22490 : tmp22515;
  assign tmp22517 = s2 ? 1 : tmp22518;
  assign tmp22516 = s3 ? tmp22517 : 1;
  assign tmp22511 = s4 ? tmp22512 : tmp22516;
  assign tmp22491 = s5 ? tmp22492 : tmp22511;
  assign tmp22474 = s6 ? tmp22475 : tmp22491;
  assign tmp22522 = s2 ? tmp22510 : tmp22489;
  assign tmp22521 = s3 ? tmp22483 : tmp22522;
  assign tmp22520 = s4 ? tmp22476 : tmp22521;
  assign tmp22527 = s1 ? tmp22486 : tmp22477;
  assign tmp22528 = s1 ? tmp22477 : tmp22481;
  assign tmp22526 = s2 ? tmp22527 : tmp22528;
  assign tmp22530 = s1 ? 1 : tmp22477;
  assign tmp22529 = s2 ? tmp22477 : tmp22530;
  assign tmp22525 = s3 ? tmp22526 : tmp22529;
  assign tmp22532 = s2 ? tmp22507 : tmp22477;
  assign tmp22531 = s3 ? tmp22532 : tmp22509;
  assign tmp22524 = s4 ? tmp22525 : tmp22531;
  assign tmp22535 = s2 ? tmp22514 : tmp22510;
  assign tmp22534 = s3 ? tmp22535 : tmp22472;
  assign tmp22538 = s1 ? tmp22477 : tmp21943;
  assign tmp22537 = s2 ? 1 : tmp22538;
  assign tmp22536 = s3 ? tmp22537 : 1;
  assign tmp22533 = s4 ? tmp22534 : tmp22536;
  assign tmp22523 = s5 ? tmp22524 : tmp22533;
  assign tmp22519 = s6 ? tmp22520 : tmp22523;
  assign tmp22473 = s7 ? tmp22474 : tmp22519;
  assign tmp22444 = s8 ? tmp22445 : tmp22473;
  assign tmp22542 = s5 ? tmp22467 : tmp22075;
  assign tmp22541 = s6 ? tmp22464 : tmp22542;
  assign tmp22540 = s7 ? tmp22446 : tmp22541;
  assign tmp22539 = s8 ? tmp22473 : tmp22540;
  assign tmp22443 = s9 ? tmp22444 : tmp22539;
  assign tmp22549 = s3 ? tmp22077 : tmp22472;
  assign tmp22548 = s4 ? tmp22549 : tmp22078;
  assign tmp22547 = s5 ? tmp22467 : tmp22548;
  assign tmp22546 = s6 ? tmp22464 : tmp22547;
  assign tmp22545 = s7 ? tmp22446 : tmp22546;
  assign tmp22544 = s8 ? tmp22545 : tmp22446;
  assign tmp22551 = s7 ? tmp22463 : tmp22541;
  assign tmp22557 = s2 ? 1 : tmp22477;
  assign tmp22556 = s3 ? tmp22557 : 1;
  assign tmp22555 = s4 ? tmp22534 : tmp22556;
  assign tmp22554 = s5 ? tmp22524 : tmp22555;
  assign tmp22553 = s6 ? tmp22520 : tmp22554;
  assign tmp22552 = s7 ? tmp22553 : tmp22546;
  assign tmp22550 = s8 ? tmp22551 : tmp22552;
  assign tmp22543 = s9 ? tmp22544 : tmp22550;
  assign tmp22442 = s10 ? tmp22443 : tmp22543;
  assign tmp22561 = s7 ? tmp22519 : tmp22546;
  assign tmp22560 = s8 ? tmp22551 : tmp22561;
  assign tmp22559 = s9 ? tmp22544 : tmp22560;
  assign tmp22558 = s10 ? tmp22443 : tmp22559;
  assign tmp22441 = s11 ? tmp22442 : tmp22558;
  assign tmp22570 = s3 ? 1 : tmp22472;
  assign tmp22569 = s4 ? tmp22570 : tmp22078;
  assign tmp22568 = s5 ? 1 : tmp22569;
  assign tmp22567 = s6 ? 1 : tmp22568;
  assign tmp22566 = s7 ? 1 : tmp22567;
  assign tmp22576 = s2 ? 1 : tmp22269;
  assign tmp22575 = s3 ? tmp22576 : 1;
  assign tmp22574 = s4 ? tmp22570 : tmp22575;
  assign tmp22573 = s5 ? 1 : tmp22574;
  assign tmp22572 = s6 ? 1 : tmp22573;
  assign tmp22571 = s7 ? 1 : tmp22572;
  assign tmp22565 = s8 ? tmp22566 : tmp22571;
  assign tmp22577 = s8 ? tmp22571 : 1;
  assign tmp22564 = s9 ? tmp22565 : tmp22577;
  assign tmp22579 = s8 ? tmp22566 : 1;
  assign tmp22584 = s4 ? tmp22570 : 1;
  assign tmp22583 = s5 ? 1 : tmp22584;
  assign tmp22582 = s6 ? 1 : tmp22583;
  assign tmp22581 = s7 ? tmp22582 : 1;
  assign tmp22580 = s8 ? tmp22581 : tmp22582;
  assign tmp22578 = s9 ? tmp22579 : tmp22580;
  assign tmp22563 = s10 ? tmp22564 : tmp22578;
  assign tmp22588 = s7 ? tmp22567 : 1;
  assign tmp22589 = s7 ? tmp22572 : tmp22567;
  assign tmp22587 = s8 ? tmp22588 : tmp22589;
  assign tmp22586 = s9 ? tmp22579 : tmp22587;
  assign tmp22585 = s10 ? tmp22564 : tmp22586;
  assign tmp22562 = s11 ? tmp22563 : tmp22585;
  assign tmp22440 = ~(s12 ? tmp22441 : tmp22562);
  assign tmp22304 = ~(s13 ? tmp22305 : tmp22440);
  assign tmp21929 = s14 ? tmp21930 : tmp22304;
  assign tmp22599 = s2 ? tmp22040 : tmp22269;
  assign tmp22598 = s3 ? 1 : tmp22599;
  assign tmp22601 = s2 ? tmp22269 : 1;
  assign tmp22603 = s1 ? 1 : tmp22040;
  assign tmp22602 = s2 ? tmp22603 : tmp21943;
  assign tmp22600 = s3 ? tmp22601 : tmp22602;
  assign tmp22597 = s4 ? tmp22598 : tmp22600;
  assign tmp22607 = s2 ? 1 : tmp22071;
  assign tmp22606 = s3 ? tmp22607 : tmp22602;
  assign tmp22608 = s3 ? tmp22074 : tmp22602;
  assign tmp22605 = s4 ? tmp22606 : tmp22608;
  assign tmp22611 = s2 ? tmp22206 : 1;
  assign tmp22612 = s2 ? tmp22603 : tmp22059;
  assign tmp22610 = s3 ? tmp22611 : tmp22612;
  assign tmp22613 = s3 ? tmp22612 : tmp22611;
  assign tmp22609 = s4 ? tmp22610 : tmp22613;
  assign tmp22604 = s5 ? tmp22605 : tmp22609;
  assign tmp22596 = s6 ? tmp22597 : tmp22604;
  assign tmp22617 = s2 ? tmp22269 : tmp21943;
  assign tmp22616 = s3 ? tmp22601 : tmp22617;
  assign tmp22615 = s4 ? tmp22598 : tmp22616;
  assign tmp22620 = s3 ? tmp22607 : tmp22617;
  assign tmp22621 = s3 ? tmp22074 : tmp22617;
  assign tmp22619 = s4 ? tmp22620 : tmp22621;
  assign tmp22623 = s3 ? tmp22611 : tmp22601;
  assign tmp22625 = s2 ? tmp22269 : tmp21951;
  assign tmp22624 = s3 ? tmp22625 : tmp21953;
  assign tmp22622 = s4 ? tmp22623 : tmp22624;
  assign tmp22618 = s5 ? tmp22619 : tmp22622;
  assign tmp22614 = s6 ? tmp22615 : tmp22618;
  assign tmp22595 = s7 ? tmp22596 : tmp22614;
  assign tmp22627 = s8 ? tmp22595 : tmp22596;
  assign tmp22631 = s3 ? tmp22601 : tmp21953;
  assign tmp22630 = s4 ? tmp22623 : tmp22631;
  assign tmp22629 = s5 ? tmp22619 : tmp22630;
  assign tmp22628 = s6 ? tmp22615 : tmp22629;
  assign tmp22626 = s9 ? tmp22627 : tmp22628;
  assign tmp22594 = s10 ? tmp22595 : tmp22626;
  assign tmp22633 = s9 ? tmp22627 : tmp22614;
  assign tmp22632 = s10 ? tmp22595 : tmp22633;
  assign tmp22593 = s11 ? tmp22594 : tmp22632;
  assign tmp22638 = s3 ? tmp22116 : tmp21943;
  assign tmp22637 = s4 ? tmp22638 : tmp21943;
  assign tmp22642 = s2 ? 1 : tmp22227;
  assign tmp22641 = s3 ? tmp22642 : tmp22049;
  assign tmp22640 = s4 ? tmp22641 : tmp22049;
  assign tmp22645 = ~(s2 ? 1 : tmp22168);
  assign tmp22644 = s3 ? tmp21943 : tmp22645;
  assign tmp22647 = ~(s1 ? tmp22046 : 0);
  assign tmp22646 = ~(s2 ? tmp22198 : tmp22647);
  assign tmp22643 = ~(s4 ? tmp22644 : tmp22646);
  assign tmp22639 = ~(s5 ? tmp22640 : tmp22643);
  assign tmp22636 = s6 ? tmp22637 : tmp22639;
  assign tmp22652 = ~(s2 ? 1 : tmp22049);
  assign tmp22651 = s3 ? tmp21943 : tmp22652;
  assign tmp22653 = ~(s2 ? tmp22227 : 1);
  assign tmp22650 = ~(s4 ? tmp22651 : tmp22653);
  assign tmp22649 = ~(s5 ? tmp22640 : tmp22650);
  assign tmp22648 = s6 ? tmp22637 : tmp22649;
  assign tmp22635 = s7 ? tmp22636 : tmp22648;
  assign tmp22655 = s8 ? tmp22635 : tmp22636;
  assign tmp22654 = s9 ? tmp22655 : tmp22648;
  assign tmp22634 = s10 ? tmp22635 : tmp22654;
  assign tmp22592 = s12 ? tmp22593 : tmp22634;
  assign tmp22662 = s2 ? tmp22168 : tmp22123;
  assign tmp22661 = s3 ? tmp22048 : tmp22662;
  assign tmp22664 = s2 ? tmp22227 : tmp22647;
  assign tmp22665 = s2 ? tmp22198 : tmp22049;
  assign tmp22663 = s3 ? tmp22664 : tmp22665;
  assign tmp22660 = s4 ? tmp22661 : tmp22663;
  assign tmp22669 = s2 ? tmp22210 : tmp22459;
  assign tmp22670 = ~(s2 ? tmp22048 : tmp22049);
  assign tmp22668 = s3 ? tmp22669 : tmp22670;
  assign tmp22672 = s2 ? tmp22116 : 0;
  assign tmp22671 = s3 ? tmp22672 : tmp22670;
  assign tmp22667 = s4 ? tmp22668 : tmp22671;
  assign tmp22675 = s2 ? tmp22039 : tmp22210;
  assign tmp22677 = ~(s1 ? tmp21943 : tmp22046);
  assign tmp22676 = ~(s2 ? tmp22198 : tmp22677);
  assign tmp22674 = s3 ? tmp22675 : tmp22676;
  assign tmp22680 = ~(s1 ? tmp22040 : 0);
  assign tmp22679 = s2 ? tmp22168 : tmp22680;
  assign tmp22681 = ~(s2 ? tmp21943 : tmp22110);
  assign tmp22678 = ~(s3 ? tmp22679 : tmp22681);
  assign tmp22673 = s4 ? tmp22674 : tmp22678;
  assign tmp22666 = ~(s5 ? tmp22667 : tmp22673);
  assign tmp22659 = s6 ? tmp22660 : tmp22666;
  assign tmp22685 = s2 ? tmp22227 : tmp22049;
  assign tmp22684 = s3 ? tmp22664 : tmp22685;
  assign tmp22683 = s4 ? tmp22661 : tmp22684;
  assign tmp22689 = s2 ? tmp22210 : tmp22045;
  assign tmp22688 = s3 ? tmp22689 : tmp21943;
  assign tmp22687 = s4 ? tmp22688 : tmp22671;
  assign tmp22692 = s2 ? tmp21943 : 0;
  assign tmp22693 = ~(s2 ? tmp22227 : tmp22677);
  assign tmp22691 = s3 ? tmp22692 : tmp22693;
  assign tmp22690 = s4 ? tmp22691 : tmp21943;
  assign tmp22686 = ~(s5 ? tmp22687 : tmp22690);
  assign tmp22682 = s6 ? tmp22683 : tmp22686;
  assign tmp22658 = s7 ? tmp22659 : tmp22682;
  assign tmp22695 = s8 ? tmp22658 : tmp22659;
  assign tmp22694 = s9 ? tmp22695 : tmp22682;
  assign tmp22657 = s10 ? tmp22658 : tmp22694;
  assign tmp22700 = s3 ? tmp21953 : tmp22599;
  assign tmp22702 = s2 ? tmp22269 : tmp22059;
  assign tmp22701 = s3 ? tmp22702 : tmp22602;
  assign tmp22699 = s4 ? tmp22700 : tmp22701;
  assign tmp22707 = ~(s1 ? 1 : tmp22119);
  assign tmp22706 = s2 ? tmp22040 : tmp22707;
  assign tmp22705 = s3 ? tmp22074 : tmp22706;
  assign tmp22704 = s4 ? tmp22606 : tmp22705;
  assign tmp22710 = s2 ? tmp22060 : tmp22206;
  assign tmp22709 = s3 ? tmp22055 : tmp22710;
  assign tmp22712 = s2 ? tmp22060 : tmp21951;
  assign tmp22711 = s3 ? tmp22702 : tmp22712;
  assign tmp22708 = s4 ? tmp22709 : tmp22711;
  assign tmp22703 = s5 ? tmp22704 : tmp22708;
  assign tmp22698 = s6 ? tmp22699 : tmp22703;
  assign tmp22715 = s3 ? tmp22702 : tmp22617;
  assign tmp22714 = s4 ? tmp22700 : tmp22715;
  assign tmp22719 = s2 ? tmp22060 : tmp22396;
  assign tmp22718 = s3 ? tmp22074 : tmp22719;
  assign tmp22717 = s4 ? tmp22620 : tmp22718;
  assign tmp22721 = s3 ? tmp22074 : tmp22262;
  assign tmp22722 = s3 ? tmp22055 : tmp21943;
  assign tmp22720 = s4 ? tmp22721 : tmp22722;
  assign tmp22716 = s5 ? tmp22717 : tmp22720;
  assign tmp22713 = s6 ? tmp22714 : tmp22716;
  assign tmp22697 = s7 ? tmp22698 : tmp22713;
  assign tmp22724 = s8 ? tmp22697 : tmp22698;
  assign tmp22723 = s9 ? tmp22724 : tmp22713;
  assign tmp22696 = ~(s10 ? tmp22697 : tmp22723);
  assign tmp22656 = ~(s12 ? tmp22657 : tmp22696);
  assign tmp22591 = s13 ? tmp22592 : tmp22656;
  assign tmp22735 = s2 ? tmp22054 : tmp21951;
  assign tmp22736 = s2 ? tmp22322 : tmp21943;
  assign tmp22734 = s3 ? tmp22735 : tmp22736;
  assign tmp22733 = s4 ? tmp22389 : tmp22734;
  assign tmp22739 = s3 ? tmp22058 : tmp22449;
  assign tmp22742 = ~(s1 ? tmp21943 : tmp21951);
  assign tmp22741 = s2 ? tmp22168 : tmp22742;
  assign tmp22740 = ~(s3 ? tmp22741 : tmp22398);
  assign tmp22738 = s4 ? tmp22739 : tmp22740;
  assign tmp22745 = s2 ? tmp22110 : tmp22059;
  assign tmp22744 = s3 ? tmp22745 : tmp22402;
  assign tmp22747 = s2 ? tmp21943 : tmp22406;
  assign tmp22748 = s2 ? tmp22134 : tmp22111;
  assign tmp22746 = s3 ? tmp22747 : tmp22748;
  assign tmp22743 = s4 ? tmp22744 : tmp22746;
  assign tmp22737 = s5 ? tmp22738 : tmp22743;
  assign tmp22732 = s6 ? tmp22733 : tmp22737;
  assign tmp22752 = s2 ? tmp22116 : tmp21943;
  assign tmp22751 = s3 ? tmp22054 : tmp22752;
  assign tmp22750 = s4 ? tmp22389 : tmp22751;
  assign tmp22755 = s3 ? tmp22415 : tmp22449;
  assign tmp22754 = s4 ? tmp22755 : tmp22397;
  assign tmp22758 = s2 ? tmp22450 : 1;
  assign tmp22759 = s2 ? tmp22210 : tmp22396;
  assign tmp22757 = s3 ? tmp22758 : tmp22759;
  assign tmp22756 = s4 ? tmp22757 : tmp21943;
  assign tmp22753 = s5 ? tmp22754 : tmp22756;
  assign tmp22749 = s6 ? tmp22750 : tmp22753;
  assign tmp22731 = s7 ? tmp22732 : tmp22749;
  assign tmp22767 = l4 ? 1 : 0;
  assign tmp22766 = l2 ? tmp22767 : 0;
  assign tmp22765 = l1 ? 1 : tmp22766;
  assign tmp22769 = l1 ? 1 : tmp22767;
  assign tmp22768 = s0 ? tmp22769 : tmp22765;
  assign tmp22764 = s1 ? tmp22765 : tmp22768;
  assign tmp22772 = s0 ? tmp22769 : 1;
  assign tmp22771 = s1 ? tmp22772 : tmp22765;
  assign tmp22770 = s2 ? tmp22765 : tmp22771;
  assign tmp22763 = s3 ? tmp22764 : tmp22770;
  assign tmp22776 = s0 ? tmp22765 : 1;
  assign tmp22775 = s1 ? tmp22776 : tmp22765;
  assign tmp22777 = s1 ? tmp22776 : tmp22772;
  assign tmp22774 = s2 ? tmp22775 : tmp22777;
  assign tmp22779 = s1 ? tmp22769 : tmp22147;
  assign tmp22778 = s2 ? tmp22779 : tmp22765;
  assign tmp22773 = s3 ? tmp22774 : tmp22778;
  assign tmp22762 = s4 ? tmp22763 : tmp22773;
  assign tmp22784 = s1 ? tmp22776 : 1;
  assign tmp22786 = s0 ? 1 : tmp22765;
  assign tmp22785 = s1 ? tmp22786 : tmp22776;
  assign tmp22783 = s2 ? tmp22784 : tmp22785;
  assign tmp22789 = s0 ? tmp22765 : 0;
  assign tmp22788 = s1 ? tmp22789 : tmp22765;
  assign tmp22787 = s2 ? tmp22786 : tmp22788;
  assign tmp22782 = s3 ? tmp22783 : tmp22787;
  assign tmp22794 = ~(l1 ? 1 : tmp22766);
  assign tmp22793 = s0 ? 1 : tmp22794;
  assign tmp22795 = ~(s0 ? 1 : tmp22769);
  assign tmp22792 = s1 ? tmp22793 : tmp22795;
  assign tmp22797 = s0 ? 1 : tmp22769;
  assign tmp22796 = ~(s1 ? tmp22797 : tmp22776);
  assign tmp22791 = s2 ? tmp22792 : tmp22796;
  assign tmp22800 = s0 ? tmp22769 : tmp21943;
  assign tmp22799 = s1 ? tmp22765 : tmp22800;
  assign tmp22798 = ~(s2 ? tmp22799 : 0);
  assign tmp22790 = ~(s3 ? tmp22791 : tmp22798);
  assign tmp22781 = s4 ? tmp22782 : tmp22790;
  assign tmp22806 = ~(l1 ? 1 : tmp22767);
  assign tmp22805 = ~(s0 ? 1 : tmp22806);
  assign tmp22804 = s1 ? tmp22789 : tmp22805;
  assign tmp22807 = s1 ? tmp22772 : 1;
  assign tmp22803 = s2 ? tmp22804 : tmp22807;
  assign tmp22802 = s3 ? tmp22803 : tmp22402;
  assign tmp22811 = s0 ? tmp21943 : tmp22765;
  assign tmp22810 = s1 ? tmp21943 : tmp22811;
  assign tmp22812 = ~(s1 ? tmp22793 : 0);
  assign tmp22809 = s2 ? tmp22810 : tmp22812;
  assign tmp22814 = s1 ? tmp22800 : tmp22111;
  assign tmp22813 = s2 ? tmp22814 : tmp22111;
  assign tmp22808 = s3 ? tmp22809 : tmp22813;
  assign tmp22801 = s4 ? tmp22802 : tmp22808;
  assign tmp22780 = s5 ? tmp22781 : tmp22801;
  assign tmp22761 = s6 ? tmp22762 : tmp22780;
  assign tmp22819 = s1 ? tmp22776 : tmp22769;
  assign tmp22818 = s2 ? tmp22775 : tmp22819;
  assign tmp22821 = s1 ? tmp22769 : 0;
  assign tmp22820 = s2 ? tmp22821 : tmp22765;
  assign tmp22817 = s3 ? tmp22818 : tmp22820;
  assign tmp22816 = s4 ? tmp22763 : tmp22817;
  assign tmp22826 = s1 ? tmp22765 : tmp22776;
  assign tmp22825 = s2 ? tmp22784 : tmp22826;
  assign tmp22827 = s2 ? tmp22765 : tmp22788;
  assign tmp22824 = s3 ? tmp22825 : tmp22827;
  assign tmp22829 = s2 ? tmp22792 : tmp22794;
  assign tmp22831 = s1 ? tmp22765 : tmp21943;
  assign tmp22830 = ~(s2 ? tmp22831 : 0);
  assign tmp22828 = ~(s3 ? tmp22829 : tmp22830);
  assign tmp22823 = s4 ? tmp22824 : tmp22828;
  assign tmp22835 = s1 ? tmp22789 : tmp22769;
  assign tmp22834 = s2 ? tmp22835 : 1;
  assign tmp22833 = s3 ? tmp22834 : tmp22759;
  assign tmp22838 = s1 ? tmp21943 : tmp22765;
  assign tmp22837 = s2 ? tmp22838 : tmp22831;
  assign tmp22836 = s3 ? tmp22837 : tmp21943;
  assign tmp22832 = s4 ? tmp22833 : tmp22836;
  assign tmp22822 = s5 ? tmp22823 : tmp22832;
  assign tmp22815 = s6 ? tmp22816 : tmp22822;
  assign tmp22760 = s7 ? tmp22761 : tmp22815;
  assign tmp22730 = s8 ? tmp22731 : tmp22760;
  assign tmp22845 = s2 ? tmp22255 : tmp22396;
  assign tmp22844 = s3 ? tmp22758 : tmp22845;
  assign tmp22843 = s4 ? tmp22844 : tmp21943;
  assign tmp22842 = s5 ? tmp22754 : tmp22843;
  assign tmp22841 = s6 ? tmp22750 : tmp22842;
  assign tmp22840 = s7 ? tmp22732 : tmp22841;
  assign tmp22839 = s8 ? tmp22760 : tmp22840;
  assign tmp22729 = s9 ? tmp22730 : tmp22839;
  assign tmp22847 = s8 ? tmp22731 : tmp22732;
  assign tmp22849 = s7 ? tmp22749 : tmp22841;
  assign tmp22855 = s2 ? tmp22838 : tmp22765;
  assign tmp22854 = s3 ? tmp22855 : tmp21943;
  assign tmp22853 = s4 ? tmp22833 : tmp22854;
  assign tmp22852 = s5 ? tmp22823 : tmp22853;
  assign tmp22851 = s6 ? tmp22816 : tmp22852;
  assign tmp22850 = s7 ? tmp22851 : tmp22749;
  assign tmp22848 = s8 ? tmp22849 : tmp22850;
  assign tmp22846 = s9 ? tmp22847 : tmp22848;
  assign tmp22728 = s10 ? tmp22729 : tmp22846;
  assign tmp22859 = s7 ? tmp22815 : tmp22749;
  assign tmp22858 = s8 ? tmp22849 : tmp22859;
  assign tmp22857 = s9 ? tmp22847 : tmp22858;
  assign tmp22856 = s10 ? tmp22729 : tmp22857;
  assign tmp22727 = s11 ? tmp22728 : tmp22856;
  assign tmp22869 = ~(l1 ? 1 : tmp21941);
  assign tmp22868 = s0 ? 1 : tmp22869;
  assign tmp22871 = s1 ? tmp21956 : tmp21940;
  assign tmp22873 = s0 ? tmp21940 : 0;
  assign tmp22872 = s1 ? tmp22873 : tmp21940;
  assign tmp22870 = ~(s2 ? tmp22871 : tmp22872);
  assign tmp22867 = s3 ? tmp22868 : tmp22870;
  assign tmp22877 = s0 ? tmp21940 : tmp22049;
  assign tmp22876 = s1 ? tmp22877 : tmp21940;
  assign tmp22878 = s1 ? tmp22873 : 0;
  assign tmp22875 = s2 ? tmp22876 : tmp22878;
  assign tmp22880 = ~(s1 ? tmp21940 : tmp21942);
  assign tmp22879 = ~(s2 ? tmp22198 : tmp22880);
  assign tmp22874 = ~(s3 ? tmp22875 : tmp22879);
  assign tmp22866 = s4 ? tmp22867 : tmp22874;
  assign tmp22885 = s1 ? tmp21950 : 1;
  assign tmp22886 = s1 ? tmp21956 : tmp22873;
  assign tmp22884 = s2 ? tmp22885 : tmp22886;
  assign tmp22888 = ~(s1 ? tmp21951 : tmp21940);
  assign tmp22887 = ~(s2 ? tmp22868 : tmp22888);
  assign tmp22883 = s3 ? tmp22884 : tmp22887;
  assign tmp22891 = s1 ? tmp21942 : tmp22140;
  assign tmp22893 = ~(s0 ? tmp21940 : tmp22049);
  assign tmp22892 = ~(s1 ? tmp21951 : tmp22893);
  assign tmp22890 = s2 ? tmp22891 : tmp22892;
  assign tmp22896 = ~(s0 ? 1 : tmp22869);
  assign tmp22895 = s1 ? tmp21940 : tmp22896;
  assign tmp22894 = s2 ? tmp22895 : tmp22071;
  assign tmp22889 = s3 ? tmp22890 : tmp22894;
  assign tmp22882 = s4 ? tmp22883 : tmp22889;
  assign tmp22900 = s1 ? tmp21950 : tmp22040;
  assign tmp22899 = s2 ? tmp22900 : tmp22059;
  assign tmp22902 = s1 ? tmp21943 : tmp21942;
  assign tmp22901 = s2 ? 1 : tmp22902;
  assign tmp22898 = s3 ? tmp22899 : tmp22901;
  assign tmp22905 = s1 ? tmp21956 : 1;
  assign tmp22904 = s2 ? tmp21988 : tmp22905;
  assign tmp22907 = s1 ? tmp21943 : tmp21956;
  assign tmp22908 = s1 ? tmp21942 : 1;
  assign tmp22906 = s2 ? tmp22907 : tmp22908;
  assign tmp22903 = s3 ? tmp22904 : tmp22906;
  assign tmp22897 = s4 ? tmp22898 : tmp22903;
  assign tmp22881 = ~(s5 ? tmp22882 : tmp22897);
  assign tmp22865 = s6 ? tmp22866 : tmp22881;
  assign tmp22912 = ~(s2 ? tmp22227 : tmp22880);
  assign tmp22911 = ~(s3 ? tmp22875 : tmp22912);
  assign tmp22910 = s4 ? tmp22867 : tmp22911;
  assign tmp22917 = s1 ? tmp21940 : tmp22873;
  assign tmp22916 = s2 ? tmp22885 : tmp22917;
  assign tmp22919 = s1 ? tmp21951 : tmp21940;
  assign tmp22918 = s2 ? tmp21940 : tmp22919;
  assign tmp22915 = s3 ? tmp22916 : tmp22918;
  assign tmp22921 = s2 ? tmp22891 : tmp21940;
  assign tmp22922 = s2 ? tmp21940 : tmp22269;
  assign tmp22920 = s3 ? tmp22921 : tmp22922;
  assign tmp22914 = s4 ? tmp22915 : tmp22920;
  assign tmp22925 = s2 ? tmp21988 : tmp22059;
  assign tmp22926 = s2 ? 1 : tmp22094;
  assign tmp22924 = s3 ? tmp22925 : tmp22926;
  assign tmp22928 = s2 ? tmp21943 : tmp21940;
  assign tmp22927 = s3 ? tmp22928 : tmp22094;
  assign tmp22923 = s4 ? tmp22924 : tmp22927;
  assign tmp22913 = ~(s5 ? tmp22914 : tmp22923);
  assign tmp22909 = s6 ? tmp22910 : tmp22913;
  assign tmp22864 = s7 ? tmp22865 : tmp22909;
  assign tmp22934 = s0 ? tmp22767 : tmp22769;
  assign tmp22933 = s1 ? tmp22769 : tmp22934;
  assign tmp22936 = s1 ? tmp22797 : tmp22769;
  assign tmp22937 = s1 ? tmp22772 : tmp22769;
  assign tmp22935 = s2 ? tmp22936 : tmp22937;
  assign tmp22932 = s3 ? tmp22933 : tmp22935;
  assign tmp22941 = s0 ? tmp22769 : 0;
  assign tmp22942 = s0 ? tmp22767 : 0;
  assign tmp22940 = s1 ? tmp22941 : tmp22942;
  assign tmp22939 = s2 ? tmp22937 : tmp22940;
  assign tmp22944 = s1 ? tmp22767 : tmp22111;
  assign tmp22943 = s2 ? tmp22944 : tmp22769;
  assign tmp22938 = s3 ? tmp22939 : tmp22943;
  assign tmp22931 = s4 ? tmp22932 : tmp22938;
  assign tmp22949 = s1 ? tmp22797 : tmp22772;
  assign tmp22948 = s2 ? tmp22807 : tmp22949;
  assign tmp22950 = s2 ? tmp22797 : tmp22937;
  assign tmp22947 = s3 ? tmp22948 : tmp22950;
  assign tmp22954 = s0 ? tmp21943 : tmp22769;
  assign tmp22955 = s0 ? 1 : tmp22767;
  assign tmp22953 = s1 ? tmp22954 : tmp22955;
  assign tmp22956 = s1 ? tmp22955 : tmp22772;
  assign tmp22952 = s2 ? tmp22953 : tmp22956;
  assign tmp22959 = s0 ? tmp22767 : tmp21940;
  assign tmp22958 = s1 ? tmp22769 : tmp22959;
  assign tmp22957 = s2 ? tmp22958 : tmp22071;
  assign tmp22951 = s3 ? tmp22952 : tmp22957;
  assign tmp22946 = s4 ? tmp22947 : tmp22951;
  assign tmp22963 = s1 ? tmp22772 : tmp22797;
  assign tmp22962 = s2 ? tmp22963 : tmp22807;
  assign tmp22961 = s3 ? tmp22962 : tmp22901;
  assign tmp22966 = s1 ? tmp21950 : tmp22797;
  assign tmp22967 = s1 ? tmp22797 : 1;
  assign tmp22965 = s2 ? tmp22966 : tmp22967;
  assign tmp22969 = s1 ? tmp22772 : tmp21956;
  assign tmp22968 = s2 ? tmp22969 : tmp22908;
  assign tmp22964 = s3 ? tmp22965 : tmp22968;
  assign tmp22960 = s4 ? tmp22961 : tmp22964;
  assign tmp22945 = s5 ? tmp22946 : tmp22960;
  assign tmp22930 = s6 ? tmp22931 : tmp22945;
  assign tmp22974 = s1 ? tmp22941 : tmp22767;
  assign tmp22973 = s2 ? tmp22937 : tmp22974;
  assign tmp22976 = s1 ? tmp22767 : tmp21943;
  assign tmp22975 = s2 ? tmp22976 : tmp22769;
  assign tmp22972 = s3 ? tmp22973 : tmp22975;
  assign tmp22971 = s4 ? tmp22932 : tmp22972;
  assign tmp22981 = s1 ? tmp22769 : tmp22772;
  assign tmp22980 = s2 ? tmp22807 : tmp22981;
  assign tmp22982 = s2 ? tmp22769 : tmp22937;
  assign tmp22979 = s3 ? tmp22980 : tmp22982;
  assign tmp22984 = s2 ? tmp22953 : tmp22769;
  assign tmp22986 = s1 ? tmp22769 : tmp21940;
  assign tmp22985 = s2 ? tmp22986 : tmp22269;
  assign tmp22983 = s3 ? tmp22984 : tmp22985;
  assign tmp22978 = s4 ? tmp22979 : tmp22983;
  assign tmp22989 = s2 ? tmp22937 : 1;
  assign tmp22988 = s3 ? tmp22989 : tmp22926;
  assign tmp22992 = s1 ? 1 : tmp22769;
  assign tmp22991 = s2 ? tmp22992 : tmp22769;
  assign tmp22993 = s1 ? 1 : tmp21940;
  assign tmp22990 = s3 ? tmp22991 : tmp22993;
  assign tmp22987 = s4 ? tmp22988 : tmp22990;
  assign tmp22977 = s5 ? tmp22978 : tmp22987;
  assign tmp22970 = s6 ? tmp22971 : tmp22977;
  assign tmp22929 = ~(s7 ? tmp22930 : tmp22970);
  assign tmp22863 = s8 ? tmp22864 : tmp22929;
  assign tmp22995 = s7 ? tmp22930 : tmp22970;
  assign tmp23000 = ~(s2 ? tmp22060 : tmp21943);
  assign tmp22999 = s3 ? tmp22048 : tmp23000;
  assign tmp23002 = s2 ? tmp22054 : tmp22210;
  assign tmp23003 = ~(s2 ? tmp22198 : tmp22049);
  assign tmp23001 = ~(s3 ? tmp23002 : tmp23003);
  assign tmp22998 = s4 ? tmp22999 : tmp23001;
  assign tmp23006 = s3 ? tmp22058 : tmp22066;
  assign tmp23009 = s1 ? tmp22147 : tmp21951;
  assign tmp23008 = s2 ? tmp22322 : tmp23009;
  assign tmp23010 = s2 ? tmp22134 : tmp22071;
  assign tmp23007 = s3 ? tmp23008 : tmp23010;
  assign tmp23005 = s4 ? tmp23006 : tmp23007;
  assign tmp23014 = s1 ? tmp21951 : tmp22040;
  assign tmp23013 = s2 ? tmp23014 : tmp22059;
  assign tmp23012 = s3 ? tmp23013 : tmp22079;
  assign tmp23017 = s1 ? tmp22040 : 1;
  assign tmp23016 = s2 ? tmp22054 : tmp23017;
  assign tmp23018 = s2 ? tmp22039 : tmp21953;
  assign tmp23015 = s3 ? tmp23016 : tmp23018;
  assign tmp23011 = s4 ? tmp23012 : tmp23015;
  assign tmp23004 = ~(s5 ? tmp23005 : tmp23011);
  assign tmp22997 = s6 ? tmp22998 : tmp23004;
  assign tmp23022 = ~(s2 ? tmp22227 : tmp22049);
  assign tmp23021 = ~(s3 ? tmp23002 : tmp23022);
  assign tmp23020 = s4 ? tmp22999 : tmp23021;
  assign tmp23025 = s3 ? tmp22415 : tmp22066;
  assign tmp23026 = s3 ? tmp22736 : tmp22268;
  assign tmp23024 = s4 ? tmp23025 : tmp23026;
  assign tmp23029 = s2 ? tmp22054 : 1;
  assign tmp23028 = s3 ? tmp23029 : tmp22079;
  assign tmp23027 = s4 ? tmp23028 : tmp21943;
  assign tmp23023 = ~(s5 ? tmp23024 : tmp23027);
  assign tmp23019 = s6 ? tmp23020 : tmp23023;
  assign tmp22996 = ~(s7 ? tmp22997 : tmp23019);
  assign tmp22994 = ~(s8 ? tmp22995 : tmp22996);
  assign tmp22862 = s9 ? tmp22863 : tmp22994;
  assign tmp23036 = ~(s2 ? tmp22871 : tmp21940);
  assign tmp23035 = s3 ? tmp22868 : tmp23036;
  assign tmp23039 = s1 ? tmp21950 : tmp21940;
  assign tmp23038 = s2 ? tmp23039 : tmp22878;
  assign tmp23037 = ~(s3 ? tmp23038 : tmp22879);
  assign tmp23034 = s4 ? tmp23035 : tmp23037;
  assign tmp23043 = s2 ? tmp22885 : tmp22871;
  assign tmp23042 = s3 ? tmp23043 : tmp22918;
  assign tmp23046 = s1 ? tmp21942 : tmp22147;
  assign tmp23047 = s1 ? tmp22147 : tmp21950;
  assign tmp23045 = s2 ? tmp23046 : tmp23047;
  assign tmp23044 = s3 ? tmp23045 : tmp22894;
  assign tmp23041 = s4 ? tmp23042 : tmp23044;
  assign tmp23040 = ~(s5 ? tmp23041 : tmp22897);
  assign tmp23033 = s6 ? tmp23034 : tmp23040;
  assign tmp23050 = ~(s3 ? tmp23038 : tmp22912);
  assign tmp23049 = s4 ? tmp23035 : tmp23050;
  assign tmp23054 = s2 ? tmp22885 : tmp21940;
  assign tmp23053 = s3 ? tmp23054 : tmp22918;
  assign tmp23056 = s2 ? tmp23046 : tmp21940;
  assign tmp23055 = s3 ? tmp23056 : tmp22922;
  assign tmp23052 = s4 ? tmp23053 : tmp23055;
  assign tmp23059 = s2 ? tmp21988 : 1;
  assign tmp23058 = s3 ? tmp23059 : tmp22926;
  assign tmp23060 = s3 ? tmp22928 : tmp22993;
  assign tmp23057 = s4 ? tmp23058 : tmp23060;
  assign tmp23051 = ~(s5 ? tmp23052 : tmp23057);
  assign tmp23048 = s6 ? tmp23049 : tmp23051;
  assign tmp23032 = s7 ? tmp23033 : tmp23048;
  assign tmp23031 = s8 ? tmp23032 : tmp23033;
  assign tmp23065 = s4 ? tmp22924 : tmp23060;
  assign tmp23064 = ~(s5 ? tmp22914 : tmp23065);
  assign tmp23063 = s6 ? tmp22910 : tmp23064;
  assign tmp23062 = s7 ? tmp23063 : tmp23019;
  assign tmp23067 = ~(s6 ? tmp23049 : tmp23051);
  assign tmp23066 = ~(s7 ? tmp22970 : tmp23067);
  assign tmp23061 = s8 ? tmp23062 : tmp23066;
  assign tmp23030 = s9 ? tmp23031 : tmp23061;
  assign tmp22861 = s10 ? tmp22862 : tmp23030;
  assign tmp23071 = s7 ? tmp22909 : tmp23019;
  assign tmp23070 = s8 ? tmp23071 : tmp23066;
  assign tmp23069 = s9 ? tmp23031 : tmp23070;
  assign tmp23068 = s10 ? tmp22862 : tmp23069;
  assign tmp22860 = ~(s11 ? tmp22861 : tmp23068);
  assign tmp22726 = s12 ? tmp22727 : tmp22860;
  assign tmp23078 = s2 ? tmp22048 : tmp22227;
  assign tmp23077 = s3 ? tmp22198 : tmp23078;
  assign tmp23080 = s2 ? tmp22227 : 1;
  assign tmp23079 = s3 ? tmp23080 : tmp22665;
  assign tmp23076 = s4 ? tmp23077 : tmp23079;
  assign tmp23083 = s3 ? tmp22669 : tmp23003;
  assign tmp23085 = s2 ? tmp22408 : 1;
  assign tmp23086 = s2 ? tmp22198 : tmp22118;
  assign tmp23084 = ~(s3 ? tmp23085 : tmp23086);
  assign tmp23082 = s4 ? tmp23083 : tmp23084;
  assign tmp23089 = ~(s2 ? tmp22168 : tmp22647);
  assign tmp23088 = s3 ? tmp22250 : tmp23089;
  assign tmp23091 = s2 ? tmp22168 : tmp22408;
  assign tmp23092 = s2 ? tmp22168 : tmp22227;
  assign tmp23090 = ~(s3 ? tmp23091 : tmp23092);
  assign tmp23087 = s4 ? tmp23088 : tmp23090;
  assign tmp23081 = ~(s5 ? tmp23082 : tmp23087);
  assign tmp23075 = s6 ? tmp23076 : tmp23081;
  assign tmp23095 = s3 ? tmp23080 : tmp22685;
  assign tmp23094 = s4 ? tmp23077 : tmp23095;
  assign tmp23098 = s3 ? tmp22689 : tmp23022;
  assign tmp23099 = ~(s3 ? tmp23085 : tmp22227);
  assign tmp23097 = s4 ? tmp23098 : tmp23099;
  assign tmp23101 = s3 ? tmp22250 : tmp22692;
  assign tmp23100 = s4 ? tmp23101 : tmp21943;
  assign tmp23096 = ~(s5 ? tmp23097 : tmp23100);
  assign tmp23093 = s6 ? tmp23094 : tmp23096;
  assign tmp23074 = s7 ? tmp23075 : tmp23093;
  assign tmp23103 = s8 ? tmp23074 : tmp23075;
  assign tmp23102 = s9 ? tmp23103 : tmp23093;
  assign tmp23073 = s10 ? tmp23074 : tmp23102;
  assign tmp23112 = s1 ? tmp22769 : tmp22797;
  assign tmp23113 = s2 ? tmp22797 : tmp22992;
  assign tmp23111 = s3 ? tmp23112 : tmp23113;
  assign tmp23116 = s1 ? tmp22769 : 1;
  assign tmp23115 = s2 ? tmp22937 : tmp23116;
  assign tmp23118 = s1 ? tmp22769 : tmp22954;
  assign tmp23117 = s2 ? tmp22269 : tmp23118;
  assign tmp23114 = s3 ? tmp23115 : tmp23117;
  assign tmp23110 = s4 ? tmp23111 : tmp23114;
  assign tmp23123 = s1 ? 1 : tmp22797;
  assign tmp23124 = s1 ? tmp21951 : tmp22769;
  assign tmp23122 = s2 ? tmp23123 : tmp23124;
  assign tmp23121 = s3 ? tmp22948 : tmp23122;
  assign tmp23127 = s1 ? tmp22954 : 1;
  assign tmp23128 = s1 ? 1 : tmp22772;
  assign tmp23126 = s2 ? tmp23127 : tmp23128;
  assign tmp23129 = s2 ? tmp23112 : tmp22071;
  assign tmp23125 = s3 ? tmp23126 : tmp23129;
  assign tmp23120 = s4 ? tmp23121 : tmp23125;
  assign tmp23132 = s2 ? tmp22807 : 1;
  assign tmp23134 = s1 ? tmp22040 : tmp22954;
  assign tmp23133 = s2 ? tmp22053 : tmp23134;
  assign tmp23131 = s3 ? tmp23132 : tmp23133;
  assign tmp23137 = s1 ? tmp22800 : tmp21943;
  assign tmp23136 = s2 ? tmp23137 : tmp22967;
  assign tmp23139 = s1 ? tmp22040 : tmp22797;
  assign tmp23140 = s1 ? tmp22954 : tmp21943;
  assign tmp23138 = s2 ? tmp23139 : tmp23140;
  assign tmp23135 = s3 ? tmp23136 : tmp23138;
  assign tmp23130 = s4 ? tmp23131 : tmp23135;
  assign tmp23119 = s5 ? tmp23120 : tmp23130;
  assign tmp23109 = s6 ? tmp23110 : tmp23119;
  assign tmp23145 = s2 ? tmp22992 : tmp23124;
  assign tmp23144 = s3 ? tmp22980 : tmp23145;
  assign tmp23147 = s2 ? tmp23127 : tmp22769;
  assign tmp23148 = s2 ? tmp22769 : tmp22269;
  assign tmp23146 = s3 ? tmp23147 : tmp23148;
  assign tmp23143 = s4 ? tmp23144 : tmp23146;
  assign tmp23152 = s1 ? tmp21943 : tmp22769;
  assign tmp23151 = s2 ? tmp21953 : tmp23152;
  assign tmp23150 = s3 ? tmp23132 : tmp23151;
  assign tmp23154 = s2 ? tmp21943 : tmp22769;
  assign tmp23155 = s2 ? tmp23152 : tmp21943;
  assign tmp23153 = s3 ? tmp23154 : tmp23155;
  assign tmp23149 = s4 ? tmp23150 : tmp23153;
  assign tmp23142 = s5 ? tmp23143 : tmp23149;
  assign tmp23141 = s6 ? tmp23110 : tmp23142;
  assign tmp23108 = s7 ? tmp23109 : tmp23141;
  assign tmp23163 = l1 ? 1 : tmp21964;
  assign tmp23162 = s0 ? tmp23163 : tmp22769;
  assign tmp23161 = s1 ? tmp22769 : tmp23162;
  assign tmp23160 = s2 ? tmp22269 : tmp23161;
  assign tmp23159 = s3 ? tmp23115 : tmp23160;
  assign tmp23158 = s4 ? tmp23111 : tmp23159;
  assign tmp23169 = s0 ? tmp23163 : 1;
  assign tmp23168 = s1 ? tmp23169 : tmp22769;
  assign tmp23167 = s2 ? tmp23123 : tmp23168;
  assign tmp23166 = s3 ? tmp22948 : tmp23167;
  assign tmp23165 = s4 ? tmp23166 : tmp23125;
  assign tmp23174 = s0 ? tmp21943 : tmp23163;
  assign tmp23173 = s1 ? tmp22800 : tmp23174;
  assign tmp23172 = s2 ? tmp23173 : tmp22967;
  assign tmp23171 = s3 ? tmp23172 : tmp23138;
  assign tmp23170 = s4 ? tmp23131 : tmp23171;
  assign tmp23164 = s5 ? tmp23165 : tmp23170;
  assign tmp23157 = s6 ? tmp23158 : tmp23164;
  assign tmp23179 = s2 ? tmp22992 : tmp23168;
  assign tmp23178 = s3 ? tmp22980 : tmp23179;
  assign tmp23177 = s4 ? tmp23178 : tmp23146;
  assign tmp23183 = s1 ? tmp21943 : tmp23174;
  assign tmp23182 = s2 ? tmp23183 : tmp22769;
  assign tmp23181 = s3 ? tmp23182 : tmp23155;
  assign tmp23180 = s4 ? tmp23150 : tmp23181;
  assign tmp23176 = s5 ? tmp23177 : tmp23180;
  assign tmp23175 = s6 ? tmp23158 : tmp23176;
  assign tmp23156 = s7 ? tmp23157 : tmp23175;
  assign tmp23107 = s8 ? tmp23108 : tmp23156;
  assign tmp23188 = s3 ? tmp22039 : tmp22599;
  assign tmp23190 = s2 ? tmp22054 : tmp21953;
  assign tmp23189 = s3 ? tmp23190 : tmp22617;
  assign tmp23187 = s4 ? tmp23188 : tmp23189;
  assign tmp23194 = s2 ? tmp22059 : tmp22053;
  assign tmp23195 = s2 ? tmp22603 : tmp22054;
  assign tmp23193 = s3 ? tmp23194 : tmp23195;
  assign tmp23197 = s2 ? tmp21953 : tmp22071;
  assign tmp23196 = s3 ? tmp23197 : tmp22070;
  assign tmp23192 = s4 ? tmp23193 : tmp23196;
  assign tmp23200 = s2 ? tmp22053 : tmp22060;
  assign tmp23199 = s3 ? tmp22472 : tmp23200;
  assign tmp23202 = s2 ? tmp21943 : tmp23017;
  assign tmp23203 = s2 ? tmp22040 : tmp21943;
  assign tmp23201 = s3 ? tmp23202 : tmp23203;
  assign tmp23198 = s4 ? tmp23199 : tmp23201;
  assign tmp23191 = s5 ? tmp23192 : tmp23198;
  assign tmp23186 = s6 ? tmp23187 : tmp23191;
  assign tmp23208 = s2 ? tmp22059 : tmp22206;
  assign tmp23209 = s2 ? tmp22269 : tmp22054;
  assign tmp23207 = s3 ? tmp23208 : tmp23209;
  assign tmp23211 = s2 ? tmp21953 : tmp21943;
  assign tmp23210 = s3 ? tmp23211 : tmp22268;
  assign tmp23206 = s4 ? tmp23207 : tmp23210;
  assign tmp23213 = s3 ? tmp22472 : tmp23211;
  assign tmp23212 = s4 ? tmp23213 : tmp21943;
  assign tmp23205 = s5 ? tmp23206 : tmp23212;
  assign tmp23204 = s6 ? tmp23187 : tmp23205;
  assign tmp23185 = s7 ? tmp23186 : tmp23204;
  assign tmp23184 = s8 ? tmp23156 : tmp23185;
  assign tmp23106 = s9 ? tmp23107 : tmp23184;
  assign tmp23221 = s2 ? tmp22769 : tmp22071;
  assign tmp23220 = s3 ? tmp23126 : tmp23221;
  assign tmp23219 = s4 ? tmp23121 : tmp23220;
  assign tmp23218 = s5 ? tmp23219 : tmp23130;
  assign tmp23217 = s6 ? tmp23110 : tmp23218;
  assign tmp23216 = s7 ? tmp23217 : tmp23141;
  assign tmp23215 = s8 ? tmp23216 : tmp23217;
  assign tmp23227 = s3 ? tmp23154 : tmp23152;
  assign tmp23226 = s4 ? tmp23150 : tmp23227;
  assign tmp23225 = s5 ? tmp23143 : tmp23226;
  assign tmp23224 = s6 ? tmp23110 : tmp23225;
  assign tmp23223 = s7 ? tmp23224 : tmp23204;
  assign tmp23232 = s3 ? tmp23182 : tmp23152;
  assign tmp23231 = s4 ? tmp23150 : tmp23232;
  assign tmp23230 = s5 ? tmp23177 : tmp23231;
  assign tmp23229 = s6 ? tmp23158 : tmp23230;
  assign tmp23228 = s7 ? tmp23229 : tmp23224;
  assign tmp23222 = s8 ? tmp23223 : tmp23228;
  assign tmp23214 = s9 ? tmp23215 : tmp23222;
  assign tmp23105 = s10 ? tmp23106 : tmp23214;
  assign tmp23236 = s7 ? tmp23141 : tmp23204;
  assign tmp23237 = s7 ? tmp23175 : tmp23141;
  assign tmp23235 = s8 ? tmp23236 : tmp23237;
  assign tmp23234 = s9 ? tmp23215 : tmp23235;
  assign tmp23233 = s10 ? tmp23106 : tmp23234;
  assign tmp23104 = ~(s11 ? tmp23105 : tmp23233);
  assign tmp23072 = ~(s12 ? tmp23073 : tmp23104);
  assign tmp22725 = s13 ? tmp22726 : tmp23072;
  assign tmp22590 = s14 ? tmp22591 : tmp22725;
  assign tmp21928 = s15 ? tmp21929 : tmp22590;
  assign tmp23249 = s3 ? tmp21996 : tmp22019;
  assign tmp23248 = s4 ? tmp22025 : tmp23249;
  assign tmp23247 = s5 ? tmp23248 : tmp21998;
  assign tmp23246 = s6 ? tmp22021 : tmp23247;
  assign tmp23245 = s7 ? tmp22004 : tmp23246;
  assign tmp23244 = s8 ? tmp21935 : tmp23245;
  assign tmp23255 = s3 ? tmp21943 : tmp22070;
  assign tmp23256 = s3 ? tmp22052 : tmp22472;
  assign tmp23254 = s4 ? tmp23255 : tmp23256;
  assign tmp23253 = s5 ? tmp23254 : tmp22056;
  assign tmp23252 = s6 ? tmp22035 : tmp23253;
  assign tmp23260 = s3 ? tmp22073 : tmp22472;
  assign tmp23259 = s4 ? tmp23255 : tmp23260;
  assign tmp23258 = s5 ? tmp23259 : tmp22075;
  assign tmp23257 = s6 ? tmp22064 : tmp23258;
  assign tmp23251 = s7 ? tmp23252 : tmp23257;
  assign tmp23250 = s8 ? tmp23245 : tmp23251;
  assign tmp23243 = s9 ? tmp23244 : tmp23250;
  assign tmp23262 = s8 ? tmp23245 : tmp22004;
  assign tmp23264 = s7 ? tmp22089 : tmp23257;
  assign tmp23268 = s3 ? tmp22093 : tmp22019;
  assign tmp23267 = s4 ? tmp22025 : tmp23268;
  assign tmp23266 = s5 ? tmp23267 : tmp21998;
  assign tmp23265 = s6 ? tmp22021 : tmp23266;
  assign tmp23263 = s8 ? tmp23264 : tmp23265;
  assign tmp23261 = s9 ? tmp23262 : tmp23263;
  assign tmp23242 = s10 ? tmp23243 : tmp23261;
  assign tmp23272 = s7 ? tmp21984 : tmp23257;
  assign tmp23271 = s8 ? tmp23272 : tmp23246;
  assign tmp23270 = s9 ? tmp23262 : tmp23271;
  assign tmp23269 = s10 ? tmp23243 : tmp23270;
  assign tmp23241 = s11 ? tmp23242 : tmp23269;
  assign tmp23283 = s1 ? tmp22046 : tmp22040;
  assign tmp23282 = s2 ? tmp22206 : tmp23283;
  assign tmp23281 = s3 ? tmp21943 : tmp23282;
  assign tmp23280 = s4 ? tmp21943 : tmp23281;
  assign tmp23287 = ~(s2 ? tmp22213 : 0);
  assign tmp23286 = s3 ? tmp22115 : tmp23287;
  assign tmp23285 = s4 ? tmp23286 : 1;
  assign tmp23284 = s5 ? tmp23285 : 1;
  assign tmp23279 = s6 ? tmp23280 : tmp23284;
  assign tmp23292 = ~(s2 ? tmp22225 : 0);
  assign tmp23291 = s3 ? tmp22224 : tmp23292;
  assign tmp23290 = s4 ? tmp23291 : 1;
  assign tmp23289 = s5 ? tmp23290 : 1;
  assign tmp23288 = s6 ? tmp23280 : tmp23289;
  assign tmp23278 = s7 ? tmp23279 : tmp23288;
  assign tmp23297 = s2 ? tmp22206 : tmp22039;
  assign tmp23296 = s3 ? tmp21943 : tmp23297;
  assign tmp23295 = s4 ? tmp21943 : tmp23296;
  assign tmp23300 = s3 ? tmp22066 : tmp22611;
  assign tmp23299 = s4 ? tmp23300 : 1;
  assign tmp23298 = s5 ? tmp23299 : 1;
  assign tmp23294 = s6 ? tmp23295 : tmp23298;
  assign tmp23304 = s3 ? tmp22268 : tmp22074;
  assign tmp23303 = s4 ? tmp23304 : 1;
  assign tmp23302 = s5 ? tmp23303 : 1;
  assign tmp23301 = s6 ? tmp23295 : tmp23302;
  assign tmp23293 = s7 ? tmp23294 : tmp23301;
  assign tmp23277 = s8 ? tmp23278 : tmp23293;
  assign tmp23276 = s9 ? tmp23277 : tmp23293;
  assign tmp23306 = s8 ? tmp23293 : tmp23294;
  assign tmp23312 = s2 ? tmp21953 : tmp23283;
  assign tmp23311 = s3 ? tmp21943 : tmp23312;
  assign tmp23310 = s4 ? tmp21943 : tmp23311;
  assign tmp23309 = s6 ? tmp23310 : tmp23289;
  assign tmp23315 = s3 ? tmp21943 : tmp22038;
  assign tmp23314 = s4 ? tmp21943 : tmp23315;
  assign tmp23313 = s6 ? tmp23314 : tmp23302;
  assign tmp23308 = s7 ? tmp23309 : tmp23313;
  assign tmp23307 = s8 ? tmp23308 : tmp23313;
  assign tmp23305 = s9 ? tmp23306 : tmp23307;
  assign tmp23275 = s10 ? tmp23276 : tmp23305;
  assign tmp23319 = s7 ? tmp23288 : tmp23301;
  assign tmp23318 = s8 ? tmp23319 : tmp23301;
  assign tmp23317 = s9 ? tmp23306 : tmp23318;
  assign tmp23316 = s10 ? tmp23276 : tmp23317;
  assign tmp23274 = s11 ? tmp23275 : tmp23316;
  assign tmp23273 = s12 ? tmp22101 : tmp23274;
  assign tmp23240 = s13 ? tmp23241 : tmp23273;
  assign tmp23332 = ~(s1 ? tmp22048 : tmp22049);
  assign tmp23331 = s2 ? tmp22110 : tmp23332;
  assign tmp23333 = s2 ? tmp22045 : tmp22396;
  assign tmp23330 = s3 ? tmp23331 : tmp23333;
  assign tmp23335 = s2 ? tmp22122 : 1;
  assign tmp23334 = ~(s3 ? tmp22167 : tmp23335);
  assign tmp23329 = s4 ? tmp23330 : tmp23334;
  assign tmp23328 = s5 ? tmp23329 : 0;
  assign tmp23327 = s6 ? tmp22131 : tmp23328;
  assign tmp23340 = s2 ? tmp22450 : tmp21943;
  assign tmp23339 = s3 ? tmp23340 : tmp23333;
  assign tmp23341 = ~(s3 ? tmp22167 : tmp23085);
  assign tmp23338 = s4 ? tmp23339 : tmp23341;
  assign tmp23337 = s5 ? tmp23338 : 0;
  assign tmp23336 = s6 ? tmp22150 : tmp23337;
  assign tmp23326 = ~(s7 ? tmp23327 : tmp23336);
  assign tmp23325 = s8 ? 1 : tmp23326;
  assign tmp23324 = s9 ? tmp23325 : tmp23326;
  assign tmp23344 = s7 ? tmp23327 : tmp23336;
  assign tmp23343 = s8 ? tmp23344 : tmp23327;
  assign tmp23351 = s2 ? tmp22116 : tmp22396;
  assign tmp23350 = s3 ? tmp23340 : tmp23351;
  assign tmp23349 = s4 ? tmp23350 : tmp23341;
  assign tmp23348 = s5 ? tmp23349 : 0;
  assign tmp23347 = ~(s6 ? tmp22150 : tmp23348);
  assign tmp23346 = s7 ? 1 : tmp23347;
  assign tmp23345 = ~(s8 ? tmp23346 : tmp23347);
  assign tmp23342 = ~(s9 ? tmp23343 : tmp23345);
  assign tmp23323 = s10 ? tmp23324 : tmp23342;
  assign tmp23356 = ~(s6 ? tmp22150 : tmp23337);
  assign tmp23355 = s7 ? 1 : tmp23356;
  assign tmp23354 = ~(s8 ? tmp23355 : tmp23356);
  assign tmp23353 = ~(s9 ? tmp23343 : tmp23354);
  assign tmp23352 = s10 ? tmp23324 : tmp23353;
  assign tmp23322 = s11 ? tmp23323 : tmp23352;
  assign tmp23364 = s4 ? tmp22379 : tmp22358;
  assign tmp23363 = s5 ? tmp23364 : tmp22361;
  assign tmp23362 = s6 ? tmp22349 : tmp23363;
  assign tmp23361 = s7 ? tmp22368 : tmp23362;
  assign tmp23369 = s2 ? tmp23039 : tmp21949;
  assign tmp23370 = s2 ? tmp22322 : tmp22895;
  assign tmp23368 = s3 ? tmp23369 : tmp23370;
  assign tmp23367 = s4 ? tmp21938 : tmp23368;
  assign tmp23375 = s1 ? tmp21950 : tmp21956;
  assign tmp23376 = s1 ? tmp21956 : tmp21946;
  assign tmp23374 = s2 ? tmp23375 : tmp23376;
  assign tmp23378 = ~(s1 ? 1 : tmp22869);
  assign tmp23377 = s2 ? tmp22015 : tmp23378;
  assign tmp23373 = s3 ? tmp23374 : tmp23377;
  assign tmp23381 = s1 ? tmp22868 : tmp22049;
  assign tmp23382 = ~(s1 ? tmp21943 : tmp21950);
  assign tmp23380 = s2 ? tmp23381 : tmp23382;
  assign tmp23385 = s0 ? tmp21964 : tmp22869;
  assign tmp23384 = s1 ? tmp23385 : tmp22315;
  assign tmp23383 = s2 ? tmp23384 : 1;
  assign tmp23379 = ~(s3 ? tmp23380 : tmp23383);
  assign tmp23372 = s4 ? tmp23373 : tmp23379;
  assign tmp23389 = s1 ? tmp21966 : tmp21964;
  assign tmp23388 = s2 ? tmp22338 : tmp23389;
  assign tmp23387 = s3 ? tmp23388 : tmp22340;
  assign tmp23390 = s3 ? tmp23388 : tmp22345;
  assign tmp23386 = ~(s4 ? tmp23387 : tmp23390);
  assign tmp23371 = s5 ? tmp23372 : tmp23386;
  assign tmp23366 = s6 ? tmp23367 : tmp23371;
  assign tmp23394 = s2 ? tmp23039 : tmp21988;
  assign tmp23395 = s2 ? tmp22116 : tmp22895;
  assign tmp23393 = s3 ? tmp23394 : tmp23395;
  assign tmp23392 = s4 ? tmp21938 : tmp23393;
  assign tmp23399 = s2 ? tmp23039 : tmp22027;
  assign tmp23400 = s2 ? tmp22029 : tmp23378;
  assign tmp23398 = s3 ? tmp23399 : tmp23400;
  assign tmp23403 = ~(s1 ? tmp21943 : tmp21940);
  assign tmp23402 = s2 ? tmp23381 : tmp23403;
  assign tmp23401 = ~(s3 ? tmp23402 : tmp23383);
  assign tmp23397 = s4 ? tmp23398 : tmp23401;
  assign tmp23406 = s2 ? tmp22338 : tmp21973;
  assign tmp23405 = s3 ? tmp23406 : tmp22364;
  assign tmp23404 = ~(s4 ? tmp23405 : tmp22365);
  assign tmp23396 = s5 ? tmp23397 : tmp23404;
  assign tmp23391 = s6 ? tmp23392 : tmp23396;
  assign tmp23365 = ~(s7 ? tmp23366 : tmp23391);
  assign tmp23360 = s8 ? tmp23361 : tmp23365;
  assign tmp23408 = s7 ? tmp23366 : tmp23391;
  assign tmp23411 = s4 ? tmp21943 : tmp22390;
  assign tmp23415 = s2 ? tmp23014 : tmp22060;
  assign tmp23414 = s3 ? tmp23415 : tmp22395;
  assign tmp23413 = s4 ? tmp23414 : tmp22397;
  assign tmp23418 = s2 ? tmp22210 : tmp23332;
  assign tmp23417 = s3 ? tmp23418 : tmp22402;
  assign tmp23419 = s3 ? tmp23418 : tmp22407;
  assign tmp23416 = s4 ? tmp23417 : tmp23419;
  assign tmp23412 = s5 ? tmp23413 : tmp23416;
  assign tmp23410 = s6 ? tmp23411 : tmp23412;
  assign tmp23421 = s4 ? tmp21943 : tmp22411;
  assign tmp23425 = s2 ? tmp22054 : tmp21943;
  assign tmp23424 = s3 ? tmp23425 : tmp22395;
  assign tmp23423 = s4 ? tmp23424 : tmp22397;
  assign tmp23427 = s3 ? tmp22234 : tmp22419;
  assign tmp23426 = s4 ? tmp23427 : tmp22420;
  assign tmp23422 = s5 ? tmp23423 : tmp23426;
  assign tmp23420 = s6 ? tmp23421 : tmp23422;
  assign tmp23409 = s7 ? tmp23410 : tmp23420;
  assign tmp23407 = ~(s8 ? tmp23408 : tmp23409);
  assign tmp23359 = s9 ? tmp23360 : tmp23407;
  assign tmp23429 = s8 ? tmp23408 : tmp23366;
  assign tmp23434 = s4 ? tmp22379 : tmp22433;
  assign tmp23433 = s5 ? tmp23434 : tmp22361;
  assign tmp23432 = s6 ? tmp22349 : tmp23433;
  assign tmp23435 = ~(s6 ? tmp23421 : tmp23422);
  assign tmp23431 = s7 ? tmp23432 : tmp23435;
  assign tmp23441 = s1 ? tmp23385 : tmp21964;
  assign tmp23440 = s2 ? tmp23441 : 1;
  assign tmp23439 = ~(s3 ? tmp23402 : tmp23440);
  assign tmp23438 = s4 ? tmp23398 : tmp23439;
  assign tmp23437 = s5 ? tmp23438 : tmp23404;
  assign tmp23436 = ~(s6 ? tmp23392 : tmp23437);
  assign tmp23430 = ~(s8 ? tmp23431 : tmp23436);
  assign tmp23428 = ~(s9 ? tmp23429 : tmp23430);
  assign tmp23358 = s10 ? tmp23359 : tmp23428;
  assign tmp23445 = s7 ? tmp23362 : tmp23435;
  assign tmp23446 = ~(s6 ? tmp23392 : tmp23396);
  assign tmp23444 = ~(s8 ? tmp23445 : tmp23446);
  assign tmp23443 = ~(s9 ? tmp23429 : tmp23444);
  assign tmp23442 = s10 ? tmp23359 : tmp23443;
  assign tmp23357 = s11 ? tmp23358 : tmp23442;
  assign tmp23321 = s12 ? tmp23322 : tmp23357;
  assign tmp23454 = s2 ? tmp21940 : tmp22872;
  assign tmp23453 = s3 ? tmp21939 : tmp23454;
  assign tmp23457 = s1 ? tmp22873 : tmp22046;
  assign tmp23456 = s2 ? tmp21945 : tmp23457;
  assign tmp23458 = s2 ? tmp22454 : tmp22008;
  assign tmp23455 = s3 ? tmp23456 : tmp23458;
  assign tmp23452 = s4 ? tmp23453 : tmp23455;
  assign tmp23463 = s1 ? tmp22873 : tmp22896;
  assign tmp23465 = ~(s0 ? tmp21940 : 0);
  assign tmp23464 = ~(s1 ? tmp22868 : tmp23465);
  assign tmp23462 = s2 ? tmp23463 : tmp23464;
  assign tmp23467 = ~(s1 ? 1 : tmp21940);
  assign tmp23466 = ~(s2 ? tmp22868 : tmp23467);
  assign tmp23461 = s3 ? tmp23462 : tmp23466;
  assign tmp23470 = s1 ? tmp21956 : tmp21943;
  assign tmp23469 = s2 ? tmp23470 : tmp21997;
  assign tmp23472 = s1 ? tmp21940 : 1;
  assign tmp23471 = s2 ? tmp23472 : 1;
  assign tmp23468 = s3 ? tmp23469 : tmp23471;
  assign tmp23460 = s4 ? tmp23461 : tmp23468;
  assign tmp23475 = s2 ? tmp23472 : tmp22871;
  assign tmp23474 = s3 ? tmp23475 : 1;
  assign tmp23477 = s2 ? 1 : tmp21940;
  assign tmp23476 = s3 ? tmp23477 : 1;
  assign tmp23473 = s4 ? tmp23474 : tmp23476;
  assign tmp23459 = s5 ? tmp23460 : tmp23473;
  assign tmp23451 = s6 ? tmp23452 : tmp23459;
  assign tmp23482 = s1 ? tmp22873 : tmp21943;
  assign tmp23481 = s2 ? tmp21945 : tmp23482;
  assign tmp23480 = s3 ? tmp23481 : tmp22007;
  assign tmp23479 = s4 ? tmp23453 : tmp23480;
  assign tmp23486 = s2 ? tmp22872 : tmp22917;
  assign tmp23487 = s2 ? tmp21940 : tmp22993;
  assign tmp23485 = s3 ? tmp23486 : tmp23487;
  assign tmp23489 = s2 ? tmp23470 : tmp21940;
  assign tmp23488 = s3 ? tmp23489 : tmp23471;
  assign tmp23484 = s4 ? tmp23485 : tmp23488;
  assign tmp23491 = s3 ? tmp23472 : 1;
  assign tmp23490 = s4 ? tmp23491 : tmp23476;
  assign tmp23483 = s5 ? tmp23484 : tmp23490;
  assign tmp23478 = s6 ? tmp23479 : tmp23483;
  assign tmp23450 = s7 ? tmp23451 : tmp23478;
  assign tmp23497 = s2 ? tmp22454 : tmp21943;
  assign tmp23496 = s3 ? tmp22452 : tmp23497;
  assign tmp23495 = s4 ? tmp22448 : tmp23496;
  assign tmp23501 = ~(s2 ? tmp22048 : tmp22144);
  assign tmp23500 = s3 ? tmp22458 : tmp23501;
  assign tmp23502 = s3 ? tmp22462 : tmp22611;
  assign tmp23499 = s4 ? tmp23500 : tmp23502;
  assign tmp23504 = s3 ? tmp21943 : 1;
  assign tmp23505 = s3 ? tmp22617 : tmp22074;
  assign tmp23503 = s4 ? tmp23504 : tmp23505;
  assign tmp23498 = s5 ? tmp23499 : tmp23503;
  assign tmp23494 = s6 ? tmp23495 : tmp23498;
  assign tmp23508 = s3 ? tmp22452 : tmp23211;
  assign tmp23507 = s4 ? tmp22448 : tmp23508;
  assign tmp23511 = s3 ? tmp22469 : tmp22066;
  assign tmp23510 = s4 ? tmp23511 : tmp22461;
  assign tmp23509 = s5 ? tmp23510 : tmp23504;
  assign tmp23506 = s6 ? tmp23507 : tmp23509;
  assign tmp23493 = s7 ? tmp23494 : tmp23506;
  assign tmp23492 = s8 ? tmp23450 : tmp23493;
  assign tmp23449 = s9 ? tmp23450 : tmp23492;
  assign tmp23518 = s2 ? tmp22454 : tmp21939;
  assign tmp23517 = s3 ? tmp23456 : tmp23518;
  assign tmp23516 = s4 ? tmp23453 : tmp23517;
  assign tmp23521 = s3 ? tmp23462 : tmp22887;
  assign tmp23524 = s1 ? tmp21940 : tmp21951;
  assign tmp23523 = s2 ? tmp23524 : 1;
  assign tmp23522 = s3 ? tmp23469 : tmp23523;
  assign tmp23520 = s4 ? tmp23521 : tmp23522;
  assign tmp23528 = s1 ? tmp21940 : tmp21943;
  assign tmp23529 = s1 ? tmp21942 : tmp21940;
  assign tmp23527 = s2 ? tmp23528 : tmp23529;
  assign tmp23526 = s3 ? tmp23527 : 1;
  assign tmp23531 = s2 ? tmp22269 : tmp21940;
  assign tmp23530 = s3 ? tmp23531 : tmp22074;
  assign tmp23525 = s4 ? tmp23526 : tmp23530;
  assign tmp23519 = s5 ? tmp23520 : tmp23525;
  assign tmp23515 = s6 ? tmp23516 : tmp23519;
  assign tmp23535 = s2 ? tmp21953 : tmp21939;
  assign tmp23534 = s3 ? tmp23481 : tmp23535;
  assign tmp23533 = s4 ? tmp23453 : tmp23534;
  assign tmp23538 = s3 ? tmp23486 : tmp22918;
  assign tmp23537 = s4 ? tmp23538 : tmp23488;
  assign tmp23541 = s2 ? tmp23528 : tmp23472;
  assign tmp23540 = s3 ? tmp23541 : 1;
  assign tmp23542 = s3 ? tmp22928 : 1;
  assign tmp23539 = s4 ? tmp23540 : tmp23542;
  assign tmp23536 = s5 ? tmp23537 : tmp23539;
  assign tmp23532 = s6 ? tmp23533 : tmp23536;
  assign tmp23514 = s7 ? tmp23515 : tmp23532;
  assign tmp23513 = s8 ? tmp23514 : tmp23515;
  assign tmp23544 = s7 ? tmp23478 : tmp23506;
  assign tmp23543 = s8 ? tmp23544 : tmp23532;
  assign tmp23512 = s9 ? tmp23513 : tmp23543;
  assign tmp23448 = s10 ? tmp23449 : tmp23512;
  assign tmp23447 = ~(s12 ? tmp23448 : 1);
  assign tmp23320 = ~(s13 ? tmp23321 : tmp23447);
  assign tmp23239 = s14 ? tmp23240 : tmp23320;
  assign tmp23559 = ~(l4 ? 1 : 0);
  assign tmp23558 = ~(l2 ? 1 : tmp23559);
  assign tmp23557 = l1 ? 1 : tmp23558;
  assign tmp23560 = s0 ? tmp21943 : tmp23557;
  assign tmp23556 = s1 ? tmp23557 : tmp23560;
  assign tmp23562 = s1 ? tmp21950 : tmp23557;
  assign tmp23561 = s2 ? tmp23557 : tmp23562;
  assign tmp23555 = s3 ? tmp23556 : tmp23561;
  assign tmp23566 = s0 ? tmp23557 : 1;
  assign tmp23565 = s1 ? tmp23566 : tmp23557;
  assign tmp23567 = s1 ? tmp23566 : tmp21951;
  assign tmp23564 = s2 ? tmp23565 : tmp23567;
  assign tmp23568 = s2 ? tmp22322 : tmp23556;
  assign tmp23563 = s3 ? tmp23564 : tmp23568;
  assign tmp23554 = s4 ? tmp23555 : tmp23563;
  assign tmp23573 = s1 ? tmp23566 : 1;
  assign tmp23575 = s0 ? 1 : tmp23557;
  assign tmp23574 = s1 ? tmp23575 : tmp23557;
  assign tmp23572 = s2 ? tmp23573 : tmp23574;
  assign tmp23577 = s1 ? tmp22046 : tmp23557;
  assign tmp23576 = s2 ? tmp23557 : tmp23577;
  assign tmp23571 = s3 ? tmp23572 : tmp23576;
  assign tmp23582 = ~(l1 ? 1 : tmp23558);
  assign tmp23581 = s0 ? 1 : tmp23582;
  assign tmp23580 = s1 ? tmp23581 : tmp22049;
  assign tmp23583 = ~(s1 ? tmp21943 : tmp23566);
  assign tmp23579 = s2 ? tmp23580 : tmp23583;
  assign tmp23584 = ~(s2 ? tmp23556 : 0);
  assign tmp23578 = ~(s3 ? tmp23579 : tmp23584);
  assign tmp23570 = s4 ? tmp23571 : tmp23578;
  assign tmp23589 = s0 ? tmp23557 : 0;
  assign tmp23588 = s1 ? tmp23589 : tmp22111;
  assign tmp23587 = s2 ? tmp23588 : tmp22059;
  assign tmp23591 = ~(s1 ? 1 : tmp23581);
  assign tmp23590 = s2 ? tmp22255 : tmp23591;
  assign tmp23586 = s3 ? tmp23587 : tmp23590;
  assign tmp23595 = s0 ? tmp23557 : tmp21943;
  assign tmp23594 = s1 ? tmp23595 : tmp21943;
  assign tmp23596 = ~(s1 ? tmp23581 : 0);
  assign tmp23593 = s2 ? tmp23594 : tmp23596;
  assign tmp23599 = ~(s0 ? 1 : tmp23582);
  assign tmp23598 = s1 ? tmp21943 : tmp23599;
  assign tmp23600 = ~(s1 ? tmp23581 : tmp22048);
  assign tmp23597 = s2 ? tmp23598 : tmp23600;
  assign tmp23592 = s3 ? tmp23593 : tmp23597;
  assign tmp23585 = s4 ? tmp23586 : tmp23592;
  assign tmp23569 = s5 ? tmp23570 : tmp23585;
  assign tmp23553 = s6 ? tmp23554 : tmp23569;
  assign tmp23605 = s1 ? tmp23566 : tmp21943;
  assign tmp23604 = s2 ? tmp23565 : tmp23605;
  assign tmp23606 = s2 ? tmp22116 : tmp23556;
  assign tmp23603 = s3 ? tmp23604 : tmp23606;
  assign tmp23602 = s4 ? tmp23555 : tmp23603;
  assign tmp23610 = s2 ? tmp23573 : tmp23557;
  assign tmp23609 = s3 ? tmp23610 : tmp23576;
  assign tmp23613 = ~(s1 ? tmp21943 : tmp23557);
  assign tmp23612 = s2 ? tmp23580 : tmp23613;
  assign tmp23611 = ~(s3 ? tmp23612 : tmp23584);
  assign tmp23608 = s4 ? tmp23609 : tmp23611;
  assign tmp23617 = s1 ? tmp23589 : tmp21943;
  assign tmp23616 = s2 ? tmp23617 : 1;
  assign tmp23619 = s1 ? 1 : tmp23582;
  assign tmp23618 = ~(s2 ? 1 : tmp23619);
  assign tmp23615 = s3 ? tmp23616 : tmp23618;
  assign tmp23621 = s2 ? tmp21943 : tmp23557;
  assign tmp23622 = s1 ? tmp21943 : tmp23557;
  assign tmp23620 = s3 ? tmp23621 : tmp23622;
  assign tmp23614 = s4 ? tmp23615 : tmp23620;
  assign tmp23607 = s5 ? tmp23608 : tmp23614;
  assign tmp23601 = s6 ? tmp23602 : tmp23607;
  assign tmp23552 = s7 ? tmp23553 : tmp23601;
  assign tmp23626 = s3 ? tmp22769 : tmp22982;
  assign tmp23628 = s2 ? tmp22937 : tmp22772;
  assign tmp23631 = s0 ? tmp22765 : tmp22769;
  assign tmp23630 = s1 ? tmp22769 : tmp23631;
  assign tmp23629 = s2 ? tmp22779 : tmp23630;
  assign tmp23627 = s3 ? tmp23628 : tmp23629;
  assign tmp23625 = s4 ? tmp23626 : tmp23627;
  assign tmp23635 = s2 ? tmp22797 : tmp22835;
  assign tmp23634 = s3 ? tmp22948 : tmp23635;
  assign tmp23639 = s0 ? 1 : tmp22806;
  assign tmp23638 = s1 ? tmp23639 : tmp22795;
  assign tmp23640 = ~(s1 ? tmp22797 : tmp22772);
  assign tmp23637 = s2 ? tmp23638 : tmp23640;
  assign tmp23643 = s0 ? tmp22769 : tmp23557;
  assign tmp23642 = s1 ? tmp22769 : tmp23643;
  assign tmp23641 = ~(s2 ? tmp23642 : 0);
  assign tmp23636 = ~(s3 ? tmp23637 : tmp23641);
  assign tmp23633 = s4 ? tmp23634 : tmp23636;
  assign tmp23647 = s1 ? tmp22941 : tmp22805;
  assign tmp23646 = s2 ? tmp23647 : tmp22807;
  assign tmp23645 = s3 ? tmp23646 : tmp23590;
  assign tmp23650 = s1 ? tmp23595 : tmp22811;
  assign tmp23651 = ~(s1 ? tmp23639 : 0);
  assign tmp23649 = s2 ? tmp23650 : tmp23651;
  assign tmp23653 = s1 ? tmp22800 : tmp23599;
  assign tmp23652 = s2 ? tmp23653 : tmp23600;
  assign tmp23648 = s3 ? tmp23649 : tmp23652;
  assign tmp23644 = s4 ? tmp23645 : tmp23648;
  assign tmp23632 = s5 ? tmp23633 : tmp23644;
  assign tmp23624 = s6 ? tmp23625 : tmp23632;
  assign tmp23657 = s2 ? tmp22821 : tmp23630;
  assign tmp23656 = s3 ? tmp22937 : tmp23657;
  assign tmp23655 = s4 ? tmp23626 : tmp23656;
  assign tmp23661 = s2 ? tmp22769 : tmp22835;
  assign tmp23660 = s3 ? tmp22980 : tmp23661;
  assign tmp23663 = s2 ? tmp23638 : tmp22806;
  assign tmp23665 = s1 ? tmp22769 : tmp23557;
  assign tmp23664 = ~(s2 ? tmp23665 : 0);
  assign tmp23662 = ~(s3 ? tmp23663 : tmp23664);
  assign tmp23659 = s4 ? tmp23660 : tmp23662;
  assign tmp23669 = s1 ? tmp22941 : tmp22769;
  assign tmp23668 = s2 ? tmp23669 : 1;
  assign tmp23667 = s3 ? tmp23668 : tmp23618;
  assign tmp23671 = s2 ? tmp22838 : tmp22769;
  assign tmp23670 = s3 ? tmp23671 : tmp23622;
  assign tmp23666 = s4 ? tmp23667 : tmp23670;
  assign tmp23658 = s5 ? tmp23659 : tmp23666;
  assign tmp23654 = s6 ? tmp23655 : tmp23658;
  assign tmp23623 = s7 ? tmp23624 : tmp23654;
  assign tmp23551 = s8 ? tmp23552 : tmp23623;
  assign tmp23672 = s8 ? tmp23623 : tmp22840;
  assign tmp23550 = s9 ? tmp23551 : tmp23672;
  assign tmp23680 = s2 ? tmp23580 : tmp23582;
  assign tmp23681 = ~(s2 ? tmp23557 : 0);
  assign tmp23679 = ~(s3 ? tmp23680 : tmp23681);
  assign tmp23678 = s4 ? tmp23609 : tmp23679;
  assign tmp23677 = s5 ? tmp23678 : tmp23614;
  assign tmp23676 = s6 ? tmp23602 : tmp23677;
  assign tmp23675 = s7 ? tmp23553 : tmp23676;
  assign tmp23674 = s8 ? tmp23675 : tmp23553;
  assign tmp23687 = ~(s3 ? tmp23612 : tmp23681);
  assign tmp23686 = s4 ? tmp23609 : tmp23687;
  assign tmp23685 = s5 ? tmp23686 : tmp23614;
  assign tmp23684 = s6 ? tmp23602 : tmp23685;
  assign tmp23683 = s7 ? tmp23684 : tmp22841;
  assign tmp23688 = s7 ? tmp23654 : tmp23676;
  assign tmp23682 = s8 ? tmp23683 : tmp23688;
  assign tmp23673 = s9 ? tmp23674 : tmp23682;
  assign tmp23549 = s10 ? tmp23550 : tmp23673;
  assign tmp23692 = s7 ? tmp23601 : tmp22841;
  assign tmp23691 = s8 ? tmp23692 : tmp23688;
  assign tmp23690 = s9 ? tmp23674 : tmp23691;
  assign tmp23689 = s10 ? tmp23550 : tmp23690;
  assign tmp23548 = s11 ? tmp23549 : tmp23689;
  assign tmp23700 = s2 ? tmp22872 : tmp22878;
  assign tmp23699 = ~(s3 ? tmp23700 : tmp22879);
  assign tmp23698 = s4 ? tmp22867 : tmp23699;
  assign tmp23704 = s2 ? tmp23472 : tmp22917;
  assign tmp23703 = s3 ? tmp23704 : tmp22887;
  assign tmp23707 = s1 ? tmp21942 : 0;
  assign tmp23708 = ~(s1 ? 1 : tmp23465);
  assign tmp23706 = s2 ? tmp23707 : tmp23708;
  assign tmp23705 = s3 ? tmp23706 : tmp22894;
  assign tmp23702 = s4 ? tmp23703 : tmp23705;
  assign tmp23701 = ~(s5 ? tmp23702 : tmp22897);
  assign tmp23697 = s6 ? tmp23698 : tmp23701;
  assign tmp23711 = ~(s3 ? tmp23700 : tmp22912);
  assign tmp23710 = s4 ? tmp22867 : tmp23711;
  assign tmp23714 = s3 ? tmp23704 : tmp22918;
  assign tmp23716 = s2 ? tmp23707 : tmp21940;
  assign tmp23715 = s3 ? tmp23716 : tmp22922;
  assign tmp23713 = s4 ? tmp23714 : tmp23715;
  assign tmp23712 = ~(s5 ? tmp23713 : tmp22923);
  assign tmp23709 = s6 ? tmp23710 : tmp23712;
  assign tmp23696 = s7 ? tmp23697 : tmp23709;
  assign tmp23722 = s2 ? tmp21940 : tmp22878;
  assign tmp23721 = ~(s3 ? tmp23722 : tmp22879);
  assign tmp23720 = s4 ? tmp23035 : tmp23721;
  assign tmp23726 = s2 ? tmp23472 : tmp21940;
  assign tmp23725 = s3 ? tmp23726 : tmp22918;
  assign tmp23728 = s2 ? tmp23707 : tmp23378;
  assign tmp23727 = s3 ? tmp23728 : tmp22894;
  assign tmp23724 = s4 ? tmp23725 : tmp23727;
  assign tmp23723 = ~(s5 ? tmp23724 : tmp22897);
  assign tmp23719 = s6 ? tmp23720 : tmp23723;
  assign tmp23731 = ~(s3 ? tmp23722 : tmp22912);
  assign tmp23730 = s4 ? tmp23035 : tmp23731;
  assign tmp23733 = s4 ? tmp23725 : tmp23715;
  assign tmp23732 = ~(s5 ? tmp23733 : tmp22923);
  assign tmp23729 = s6 ? tmp23730 : tmp23732;
  assign tmp23718 = s7 ? tmp23719 : tmp23729;
  assign tmp23738 = ~(s2 ? tmp21943 : tmp22450);
  assign tmp23737 = s3 ? tmp22048 : tmp23738;
  assign tmp23740 = s2 ? tmp21943 : tmp22210;
  assign tmp23739 = ~(s3 ? tmp23740 : tmp23003);
  assign tmp23736 = s4 ? tmp23737 : tmp23739;
  assign tmp23743 = s3 ? tmp22044 : tmp23501;
  assign tmp23744 = s3 ? tmp23351 : tmp23010;
  assign tmp23742 = s4 ? tmp23743 : tmp23744;
  assign tmp23747 = s2 ? tmp23014 : tmp21943;
  assign tmp23746 = s3 ? tmp23747 : tmp22079;
  assign tmp23749 = s2 ? tmp22054 : tmp22060;
  assign tmp23748 = s3 ? tmp23749 : tmp23018;
  assign tmp23745 = s4 ? tmp23746 : tmp23748;
  assign tmp23741 = ~(s5 ? tmp23742 : tmp23745);
  assign tmp23735 = s6 ? tmp23736 : tmp23741;
  assign tmp23752 = ~(s3 ? tmp23740 : tmp23022);
  assign tmp23751 = s4 ? tmp23737 : tmp23752;
  assign tmp23755 = s3 ? tmp22044 : tmp22066;
  assign tmp23756 = s3 ? tmp22752 : tmp22268;
  assign tmp23754 = s4 ? tmp23755 : tmp23756;
  assign tmp23758 = s3 ? tmp23190 : tmp22079;
  assign tmp23757 = s4 ? tmp23758 : tmp21943;
  assign tmp23753 = ~(s5 ? tmp23754 : tmp23757);
  assign tmp23750 = s6 ? tmp23751 : tmp23753;
  assign tmp23734 = s7 ? tmp23735 : tmp23750;
  assign tmp23717 = s8 ? tmp23718 : tmp23734;
  assign tmp23695 = s9 ? tmp23696 : tmp23717;
  assign tmp23765 = ~(s2 ? tmp21940 : tmp22872);
  assign tmp23764 = s3 ? tmp22868 : tmp23765;
  assign tmp23763 = s4 ? tmp23764 : tmp23721;
  assign tmp23769 = s2 ? tmp21940 : tmp22917;
  assign tmp23768 = s3 ? tmp23769 : tmp22887;
  assign tmp23767 = s4 ? tmp23768 : tmp23727;
  assign tmp23772 = s2 ? tmp22900 : tmp23529;
  assign tmp23771 = s3 ? tmp23772 : tmp22901;
  assign tmp23774 = s2 ? tmp21988 : tmp22871;
  assign tmp23773 = s3 ? tmp23774 : tmp22906;
  assign tmp23770 = s4 ? tmp23771 : tmp23773;
  assign tmp23766 = ~(s5 ? tmp23767 : tmp23770);
  assign tmp23762 = s6 ? tmp23763 : tmp23766;
  assign tmp23776 = s4 ? tmp23764 : tmp23731;
  assign tmp23779 = s3 ? tmp23769 : tmp22918;
  assign tmp23778 = s4 ? tmp23779 : tmp23715;
  assign tmp23782 = s2 ? tmp21988 : tmp22908;
  assign tmp23781 = s3 ? tmp23782 : tmp22926;
  assign tmp23780 = s4 ? tmp23781 : tmp22927;
  assign tmp23777 = ~(s5 ? tmp23778 : tmp23780);
  assign tmp23775 = s6 ? tmp23776 : tmp23777;
  assign tmp23761 = s7 ? tmp23762 : tmp23775;
  assign tmp23760 = s8 ? tmp23761 : tmp23762;
  assign tmp23786 = ~(s5 ? tmp23713 : tmp23065);
  assign tmp23785 = s6 ? tmp23710 : tmp23786;
  assign tmp23784 = s7 ? tmp23785 : tmp23750;
  assign tmp23789 = s4 ? tmp23781 : tmp23060;
  assign tmp23788 = ~(s5 ? tmp23778 : tmp23789);
  assign tmp23787 = s6 ? tmp23776 : tmp23788;
  assign tmp23783 = s8 ? tmp23784 : tmp23787;
  assign tmp23759 = s9 ? tmp23760 : tmp23783;
  assign tmp23694 = s10 ? tmp23695 : tmp23759;
  assign tmp23793 = s7 ? tmp23709 : tmp23750;
  assign tmp23792 = s8 ? tmp23793 : tmp23775;
  assign tmp23791 = s9 ? tmp23760 : tmp23792;
  assign tmp23790 = s10 ? tmp23695 : tmp23791;
  assign tmp23693 = ~(s11 ? tmp23694 : tmp23790);
  assign tmp23547 = s12 ? tmp23548 : tmp23693;
  assign tmp23546 = s13 ? tmp23547 : tmp23072;
  assign tmp23545 = s14 ? tmp22591 : tmp23546;
  assign tmp23238 = s15 ? tmp23239 : tmp23545;
  assign tmp21927 = s16 ? tmp21928 : tmp23238;
  assign tmp23801 = s8 ? tmp23245 : tmp22033;
  assign tmp23800 = s9 ? tmp23244 : tmp23801;
  assign tmp23804 = s7 ? tmp23265 : tmp22083;
  assign tmp23803 = s8 ? tmp22088 : tmp23804;
  assign tmp23802 = s9 ? tmp22081 : tmp23803;
  assign tmp23799 = s10 ? tmp23800 : tmp23802;
  assign tmp23808 = s7 ? tmp23246 : tmp22083;
  assign tmp23807 = s8 ? tmp22099 : tmp23808;
  assign tmp23806 = s9 ? tmp22081 : tmp23807;
  assign tmp23805 = s10 ? tmp23800 : tmp23806;
  assign tmp23798 = s11 ? tmp23799 : tmp23805;
  assign tmp23817 = s3 ? tmp22262 : tmp23312;
  assign tmp23816 = s4 ? tmp21943 : tmp23817;
  assign tmp23815 = s6 ? tmp23816 : tmp23289;
  assign tmp23814 = s7 ? tmp23279 : tmp23815;
  assign tmp23813 = s8 ? tmp23293 : tmp23814;
  assign tmp23812 = s9 ? tmp23277 : tmp23813;
  assign tmp23819 = s8 ? tmp23814 : tmp23279;
  assign tmp23821 = s7 ? tmp23309 : tmp23815;
  assign tmp23822 = s7 ? tmp23313 : tmp23815;
  assign tmp23820 = s8 ? tmp23821 : tmp23822;
  assign tmp23818 = s9 ? tmp23819 : tmp23820;
  assign tmp23811 = s10 ? tmp23812 : tmp23818;
  assign tmp23826 = s7 ? tmp23288 : tmp23815;
  assign tmp23827 = s7 ? tmp23301 : tmp23815;
  assign tmp23825 = s8 ? tmp23826 : tmp23827;
  assign tmp23824 = s9 ? tmp23819 : tmp23825;
  assign tmp23823 = s10 ? tmp23812 : tmp23824;
  assign tmp23810 = s11 ? tmp23811 : tmp23823;
  assign tmp23809 = s12 ? tmp22101 : tmp23810;
  assign tmp23797 = s13 ? tmp23798 : tmp23809;
  assign tmp23833 = ~(s8 ? tmp23344 : 0);
  assign tmp23832 = s9 ? tmp23325 : tmp23833;
  assign tmp23837 = s6 ? tmp22150 : tmp23348;
  assign tmp23836 = ~(s7 ? tmp23837 : 0);
  assign tmp23835 = s8 ? 1 : tmp23836;
  assign tmp23834 = s9 ? 1 : tmp23835;
  assign tmp23831 = s10 ? tmp23832 : tmp23834;
  assign tmp23841 = ~(s7 ? tmp23336 : 0);
  assign tmp23840 = s8 ? 1 : tmp23841;
  assign tmp23839 = s9 ? 1 : tmp23840;
  assign tmp23838 = s10 ? tmp23832 : tmp23839;
  assign tmp23830 = s11 ? tmp23831 : tmp23838;
  assign tmp23851 = s2 ? tmp22040 : tmp22396;
  assign tmp23850 = s3 ? tmp23194 : tmp23851;
  assign tmp23849 = s4 ? tmp23850 : tmp22397;
  assign tmp23848 = s5 ? tmp23849 : tmp22399;
  assign tmp23847 = s6 ? tmp22388 : tmp23848;
  assign tmp23855 = s3 ? tmp23208 : tmp22395;
  assign tmp23854 = s4 ? tmp23855 : tmp22397;
  assign tmp23853 = s5 ? tmp23854 : tmp22416;
  assign tmp23852 = s6 ? tmp22410 : tmp23853;
  assign tmp23846 = s7 ? tmp23847 : tmp23852;
  assign tmp23845 = ~(s8 ? tmp23408 : tmp23846);
  assign tmp23844 = s9 ? tmp23360 : tmp23845;
  assign tmp23857 = s8 ? tmp22367 : tmp22368;
  assign tmp23860 = ~(s6 ? tmp22410 : tmp23853);
  assign tmp23859 = s7 ? tmp23432 : tmp23860;
  assign tmp23862 = s6 ? tmp23392 : tmp23437;
  assign tmp23863 = ~(s6 ? tmp22349 : tmp22377);
  assign tmp23861 = ~(s7 ? tmp23862 : tmp23863);
  assign tmp23858 = s8 ? tmp23859 : tmp23861;
  assign tmp23856 = s9 ? tmp23857 : tmp23858;
  assign tmp23843 = s10 ? tmp23844 : tmp23856;
  assign tmp23867 = s7 ? tmp23362 : tmp23860;
  assign tmp23868 = ~(s7 ? tmp23391 : tmp23863);
  assign tmp23866 = s8 ? tmp23867 : tmp23868;
  assign tmp23865 = s9 ? tmp23857 : tmp23866;
  assign tmp23864 = s10 ? tmp23844 : tmp23865;
  assign tmp23842 = s11 ? tmp23843 : tmp23864;
  assign tmp23829 = s12 ? tmp23830 : tmp23842;
  assign tmp23876 = s3 ? tmp21943 : tmp22074;
  assign tmp23875 = s4 ? tmp22457 : tmp23876;
  assign tmp23879 = s2 ? tmp21953 : tmp22060;
  assign tmp23878 = s3 ? tmp23879 : 1;
  assign tmp23877 = s4 ? tmp23878 : tmp22078;
  assign tmp23874 = s5 ? tmp23875 : tmp23877;
  assign tmp23873 = s6 ? tmp22447 : tmp23874;
  assign tmp23882 = s4 ? tmp22468 : tmp23876;
  assign tmp23884 = s3 ? tmp23211 : tmp22472;
  assign tmp23883 = s4 ? tmp23884 : tmp22078;
  assign tmp23881 = s5 ? tmp23882 : tmp23883;
  assign tmp23880 = s6 ? tmp22464 : tmp23881;
  assign tmp23872 = s7 ? tmp23873 : tmp23880;
  assign tmp23890 = s3 ? tmp21953 : 1;
  assign tmp23889 = s4 ? tmp23890 : tmp22078;
  assign tmp23888 = s5 ? tmp23882 : tmp23889;
  assign tmp23887 = s6 ? tmp22464 : tmp23888;
  assign tmp23886 = s7 ? tmp23873 : tmp23887;
  assign tmp23885 = s8 ? tmp23872 : tmp23886;
  assign tmp23871 = s9 ? tmp23872 : tmp23885;
  assign tmp23897 = s3 ? tmp21953 : tmp22472;
  assign tmp23896 = s4 ? tmp23897 : tmp22078;
  assign tmp23895 = s5 ? tmp23882 : tmp23896;
  assign tmp23894 = s6 ? tmp22464 : tmp23895;
  assign tmp23893 = s7 ? tmp23873 : tmp23894;
  assign tmp23892 = s8 ? tmp23893 : tmp23873;
  assign tmp23898 = s7 ? tmp23880 : tmp23894;
  assign tmp23891 = s9 ? tmp23892 : tmp23898;
  assign tmp23870 = s10 ? tmp23871 : tmp23891;
  assign tmp23869 = ~(s12 ? tmp23870 : tmp22562);
  assign tmp23828 = ~(s13 ? tmp23829 : tmp23869);
  assign tmp23796 = s14 ? tmp23797 : tmp23828;
  assign tmp23908 = s4 ? tmp22999 : tmp23739;
  assign tmp23911 = s3 ? tmp23211 : tmp22066;
  assign tmp23910 = s4 ? tmp23911 : tmp23744;
  assign tmp23909 = ~(s5 ? tmp23910 : tmp23011);
  assign tmp23907 = s6 ? tmp23908 : tmp23909;
  assign tmp23913 = s4 ? tmp22999 : tmp23752;
  assign tmp23915 = s4 ? tmp23911 : tmp23756;
  assign tmp23914 = ~(s5 ? tmp23915 : tmp23027);
  assign tmp23912 = s6 ? tmp23913 : tmp23914;
  assign tmp23906 = s7 ? tmp23907 : tmp23912;
  assign tmp23905 = s8 ? tmp23718 : tmp23906;
  assign tmp23904 = s9 ? tmp23696 : tmp23905;
  assign tmp23920 = ~(s5 ? tmp23733 : tmp23057);
  assign tmp23919 = s6 ? tmp23730 : tmp23920;
  assign tmp23918 = s7 ? tmp23719 : tmp23919;
  assign tmp23917 = s8 ? tmp23918 : tmp23719;
  assign tmp23922 = s7 ? tmp23785 : tmp23912;
  assign tmp23925 = ~(s5 ? tmp23733 : tmp23065);
  assign tmp23924 = s6 ? tmp23730 : tmp23925;
  assign tmp23923 = s7 ? tmp23924 : tmp23919;
  assign tmp23921 = s8 ? tmp23922 : tmp23923;
  assign tmp23916 = s9 ? tmp23917 : tmp23921;
  assign tmp23903 = s10 ? tmp23904 : tmp23916;
  assign tmp23929 = s7 ? tmp23709 : tmp23912;
  assign tmp23930 = s7 ? tmp23729 : tmp23919;
  assign tmp23928 = s8 ? tmp23929 : tmp23930;
  assign tmp23927 = s9 ? tmp23917 : tmp23928;
  assign tmp23926 = s10 ? tmp23904 : tmp23927;
  assign tmp23902 = ~(s11 ? tmp23903 : tmp23926);
  assign tmp23901 = s12 ? tmp22727 : tmp23902;
  assign tmp23900 = s13 ? tmp23901 : tmp23072;
  assign tmp23899 = s14 ? tmp22591 : tmp23900;
  assign tmp23795 = s15 ? tmp23796 : tmp23899;
  assign tmp23940 = s3 ? tmp21943 : tmp22611;
  assign tmp23939 = s4 ? tmp23500 : tmp23940;
  assign tmp23938 = s5 ? tmp23939 : tmp23503;
  assign tmp23937 = s6 ? tmp23495 : tmp23938;
  assign tmp23943 = s4 ? tmp23511 : tmp23876;
  assign tmp23945 = s3 ? tmp21943 : tmp22472;
  assign tmp23944 = s4 ? tmp23945 : tmp23504;
  assign tmp23942 = s5 ? tmp23943 : tmp23944;
  assign tmp23941 = s6 ? tmp23507 : tmp23942;
  assign tmp23936 = s7 ? tmp23937 : tmp23941;
  assign tmp23947 = s8 ? tmp23936 : tmp23937;
  assign tmp23946 = s9 ? tmp23947 : tmp23941;
  assign tmp23935 = s10 ? tmp23936 : tmp23946;
  assign tmp23934 = ~(s12 ? tmp23935 : tmp22562);
  assign tmp23933 = ~(s13 ? tmp23321 : tmp23934);
  assign tmp23932 = s14 ? tmp23240 : tmp23933;
  assign tmp23950 = s12 ? tmp22727 : tmp23693;
  assign tmp23949 = s13 ? tmp23950 : tmp23072;
  assign tmp23948 = s14 ? tmp22591 : tmp23949;
  assign tmp23931 = s15 ? tmp23932 : tmp23948;
  assign tmp23794 = s16 ? tmp23795 : tmp23931;
  assign tmp21926 = s17 ? tmp21927 : tmp23794;
  assign s12n = tmp21926;

  assign tmp23965 = ~(l4 ? 1 : 0);
  assign tmp23964 = l2 ? 1 : tmp23965;
  assign tmp23968 = l4 ? 1 : 0;
  assign tmp23967 = l3 ? tmp23968 : 0;
  assign tmp23966 = ~(l2 ? tmp23967 : 0);
  assign tmp23963 = l1 ? tmp23964 : tmp23966;
  assign tmp23974 = ~(l3 ? tmp23968 : 0);
  assign tmp23973 = l2 ? 1 : tmp23974;
  assign tmp23972 = l1 ? tmp23973 : tmp23966;
  assign tmp23971 = s0 ? tmp23963 : tmp23972;
  assign tmp23970 = s1 ? tmp23971 : tmp23963;
  assign tmp23969 = s2 ? tmp23963 : tmp23970;
  assign tmp23962 = s3 ? tmp23963 : tmp23969;
  assign tmp23978 = l1 ? tmp23973 : 1;
  assign tmp23977 = s0 ? tmp23963 : tmp23978;
  assign tmp23976 = s2 ? tmp23963 : tmp23977;
  assign tmp23984 = l3 ? 1 : tmp23965;
  assign tmp23983 = l2 ? 1 : tmp23984;
  assign tmp23982 = l1 ? tmp23983 : 1;
  assign tmp23981 = s0 ? tmp23978 : tmp23982;
  assign tmp23980 = s1 ? tmp23963 : tmp23981;
  assign tmp23987 = l1 ? tmp23983 : tmp23966;
  assign tmp23986 = s0 ? tmp23963 : tmp23987;
  assign tmp23988 = s0 ? tmp23982 : tmp23963;
  assign tmp23985 = s1 ? tmp23986 : tmp23988;
  assign tmp23979 = s2 ? tmp23980 : tmp23985;
  assign tmp23975 = s3 ? tmp23976 : tmp23979;
  assign tmp23961 = s4 ? tmp23962 : tmp23975;
  assign tmp23994 = s0 ? tmp23972 : tmp23963;
  assign tmp23993 = s1 ? tmp23971 : tmp23994;
  assign tmp23997 = l1 ? 1 : tmp23966;
  assign tmp23996 = s0 ? tmp23987 : tmp23997;
  assign tmp23995 = s1 ? tmp23994 : tmp23996;
  assign tmp23992 = s2 ? tmp23993 : tmp23995;
  assign tmp23999 = s0 ? tmp23997 : tmp23987;
  assign tmp24001 = s0 ? tmp23963 : tmp23982;
  assign tmp24000 = s1 ? tmp23982 : tmp24001;
  assign tmp23998 = s2 ? tmp23999 : tmp24000;
  assign tmp23991 = s3 ? tmp23992 : tmp23998;
  assign tmp24004 = s1 ? tmp23988 : tmp24001;
  assign tmp24005 = s1 ? tmp24001 : tmp23963;
  assign tmp24003 = s2 ? tmp24004 : tmp24005;
  assign tmp24007 = s1 ? tmp23987 : tmp23982;
  assign tmp24006 = s2 ? tmp24007 : tmp23982;
  assign tmp24002 = s3 ? tmp24003 : tmp24006;
  assign tmp23990 = s4 ? tmp23991 : tmp24002;
  assign tmp24012 = s0 ? tmp23987 : tmp23982;
  assign tmp24011 = s1 ? tmp24012 : tmp23982;
  assign tmp24014 = s0 ? tmp23982 : tmp23987;
  assign tmp24013 = s1 ? tmp24014 : tmp23987;
  assign tmp24010 = s2 ? tmp24011 : tmp24013;
  assign tmp24009 = s3 ? tmp24010 : tmp23982;
  assign tmp24016 = s2 ? tmp23982 : tmp24013;
  assign tmp24015 = s3 ? tmp24016 : tmp23982;
  assign tmp24008 = s4 ? tmp24009 : tmp24015;
  assign tmp23989 = s5 ? tmp23990 : tmp24008;
  assign tmp23960 = s6 ? tmp23961 : tmp23989;
  assign tmp24021 = s1 ? tmp23977 : tmp23963;
  assign tmp24020 = s2 ? tmp23963 : tmp24021;
  assign tmp24023 = s1 ? tmp23963 : tmp23982;
  assign tmp24022 = s2 ? tmp24023 : tmp23985;
  assign tmp24019 = s3 ? tmp24020 : tmp24022;
  assign tmp24018 = s4 ? tmp23962 : tmp24019;
  assign tmp24028 = s1 ? tmp23963 : tmp23996;
  assign tmp24027 = s2 ? tmp23970 : tmp24028;
  assign tmp24029 = s2 ? tmp23987 : tmp24000;
  assign tmp24026 = s3 ? tmp24027 : tmp24029;
  assign tmp24031 = s2 ? tmp24004 : tmp23963;
  assign tmp24030 = s3 ? tmp24031 : tmp24006;
  assign tmp24025 = s4 ? tmp24026 : tmp24030;
  assign tmp24034 = s2 ? tmp24011 : tmp24007;
  assign tmp24033 = s3 ? tmp24034 : tmp23982;
  assign tmp24036 = s2 ? tmp23982 : tmp23987;
  assign tmp24035 = s3 ? tmp24036 : tmp23982;
  assign tmp24032 = s4 ? tmp24033 : tmp24035;
  assign tmp24024 = s5 ? tmp24025 : tmp24032;
  assign tmp24017 = s6 ? tmp24018 : tmp24024;
  assign tmp23959 = s7 ? tmp23960 : tmp24017;
  assign tmp24044 = s0 ? tmp23987 : tmp23972;
  assign tmp24043 = s1 ? tmp23994 : tmp24044;
  assign tmp24042 = s2 ? tmp23993 : tmp24043;
  assign tmp24046 = s0 ? tmp23972 : tmp23987;
  assign tmp24045 = s2 ? tmp24046 : tmp24000;
  assign tmp24041 = s3 ? tmp24042 : tmp24045;
  assign tmp24048 = s2 ? tmp24011 : tmp23982;
  assign tmp24047 = s3 ? tmp24003 : tmp24048;
  assign tmp24040 = s4 ? tmp24041 : tmp24047;
  assign tmp24039 = s5 ? tmp24040 : tmp24008;
  assign tmp24038 = s6 ? tmp23961 : tmp24039;
  assign tmp24054 = s1 ? tmp23963 : tmp24044;
  assign tmp24053 = s2 ? tmp23970 : tmp24054;
  assign tmp24052 = s3 ? tmp24053 : tmp24029;
  assign tmp24055 = s3 ? tmp24031 : tmp24048;
  assign tmp24051 = s4 ? tmp24052 : tmp24055;
  assign tmp24050 = s5 ? tmp24051 : tmp24032;
  assign tmp24049 = s6 ? tmp24018 : tmp24050;
  assign tmp24037 = s7 ? tmp24038 : tmp24049;
  assign tmp23958 = s8 ? tmp23959 : tmp24037;
  assign tmp24059 = s4 ? tmp23963 : tmp23975;
  assign tmp24063 = s2 ? tmp23963 : tmp24028;
  assign tmp24062 = s3 ? tmp24063 : tmp23998;
  assign tmp24065 = s2 ? tmp23987 : tmp23982;
  assign tmp24064 = s3 ? tmp24003 : tmp24065;
  assign tmp24061 = s4 ? tmp24062 : tmp24064;
  assign tmp24060 = s5 ? tmp24061 : tmp24008;
  assign tmp24058 = s6 ? tmp24059 : tmp24060;
  assign tmp24067 = s4 ? tmp23963 : tmp24019;
  assign tmp24070 = s3 ? tmp24063 : tmp24029;
  assign tmp24069 = s4 ? tmp24070 : tmp24030;
  assign tmp24068 = s5 ? tmp24069 : tmp24032;
  assign tmp24066 = s6 ? tmp24067 : tmp24068;
  assign tmp24057 = s7 ? tmp24058 : tmp24066;
  assign tmp24056 = s8 ? tmp24037 : tmp24057;
  assign tmp23957 = s9 ? tmp23958 : tmp24056;
  assign tmp24072 = s8 ? tmp23959 : tmp23960;
  assign tmp24074 = s7 ? tmp24017 : tmp24066;
  assign tmp24075 = s7 ? tmp24049 : tmp24017;
  assign tmp24073 = s8 ? tmp24074 : tmp24075;
  assign tmp24071 = s9 ? tmp24072 : tmp24073;
  assign tmp23956 = s10 ? tmp23957 : tmp24071;
  assign tmp24084 = l1 ? tmp23973 : tmp23974;
  assign tmp24087 = s0 ? tmp24084 : tmp23973;
  assign tmp24086 = s2 ? tmp24084 : tmp24087;
  assign tmp24090 = s0 ? tmp23973 : tmp23997;
  assign tmp24089 = s1 ? tmp24084 : tmp24090;
  assign tmp24093 = l1 ? 1 : tmp23974;
  assign tmp24092 = s0 ? tmp24084 : tmp24093;
  assign tmp24094 = s0 ? tmp23997 : tmp24084;
  assign tmp24091 = s1 ? tmp24092 : tmp24094;
  assign tmp24088 = s2 ? tmp24089 : tmp24091;
  assign tmp24085 = s3 ? tmp24086 : tmp24088;
  assign tmp24083 = s4 ? tmp24084 : tmp24085;
  assign tmp24099 = s1 ? tmp24084 : tmp24093;
  assign tmp24098 = s2 ? tmp24084 : tmp24099;
  assign tmp24102 = s0 ? tmp23972 : tmp23997;
  assign tmp24101 = s1 ? tmp23997 : tmp24102;
  assign tmp24100 = s2 ? tmp24093 : tmp24101;
  assign tmp24097 = s3 ? tmp24098 : tmp24100;
  assign tmp24106 = s0 ? tmp23997 : tmp23972;
  assign tmp24105 = s1 ? tmp24106 : tmp24102;
  assign tmp24107 = s1 ? tmp24102 : tmp23972;
  assign tmp24104 = s2 ? tmp24105 : tmp24107;
  assign tmp24103 = s3 ? tmp24104 : tmp23997;
  assign tmp24096 = s4 ? tmp24097 : tmp24103;
  assign tmp24095 = s5 ? tmp24096 : tmp23997;
  assign tmp24082 = s6 ? tmp24083 : tmp24095;
  assign tmp24112 = s2 ? tmp24105 : tmp23972;
  assign tmp24111 = s3 ? tmp24112 : tmp23997;
  assign tmp24110 = s4 ? tmp24097 : tmp24111;
  assign tmp24109 = s5 ? tmp24110 : tmp23997;
  assign tmp24108 = s6 ? tmp24083 : tmp24109;
  assign tmp24081 = s7 ? tmp24082 : tmp24108;
  assign tmp24118 = s1 ? tmp24084 : tmp24094;
  assign tmp24117 = s2 ? tmp24089 : tmp24118;
  assign tmp24116 = s3 ? tmp24086 : tmp24117;
  assign tmp24115 = s4 ? tmp24084 : tmp24116;
  assign tmp24123 = s1 ? tmp24084 : tmp24092;
  assign tmp24125 = s0 ? tmp23972 : tmp23978;
  assign tmp24124 = s1 ? tmp23997 : tmp24125;
  assign tmp24122 = s2 ? tmp24123 : tmp24124;
  assign tmp24121 = s3 ? tmp24084 : tmp24122;
  assign tmp24128 = s1 ? tmp24106 : tmp24125;
  assign tmp24129 = s1 ? tmp24125 : tmp23972;
  assign tmp24127 = s2 ? tmp24128 : tmp24129;
  assign tmp24132 = s0 ? tmp23997 : tmp23978;
  assign tmp24133 = s0 ? tmp23978 : tmp23997;
  assign tmp24131 = s1 ? tmp24132 : tmp24133;
  assign tmp24130 = s2 ? tmp24131 : tmp23997;
  assign tmp24126 = s3 ? tmp24127 : tmp24130;
  assign tmp24120 = s4 ? tmp24121 : tmp24126;
  assign tmp24119 = s5 ? tmp24120 : tmp23997;
  assign tmp24114 = s6 ? tmp24115 : tmp24119;
  assign tmp24138 = s1 ? tmp24087 : tmp24084;
  assign tmp24137 = s2 ? tmp24084 : tmp24138;
  assign tmp24140 = s1 ? tmp24084 : tmp23997;
  assign tmp24139 = s2 ? tmp24140 : tmp24118;
  assign tmp24136 = s3 ? tmp24137 : tmp24139;
  assign tmp24135 = s4 ? tmp24084 : tmp24136;
  assign tmp24144 = s2 ? tmp24099 : tmp24124;
  assign tmp24143 = s3 ? tmp24084 : tmp24144;
  assign tmp24146 = s2 ? tmp24128 : tmp23972;
  assign tmp24148 = s1 ? tmp24132 : tmp23997;
  assign tmp24147 = s2 ? tmp24148 : tmp23997;
  assign tmp24145 = s3 ? tmp24146 : tmp24147;
  assign tmp24142 = s4 ? tmp24143 : tmp24145;
  assign tmp24141 = s5 ? tmp24142 : tmp23997;
  assign tmp24134 = s6 ? tmp24135 : tmp24141;
  assign tmp24113 = s7 ? tmp24114 : tmp24134;
  assign tmp24080 = s8 ? tmp24081 : tmp24113;
  assign tmp24157 = s0 ? tmp23972 : tmp23973;
  assign tmp24156 = s1 ? tmp24106 : tmp24157;
  assign tmp24158 = s1 ? tmp24157 : tmp23972;
  assign tmp24155 = s2 ? tmp24156 : tmp24158;
  assign tmp24154 = s3 ? tmp24155 : tmp23997;
  assign tmp24153 = s4 ? tmp24097 : tmp24154;
  assign tmp24152 = s5 ? tmp24153 : tmp23997;
  assign tmp24151 = s6 ? tmp24083 : tmp24152;
  assign tmp24162 = s2 ? tmp24140 : tmp24091;
  assign tmp24161 = s3 ? tmp24137 : tmp24162;
  assign tmp24160 = s4 ? tmp24084 : tmp24161;
  assign tmp24166 = s2 ? tmp24156 : tmp23972;
  assign tmp24165 = s3 ? tmp24166 : tmp23997;
  assign tmp24164 = s4 ? tmp24097 : tmp24165;
  assign tmp24163 = s5 ? tmp24164 : tmp23997;
  assign tmp24159 = s6 ? tmp24160 : tmp24163;
  assign tmp24150 = s7 ? tmp24151 : tmp24159;
  assign tmp24149 = s8 ? tmp24113 : tmp24150;
  assign tmp24079 = s9 ? tmp24080 : tmp24149;
  assign tmp24168 = s8 ? tmp24150 : tmp24151;
  assign tmp24173 = s3 ? tmp24086 : tmp24162;
  assign tmp24172 = s4 ? tmp24084 : tmp24173;
  assign tmp24178 = s1 ? tmp23972 : tmp24093;
  assign tmp24177 = s2 ? tmp24084 : tmp24178;
  assign tmp24180 = s1 ? tmp24093 : tmp23997;
  assign tmp24179 = s2 ? tmp24180 : tmp24101;
  assign tmp24176 = s3 ? tmp24177 : tmp24179;
  assign tmp24175 = s4 ? tmp24176 : tmp24111;
  assign tmp24174 = s5 ? tmp24175 : tmp23997;
  assign tmp24171 = s6 ? tmp24172 : tmp24174;
  assign tmp24184 = s3 ? tmp24177 : tmp24100;
  assign tmp24183 = s4 ? tmp24184 : tmp24165;
  assign tmp24182 = s5 ? tmp24183 : tmp23997;
  assign tmp24181 = s6 ? tmp24160 : tmp24182;
  assign tmp24170 = s7 ? tmp24171 : tmp24181;
  assign tmp24191 = s1 ? tmp23972 : tmp24084;
  assign tmp24190 = s2 ? tmp24084 : tmp24191;
  assign tmp24189 = s3 ? tmp24190 : tmp24144;
  assign tmp24188 = s4 ? tmp24189 : tmp24145;
  assign tmp24187 = s5 ? tmp24188 : tmp23997;
  assign tmp24186 = s6 ? tmp24135 : tmp24187;
  assign tmp24185 = s7 ? tmp24186 : tmp24181;
  assign tmp24169 = s8 ? tmp24170 : tmp24185;
  assign tmp24167 = s9 ? tmp24168 : tmp24169;
  assign tmp24078 = s10 ? tmp24079 : tmp24167;
  assign tmp24195 = s7 ? tmp24108 : tmp24159;
  assign tmp24196 = s7 ? tmp24134 : tmp24159;
  assign tmp24194 = s8 ? tmp24195 : tmp24196;
  assign tmp24193 = s9 ? tmp24168 : tmp24194;
  assign tmp24192 = s10 ? tmp24079 : tmp24193;
  assign tmp24077 = s11 ? tmp24078 : tmp24192;
  assign tmp24207 = s0 ? tmp23973 : 1;
  assign tmp24206 = s1 ? tmp23973 : tmp24207;
  assign tmp24210 = l1 ? 1 : tmp23973;
  assign tmp24209 = s0 ? tmp23973 : tmp24210;
  assign tmp24211 = s0 ? tmp24210 : tmp23973;
  assign tmp24208 = s1 ? tmp24209 : tmp24211;
  assign tmp24205 = s2 ? tmp24206 : tmp24208;
  assign tmp24204 = s3 ? tmp23973 : tmp24205;
  assign tmp24203 = s4 ? tmp23973 : tmp24204;
  assign tmp24216 = s1 ? tmp23973 : tmp24210;
  assign tmp24215 = s2 ? tmp23973 : tmp24216;
  assign tmp24218 = s1 ? tmp24210 : tmp24211;
  assign tmp24220 = s0 ? tmp23978 : tmp23973;
  assign tmp24219 = s1 ? tmp24210 : tmp24220;
  assign tmp24217 = s2 ? tmp24218 : tmp24219;
  assign tmp24214 = s3 ? tmp24215 : tmp24217;
  assign tmp24224 = s0 ? 1 : tmp23978;
  assign tmp24223 = s1 ? tmp24224 : tmp24220;
  assign tmp24225 = s1 ? tmp24220 : tmp23978;
  assign tmp24222 = s2 ? tmp24223 : tmp24225;
  assign tmp24228 = s0 ? tmp23973 : tmp23978;
  assign tmp24227 = s1 ? tmp23973 : tmp24228;
  assign tmp24230 = s0 ? 1 : tmp24210;
  assign tmp24229 = s1 ? tmp24210 : tmp24230;
  assign tmp24226 = s2 ? tmp24227 : tmp24229;
  assign tmp24221 = s3 ? tmp24222 : tmp24226;
  assign tmp24213 = s4 ? tmp24214 : tmp24221;
  assign tmp24234 = s1 ? tmp24209 : tmp24210;
  assign tmp24235 = s1 ? tmp24211 : tmp24220;
  assign tmp24233 = s2 ? tmp24234 : tmp24235;
  assign tmp24238 = s0 ? tmp23978 : tmp24210;
  assign tmp24237 = s1 ? tmp23978 : tmp24238;
  assign tmp24240 = s0 ? tmp24210 : 1;
  assign tmp24239 = s1 ? tmp24240 : tmp24224;
  assign tmp24236 = s2 ? tmp24237 : tmp24239;
  assign tmp24232 = s3 ? tmp24233 : tmp24236;
  assign tmp24244 = s0 ? tmp23978 : 1;
  assign tmp24243 = s1 ? tmp24244 : tmp24230;
  assign tmp24245 = s1 ? tmp24211 : tmp24228;
  assign tmp24242 = s2 ? tmp24243 : tmp24245;
  assign tmp24248 = s0 ? tmp24210 : tmp23978;
  assign tmp24247 = s1 ? tmp24240 : tmp24248;
  assign tmp24249 = s1 ? tmp24224 : tmp24244;
  assign tmp24246 = s2 ? tmp24247 : tmp24249;
  assign tmp24241 = s3 ? tmp24242 : tmp24246;
  assign tmp24231 = s4 ? tmp24232 : tmp24241;
  assign tmp24212 = s5 ? tmp24213 : tmp24231;
  assign tmp24202 = s6 ? tmp24203 : tmp24212;
  assign tmp24255 = s1 ? tmp23978 : tmp24210;
  assign tmp24254 = s2 ? tmp23973 : tmp24255;
  assign tmp24257 = s1 ? tmp24210 : tmp23973;
  assign tmp24256 = s2 ? tmp24257 : tmp24219;
  assign tmp24253 = s3 ? tmp24254 : tmp24256;
  assign tmp24259 = s2 ? tmp24223 : tmp23978;
  assign tmp24261 = s1 ? tmp23973 : tmp23978;
  assign tmp24262 = s1 ? tmp24210 : 1;
  assign tmp24260 = s2 ? tmp24261 : tmp24262;
  assign tmp24258 = s3 ? tmp24259 : tmp24260;
  assign tmp24252 = s4 ? tmp24253 : tmp24258;
  assign tmp24265 = s2 ? tmp24234 : tmp24261;
  assign tmp24267 = s1 ? 1 : tmp23978;
  assign tmp24266 = s2 ? tmp24255 : tmp24267;
  assign tmp24264 = s3 ? tmp24265 : tmp24266;
  assign tmp24270 = s1 ? 1 : tmp24210;
  assign tmp24269 = s2 ? tmp24270 : tmp23973;
  assign tmp24268 = s3 ? tmp24269 : tmp24267;
  assign tmp24263 = s4 ? tmp24264 : tmp24268;
  assign tmp24251 = s5 ? tmp24252 : tmp24263;
  assign tmp24250 = s6 ? tmp24203 : tmp24251;
  assign tmp24201 = s7 ? tmp24202 : tmp24250;
  assign tmp24276 = s1 ? tmp23973 : tmp24211;
  assign tmp24275 = s2 ? tmp24206 : tmp24276;
  assign tmp24274 = s3 ? tmp23973 : tmp24275;
  assign tmp24273 = s4 ? tmp23973 : tmp24274;
  assign tmp24281 = s1 ? tmp24228 : tmp23973;
  assign tmp24280 = s2 ? tmp23973 : tmp24281;
  assign tmp24283 = s1 ? tmp24210 : tmp23978;
  assign tmp24282 = s2 ? tmp24227 : tmp24283;
  assign tmp24279 = s3 ? tmp24280 : tmp24282;
  assign tmp24286 = s1 ? tmp24224 : tmp23978;
  assign tmp24285 = s2 ? tmp24286 : tmp23978;
  assign tmp24287 = s2 ? tmp23978 : tmp24229;
  assign tmp24284 = s3 ? tmp24285 : tmp24287;
  assign tmp24278 = s4 ? tmp24279 : tmp24284;
  assign tmp24291 = s1 ? tmp24238 : tmp24210;
  assign tmp24292 = s1 ? tmp24248 : tmp23978;
  assign tmp24290 = s2 ? tmp24291 : tmp24292;
  assign tmp24289 = s3 ? tmp24290 : tmp24236;
  assign tmp24294 = s2 ? tmp24243 : tmp24292;
  assign tmp24293 = s3 ? tmp24294 : tmp24246;
  assign tmp24288 = s4 ? tmp24289 : tmp24293;
  assign tmp24277 = s5 ? tmp24278 : tmp24288;
  assign tmp24272 = s6 ? tmp24273 : tmp24277;
  assign tmp24298 = s2 ? tmp23973 : tmp24261;
  assign tmp24300 = s1 ? tmp23973 : 1;
  assign tmp24299 = s2 ? tmp24300 : tmp24276;
  assign tmp24297 = s3 ? tmp24298 : tmp24299;
  assign tmp24296 = s4 ? tmp23973 : tmp24297;
  assign tmp24305 = s1 ? tmp23978 : tmp23973;
  assign tmp24304 = s2 ? tmp23973 : tmp24305;
  assign tmp24306 = s2 ? tmp24261 : tmp24283;
  assign tmp24303 = s3 ? tmp24304 : tmp24306;
  assign tmp24308 = s2 ? tmp23978 : tmp24262;
  assign tmp24307 = s3 ? tmp24285 : tmp24308;
  assign tmp24302 = s4 ? tmp24303 : tmp24307;
  assign tmp24311 = s2 ? tmp24291 : tmp23978;
  assign tmp24310 = s3 ? tmp24311 : tmp24266;
  assign tmp24313 = s2 ? tmp24270 : tmp23978;
  assign tmp24312 = s3 ? tmp24313 : tmp24267;
  assign tmp24309 = s4 ? tmp24310 : tmp24312;
  assign tmp24301 = s5 ? tmp24302 : tmp24309;
  assign tmp24295 = s6 ? tmp24296 : tmp24301;
  assign tmp24271 = s7 ? tmp24272 : tmp24295;
  assign tmp24200 = s8 ? tmp24201 : tmp24271;
  assign tmp24321 = s1 ? tmp24210 : tmp24248;
  assign tmp24320 = s2 ? tmp24321 : tmp24283;
  assign tmp24319 = s3 ? tmp24215 : tmp24320;
  assign tmp24318 = s4 ? tmp24319 : tmp24284;
  assign tmp24317 = s5 ? tmp24318 : tmp24288;
  assign tmp24316 = s6 ? tmp24203 : tmp24317;
  assign tmp24325 = s2 ? tmp24300 : tmp24208;
  assign tmp24324 = s3 ? tmp24298 : tmp24325;
  assign tmp24323 = s4 ? tmp23973 : tmp24324;
  assign tmp24328 = s3 ? tmp24254 : tmp24283;
  assign tmp24327 = s4 ? tmp24328 : tmp24307;
  assign tmp24326 = s5 ? tmp24327 : tmp24309;
  assign tmp24322 = s6 ? tmp24323 : tmp24326;
  assign tmp24315 = s7 ? tmp24316 : tmp24322;
  assign tmp24314 = s8 ? tmp24271 : tmp24315;
  assign tmp24199 = s9 ? tmp24200 : tmp24314;
  assign tmp24330 = s8 ? tmp24315 : tmp24316;
  assign tmp24335 = s3 ? tmp23973 : tmp24325;
  assign tmp24334 = s4 ? tmp23973 : tmp24335;
  assign tmp24333 = s6 ? tmp24334 : tmp24251;
  assign tmp24332 = s7 ? tmp24333 : tmp24322;
  assign tmp24336 = s7 ? tmp24295 : tmp24322;
  assign tmp24331 = s8 ? tmp24332 : tmp24336;
  assign tmp24329 = s9 ? tmp24330 : tmp24331;
  assign tmp24198 = s10 ? tmp24199 : tmp24329;
  assign tmp24340 = s7 ? tmp24250 : tmp24322;
  assign tmp24339 = s8 ? tmp24340 : tmp24336;
  assign tmp24338 = s9 ? tmp24330 : tmp24339;
  assign tmp24337 = s10 ? tmp24199 : tmp24338;
  assign tmp24197 = s11 ? tmp24198 : tmp24337;
  assign tmp24076 = s12 ? tmp24077 : tmp24197;
  assign tmp23955 = s13 ? tmp23956 : tmp24076;
  assign tmp24352 = s0 ? tmp24093 : tmp24210;
  assign tmp24351 = s2 ? tmp24093 : tmp24352;
  assign tmp24355 = s0 ? tmp24210 : tmp23997;
  assign tmp24354 = s1 ? tmp24093 : tmp24355;
  assign tmp24357 = s0 ? tmp23997 : tmp24093;
  assign tmp24356 = s1 ? tmp24093 : tmp24357;
  assign tmp24353 = s2 ? tmp24354 : tmp24356;
  assign tmp24350 = s3 ? tmp24351 : tmp24353;
  assign tmp24349 = s4 ? tmp24093 : tmp24350;
  assign tmp24361 = s2 ? tmp24093 : tmp23997;
  assign tmp24360 = s3 ? tmp24093 : tmp24361;
  assign tmp24359 = s4 ? tmp24360 : tmp23997;
  assign tmp24358 = s5 ? tmp24359 : tmp23997;
  assign tmp24348 = s6 ? tmp24349 : tmp24358;
  assign tmp24366 = s1 ? tmp24352 : tmp24093;
  assign tmp24365 = s2 ? tmp24093 : tmp24366;
  assign tmp24367 = s2 ? tmp24180 : tmp24356;
  assign tmp24364 = s3 ? tmp24365 : tmp24367;
  assign tmp24363 = s4 ? tmp24093 : tmp24364;
  assign tmp24372 = s1 ? tmp23997 : tmp24093;
  assign tmp24371 = s2 ? tmp24093 : tmp24372;
  assign tmp24370 = s3 ? tmp24371 : tmp24361;
  assign tmp24369 = s4 ? tmp24370 : tmp23997;
  assign tmp24368 = s5 ? tmp24369 : tmp23997;
  assign tmp24362 = s6 ? tmp24363 : tmp24368;
  assign tmp24347 = s7 ? tmp24348 : tmp24362;
  assign tmp24380 = s0 ? tmp24093 : tmp23997;
  assign tmp24379 = s1 ? tmp24380 : tmp24093;
  assign tmp24378 = s2 ? tmp24093 : tmp24379;
  assign tmp24377 = s3 ? tmp24378 : tmp24361;
  assign tmp24376 = s4 ? tmp24377 : tmp23997;
  assign tmp24375 = s5 ? tmp24376 : tmp23997;
  assign tmp24374 = s6 ? tmp24349 : tmp24375;
  assign tmp24373 = s7 ? tmp24374 : tmp24362;
  assign tmp24346 = s8 ? tmp24347 : tmp24373;
  assign tmp24345 = s9 ? tmp24346 : tmp24373;
  assign tmp24382 = s8 ? tmp24373 : tmp24374;
  assign tmp24389 = s2 ? tmp24180 : tmp23997;
  assign tmp24388 = s3 ? tmp24371 : tmp24389;
  assign tmp24387 = s4 ? tmp24388 : tmp23997;
  assign tmp24386 = s5 ? tmp24387 : tmp23997;
  assign tmp24385 = s6 ? tmp24363 : tmp24386;
  assign tmp24384 = s7 ? tmp24385 : tmp24362;
  assign tmp24383 = s8 ? tmp24384 : tmp24362;
  assign tmp24381 = s9 ? tmp24382 : tmp24383;
  assign tmp24344 = s10 ? tmp24345 : tmp24381;
  assign tmp24391 = s9 ? tmp24382 : tmp24362;
  assign tmp24390 = s10 ? tmp24345 : tmp24391;
  assign tmp24343 = s11 ? tmp24344 : tmp24390;
  assign tmp24401 = l3 ? 1 : tmp23968;
  assign tmp24400 = l2 ? tmp24401 : 1;
  assign tmp24399 = l1 ? tmp23983 : tmp24400;
  assign tmp24404 = s0 ? tmp24399 : tmp23982;
  assign tmp24403 = s1 ? tmp24404 : tmp24399;
  assign tmp24402 = s2 ? tmp24399 : tmp24403;
  assign tmp24398 = s3 ? tmp24399 : tmp24402;
  assign tmp24406 = s2 ? tmp24403 : tmp24404;
  assign tmp24410 = l1 ? 1 : tmp24400;
  assign tmp24409 = s0 ? tmp23982 : tmp24410;
  assign tmp24408 = s1 ? tmp24399 : tmp24409;
  assign tmp24412 = s0 ? tmp24410 : tmp24399;
  assign tmp24411 = s1 ? tmp24399 : tmp24412;
  assign tmp24407 = s2 ? tmp24408 : tmp24411;
  assign tmp24405 = s3 ? tmp24406 : tmp24407;
  assign tmp24397 = s4 ? tmp24398 : tmp24405;
  assign tmp24417 = s1 ? tmp24404 : tmp23982;
  assign tmp24419 = s0 ? tmp23982 : tmp24399;
  assign tmp24418 = s1 ? tmp24419 : tmp24399;
  assign tmp24416 = s2 ? tmp24417 : tmp24418;
  assign tmp24421 = s1 ? tmp24410 : tmp24399;
  assign tmp24420 = s2 ? tmp24399 : tmp24421;
  assign tmp24415 = s3 ? tmp24416 : tmp24420;
  assign tmp24424 = s1 ? tmp24412 : tmp24399;
  assign tmp24425 = s1 ? tmp24399 : tmp24404;
  assign tmp24423 = s2 ? tmp24424 : tmp24425;
  assign tmp24426 = s2 ? tmp24399 : tmp24410;
  assign tmp24422 = s3 ? tmp24423 : tmp24426;
  assign tmp24414 = s4 ? tmp24415 : tmp24422;
  assign tmp24431 = s0 ? tmp24399 : tmp24410;
  assign tmp24430 = s1 ? tmp24431 : tmp24410;
  assign tmp24433 = s0 ? tmp24410 : tmp23982;
  assign tmp24432 = s1 ? tmp24433 : tmp23982;
  assign tmp24429 = s2 ? tmp24430 : tmp24432;
  assign tmp24435 = s1 ? tmp24409 : tmp24410;
  assign tmp24436 = s1 ? tmp24410 : tmp24412;
  assign tmp24434 = s2 ? tmp24435 : tmp24436;
  assign tmp24428 = s3 ? tmp24429 : tmp24434;
  assign tmp24439 = s1 ? tmp24412 : tmp23982;
  assign tmp24438 = s2 ? tmp24430 : tmp24439;
  assign tmp24441 = s1 ? tmp24412 : tmp24410;
  assign tmp24440 = s2 ? tmp24436 : tmp24441;
  assign tmp24437 = s3 ? tmp24438 : tmp24440;
  assign tmp24427 = s4 ? tmp24428 : tmp24437;
  assign tmp24413 = s5 ? tmp24414 : tmp24427;
  assign tmp24396 = s6 ? tmp24397 : tmp24413;
  assign tmp24446 = s1 ? tmp24399 : tmp24410;
  assign tmp24445 = s2 ? tmp24446 : tmp24411;
  assign tmp24444 = s3 ? tmp24403 : tmp24445;
  assign tmp24443 = s4 ? tmp24398 : tmp24444;
  assign tmp24450 = s2 ? tmp24417 : tmp24399;
  assign tmp24449 = s3 ? tmp24450 : tmp24420;
  assign tmp24452 = s2 ? tmp24424 : tmp24399;
  assign tmp24451 = s3 ? tmp24452 : tmp24426;
  assign tmp24448 = s4 ? tmp24449 : tmp24451;
  assign tmp24455 = s2 ? tmp24430 : tmp23982;
  assign tmp24456 = s2 ? tmp24410 : tmp24421;
  assign tmp24454 = s3 ? tmp24455 : tmp24456;
  assign tmp24458 = s2 ? tmp24410 : tmp24399;
  assign tmp24457 = s3 ? tmp24458 : tmp24421;
  assign tmp24453 = s4 ? tmp24454 : tmp24457;
  assign tmp24447 = s5 ? tmp24448 : tmp24453;
  assign tmp24442 = s6 ? tmp24443 : tmp24447;
  assign tmp24395 = s7 ? tmp24396 : tmp24442;
  assign tmp24465 = s1 ? tmp24419 : tmp24404;
  assign tmp24464 = s2 ? tmp24417 : tmp24465;
  assign tmp24466 = s2 ? tmp24419 : tmp24421;
  assign tmp24463 = s3 ? tmp24464 : tmp24466;
  assign tmp24462 = s4 ? tmp24463 : tmp24422;
  assign tmp24461 = s5 ? tmp24462 : tmp24427;
  assign tmp24460 = s6 ? tmp24397 : tmp24461;
  assign tmp24471 = s2 ? tmp24417 : tmp24425;
  assign tmp24470 = s3 ? tmp24471 : tmp24420;
  assign tmp24469 = s4 ? tmp24470 : tmp24451;
  assign tmp24468 = s5 ? tmp24469 : tmp24453;
  assign tmp24467 = s6 ? tmp24443 : tmp24468;
  assign tmp24459 = s7 ? tmp24460 : tmp24467;
  assign tmp24394 = s8 ? tmp24395 : tmp24459;
  assign tmp24477 = s2 ? tmp24399 : tmp24404;
  assign tmp24476 = s3 ? tmp24477 : tmp24407;
  assign tmp24475 = s4 ? tmp24398 : tmp24476;
  assign tmp24479 = s4 ? tmp24415 : tmp24451;
  assign tmp24478 = s5 ? tmp24479 : tmp24427;
  assign tmp24474 = s6 ? tmp24475 : tmp24478;
  assign tmp24482 = s3 ? tmp24402 : tmp24445;
  assign tmp24481 = s4 ? tmp24398 : tmp24482;
  assign tmp24480 = s6 ? tmp24481 : tmp24447;
  assign tmp24473 = s7 ? tmp24474 : tmp24480;
  assign tmp24472 = s8 ? tmp24459 : tmp24473;
  assign tmp24393 = s9 ? tmp24394 : tmp24472;
  assign tmp24484 = s8 ? tmp24395 : tmp24396;
  assign tmp24486 = s7 ? tmp24442 : tmp24480;
  assign tmp24487 = s7 ? tmp24467 : tmp24442;
  assign tmp24485 = s8 ? tmp24486 : tmp24487;
  assign tmp24483 = s9 ? tmp24484 : tmp24485;
  assign tmp24392 = s10 ? tmp24393 : tmp24483;
  assign tmp24342 = s12 ? tmp24343 : tmp24392;
  assign tmp24499 = l2 ? tmp24401 : tmp23984;
  assign tmp24501 = ~(l3 ? 1 : tmp23965);
  assign tmp24500 = ~(l2 ? tmp23967 : tmp24501);
  assign tmp24498 = l1 ? tmp24499 : tmp24500;
  assign tmp24502 = s0 ? tmp23987 : tmp24498;
  assign tmp24497 = s1 ? tmp24498 : tmp24502;
  assign tmp24505 = s0 ? tmp24498 : tmp23997;
  assign tmp24504 = s1 ? tmp24505 : tmp24498;
  assign tmp24503 = s2 ? tmp24498 : tmp24504;
  assign tmp24496 = s3 ? tmp24497 : tmp24503;
  assign tmp24509 = s0 ? tmp24498 : tmp23987;
  assign tmp24508 = s1 ? tmp24509 : tmp24498;
  assign tmp24510 = s1 ? tmp24505 : tmp23996;
  assign tmp24507 = s2 ? tmp24508 : tmp24510;
  assign tmp24514 = l1 ? tmp24400 : 1;
  assign tmp24513 = s0 ? tmp23997 : tmp24514;
  assign tmp24512 = s1 ? tmp23987 : tmp24513;
  assign tmp24516 = s0 ? tmp24514 : tmp24498;
  assign tmp24515 = s1 ? tmp24498 : tmp24516;
  assign tmp24511 = s2 ? tmp24512 : tmp24515;
  assign tmp24506 = s3 ? tmp24507 : tmp24511;
  assign tmp24495 = s4 ? tmp24496 : tmp24506;
  assign tmp24522 = s0 ? tmp23997 : tmp24498;
  assign tmp24521 = s1 ? tmp24505 : tmp24522;
  assign tmp24523 = s1 ? tmp24522 : tmp24505;
  assign tmp24520 = s2 ? tmp24521 : tmp24523;
  assign tmp24527 = l1 ? tmp24499 : tmp23983;
  assign tmp24526 = s0 ? tmp24498 : tmp24527;
  assign tmp24525 = s1 ? tmp24514 : tmp24526;
  assign tmp24524 = s2 ? tmp24522 : tmp24525;
  assign tmp24519 = s3 ? tmp24520 : tmp24524;
  assign tmp24531 = s0 ? tmp23987 : tmp23983;
  assign tmp24530 = s1 ? tmp24516 : tmp24531;
  assign tmp24532 = s1 ? tmp24531 : tmp24509;
  assign tmp24529 = s2 ? tmp24530 : tmp24532;
  assign tmp24536 = l1 ? tmp24499 : 1;
  assign tmp24535 = s0 ? tmp23982 : tmp24536;
  assign tmp24534 = s1 ? tmp24526 : tmp24535;
  assign tmp24533 = s2 ? tmp24534 : tmp24514;
  assign tmp24528 = s3 ? tmp24529 : tmp24533;
  assign tmp24518 = s4 ? tmp24519 : tmp24528;
  assign tmp24541 = s0 ? tmp24498 : tmp24514;
  assign tmp24540 = s1 ? tmp24541 : tmp24514;
  assign tmp24543 = s0 ? tmp24536 : tmp24498;
  assign tmp24544 = s0 ? tmp24527 : tmp24498;
  assign tmp24542 = s1 ? tmp24543 : tmp24544;
  assign tmp24539 = s2 ? tmp24540 : tmp24542;
  assign tmp24547 = s0 ? tmp24536 : tmp24514;
  assign tmp24546 = s1 ? tmp24547 : tmp24514;
  assign tmp24549 = s0 ? tmp24514 : tmp24536;
  assign tmp24548 = s1 ? tmp24514 : tmp24549;
  assign tmp24545 = s2 ? tmp24546 : tmp24548;
  assign tmp24538 = s3 ? tmp24539 : tmp24545;
  assign tmp24552 = s1 ? tmp24516 : tmp24526;
  assign tmp24551 = s2 ? tmp24536 : tmp24552;
  assign tmp24554 = s1 ? tmp24549 : tmp24514;
  assign tmp24553 = s2 ? tmp24548 : tmp24554;
  assign tmp24550 = s3 ? tmp24551 : tmp24553;
  assign tmp24537 = s4 ? tmp24538 : tmp24550;
  assign tmp24517 = s5 ? tmp24518 : tmp24537;
  assign tmp24494 = s6 ? tmp24495 : tmp24517;
  assign tmp24559 = s1 ? tmp24505 : tmp23987;
  assign tmp24558 = s2 ? tmp24508 : tmp24559;
  assign tmp24561 = s1 ? tmp23987 : tmp24514;
  assign tmp24560 = s2 ? tmp24561 : tmp24515;
  assign tmp24557 = s3 ? tmp24558 : tmp24560;
  assign tmp24556 = s4 ? tmp24496 : tmp24557;
  assign tmp24566 = s1 ? tmp24498 : tmp24505;
  assign tmp24565 = s2 ? tmp24504 : tmp24566;
  assign tmp24567 = s2 ? tmp24498 : tmp24525;
  assign tmp24564 = s3 ? tmp24565 : tmp24567;
  assign tmp24569 = s2 ? tmp24530 : tmp24498;
  assign tmp24571 = s1 ? tmp24526 : tmp24536;
  assign tmp24570 = s2 ? tmp24571 : tmp24514;
  assign tmp24568 = s3 ? tmp24569 : tmp24570;
  assign tmp24563 = s4 ? tmp24564 : tmp24568;
  assign tmp24575 = s1 ? tmp24498 : tmp24544;
  assign tmp24574 = s2 ? tmp24540 : tmp24575;
  assign tmp24578 = s0 ? tmp24527 : tmp24514;
  assign tmp24577 = s1 ? tmp24578 : tmp24514;
  assign tmp24579 = s1 ? tmp24514 : tmp24536;
  assign tmp24576 = s2 ? tmp24577 : tmp24579;
  assign tmp24573 = s3 ? tmp24574 : tmp24576;
  assign tmp24582 = s1 ? tmp24498 : tmp24526;
  assign tmp24581 = s2 ? tmp24514 : tmp24582;
  assign tmp24580 = s3 ? tmp24581 : tmp24536;
  assign tmp24572 = s4 ? tmp24573 : tmp24580;
  assign tmp24562 = s5 ? tmp24563 : tmp24572;
  assign tmp24555 = s6 ? tmp24556 : tmp24562;
  assign tmp24493 = s7 ? tmp24494 : tmp24555;
  assign tmp24588 = l1 ? tmp24499 : tmp23966;
  assign tmp24589 = s0 ? tmp23987 : tmp24588;
  assign tmp24587 = s1 ? tmp24588 : tmp24589;
  assign tmp24593 = l1 ? tmp24400 : tmp23966;
  assign tmp24592 = s0 ? tmp24588 : tmp24593;
  assign tmp24591 = s1 ? tmp24592 : tmp24588;
  assign tmp24590 = s2 ? tmp24588 : tmp24591;
  assign tmp24586 = s3 ? tmp24587 : tmp24590;
  assign tmp24597 = s0 ? tmp24588 : tmp23987;
  assign tmp24596 = s1 ? tmp24597 : tmp24588;
  assign tmp24599 = s0 ? tmp24588 : tmp23997;
  assign tmp24598 = s1 ? tmp24599 : tmp23996;
  assign tmp24595 = s2 ? tmp24596 : tmp24598;
  assign tmp24602 = s0 ? tmp24514 : tmp24588;
  assign tmp24601 = s1 ? tmp24588 : tmp24602;
  assign tmp24600 = s2 ? tmp24512 : tmp24601;
  assign tmp24594 = s3 ? tmp24595 : tmp24600;
  assign tmp24585 = s4 ? tmp24586 : tmp24594;
  assign tmp24608 = s0 ? tmp23997 : tmp24588;
  assign tmp24607 = s1 ? tmp24599 : tmp24608;
  assign tmp24609 = s1 ? tmp24608 : tmp24592;
  assign tmp24606 = s2 ? tmp24607 : tmp24609;
  assign tmp24611 = s0 ? tmp24593 : tmp24588;
  assign tmp24612 = s1 ? tmp24514 : tmp24588;
  assign tmp24610 = s2 ? tmp24611 : tmp24612;
  assign tmp24605 = s3 ? tmp24606 : tmp24610;
  assign tmp24615 = s1 ? tmp24602 : tmp24012;
  assign tmp24616 = s1 ? tmp24012 : tmp24597;
  assign tmp24614 = s2 ? tmp24615 : tmp24616;
  assign tmp24618 = s1 ? tmp24588 : tmp24535;
  assign tmp24617 = s2 ? tmp24618 : tmp24514;
  assign tmp24613 = s3 ? tmp24614 : tmp24617;
  assign tmp24604 = s4 ? tmp24605 : tmp24613;
  assign tmp24623 = s0 ? tmp24588 : tmp24514;
  assign tmp24622 = s1 ? tmp24623 : tmp24514;
  assign tmp24625 = s0 ? tmp24536 : tmp24588;
  assign tmp24624 = s1 ? tmp24602 : tmp24625;
  assign tmp24621 = s2 ? tmp24622 : tmp24624;
  assign tmp24620 = s3 ? tmp24621 : tmp24545;
  assign tmp24628 = s1 ? tmp24536 : tmp24514;
  assign tmp24630 = s0 ? tmp24588 : tmp24536;
  assign tmp24629 = s1 ? tmp24602 : tmp24630;
  assign tmp24627 = s2 ? tmp24628 : tmp24629;
  assign tmp24626 = s3 ? tmp24627 : tmp24553;
  assign tmp24619 = s4 ? tmp24620 : tmp24626;
  assign tmp24603 = s5 ? tmp24604 : tmp24619;
  assign tmp24584 = s6 ? tmp24585 : tmp24603;
  assign tmp24635 = s1 ? tmp24599 : tmp23987;
  assign tmp24634 = s2 ? tmp24596 : tmp24635;
  assign tmp24636 = s2 ? tmp24561 : tmp24601;
  assign tmp24633 = s3 ? tmp24634 : tmp24636;
  assign tmp24632 = s4 ? tmp24586 : tmp24633;
  assign tmp24641 = s1 ? tmp24599 : tmp24588;
  assign tmp24642 = s1 ? tmp24588 : tmp24592;
  assign tmp24640 = s2 ? tmp24641 : tmp24642;
  assign tmp24643 = s2 ? tmp24588 : tmp24612;
  assign tmp24639 = s3 ? tmp24640 : tmp24643;
  assign tmp24645 = s2 ? tmp24615 : tmp24588;
  assign tmp24647 = s1 ? tmp24588 : tmp24536;
  assign tmp24646 = s2 ? tmp24647 : tmp24514;
  assign tmp24644 = s3 ? tmp24645 : tmp24646;
  assign tmp24638 = s4 ? tmp24639 : tmp24644;
  assign tmp24650 = s2 ? tmp24622 : tmp24647;
  assign tmp24649 = s3 ? tmp24650 : tmp24576;
  assign tmp24653 = s1 ? tmp24588 : tmp24527;
  assign tmp24652 = s2 ? tmp24514 : tmp24653;
  assign tmp24651 = s3 ? tmp24652 : tmp24536;
  assign tmp24648 = s4 ? tmp24649 : tmp24651;
  assign tmp24637 = s5 ? tmp24638 : tmp24648;
  assign tmp24631 = s6 ? tmp24632 : tmp24637;
  assign tmp24583 = s7 ? tmp24584 : tmp24631;
  assign tmp24492 = s8 ? tmp24493 : tmp24583;
  assign tmp24659 = s2 ? tmp24588 : tmp24641;
  assign tmp24658 = s3 ? tmp24587 : tmp24659;
  assign tmp24657 = s4 ? tmp24658 : tmp24594;
  assign tmp24664 = s1 ? tmp24608 : tmp24599;
  assign tmp24663 = s2 ? tmp24607 : tmp24664;
  assign tmp24667 = s0 ? tmp24588 : tmp24498;
  assign tmp24666 = s1 ? tmp24514 : tmp24667;
  assign tmp24665 = s2 ? tmp24608 : tmp24666;
  assign tmp24662 = s3 ? tmp24663 : tmp24665;
  assign tmp24670 = s1 ? tmp24602 : tmp24531;
  assign tmp24671 = s1 ? tmp24531 : tmp24597;
  assign tmp24669 = s2 ? tmp24670 : tmp24671;
  assign tmp24673 = s1 ? tmp24667 : tmp24535;
  assign tmp24672 = s2 ? tmp24673 : tmp24514;
  assign tmp24668 = s3 ? tmp24669 : tmp24672;
  assign tmp24661 = s4 ? tmp24662 : tmp24668;
  assign tmp24678 = s0 ? tmp24498 : tmp24588;
  assign tmp24677 = s1 ? tmp24625 : tmp24678;
  assign tmp24676 = s2 ? tmp24622 : tmp24677;
  assign tmp24675 = s3 ? tmp24676 : tmp24545;
  assign tmp24681 = s1 ? tmp24602 : tmp24667;
  assign tmp24680 = s2 ? tmp24536 : tmp24681;
  assign tmp24679 = s3 ? tmp24680 : tmp24553;
  assign tmp24674 = s4 ? tmp24675 : tmp24679;
  assign tmp24660 = s5 ? tmp24661 : tmp24674;
  assign tmp24656 = s6 ? tmp24657 : tmp24660;
  assign tmp24683 = s4 ? tmp24658 : tmp24633;
  assign tmp24688 = s1 ? tmp24588 : tmp24599;
  assign tmp24687 = s2 ? tmp24641 : tmp24688;
  assign tmp24689 = s2 ? tmp24588 : tmp24666;
  assign tmp24686 = s3 ? tmp24687 : tmp24689;
  assign tmp24691 = s2 ? tmp24670 : tmp24588;
  assign tmp24693 = s1 ? tmp24667 : tmp24536;
  assign tmp24692 = s2 ? tmp24693 : tmp24514;
  assign tmp24690 = s3 ? tmp24691 : tmp24692;
  assign tmp24685 = s4 ? tmp24686 : tmp24690;
  assign tmp24696 = s2 ? tmp24546 : tmp24579;
  assign tmp24695 = s3 ? tmp24650 : tmp24696;
  assign tmp24699 = s1 ? tmp24588 : tmp24498;
  assign tmp24698 = s2 ? tmp24514 : tmp24699;
  assign tmp24697 = s3 ? tmp24698 : tmp24536;
  assign tmp24694 = s4 ? tmp24695 : tmp24697;
  assign tmp24684 = s5 ? tmp24685 : tmp24694;
  assign tmp24682 = s6 ? tmp24683 : tmp24684;
  assign tmp24655 = s7 ? tmp24656 : tmp24682;
  assign tmp24654 = s8 ? tmp24583 : tmp24655;
  assign tmp24491 = s9 ? tmp24492 : tmp24654;
  assign tmp24708 = s1 ? tmp24498 : tmp24536;
  assign tmp24707 = s2 ? tmp24540 : tmp24708;
  assign tmp24706 = s3 ? tmp24707 : tmp24576;
  assign tmp24711 = s1 ? tmp24498 : tmp24527;
  assign tmp24710 = s2 ? tmp24514 : tmp24711;
  assign tmp24709 = s3 ? tmp24710 : tmp24536;
  assign tmp24705 = s4 ? tmp24706 : tmp24709;
  assign tmp24704 = s5 ? tmp24563 : tmp24705;
  assign tmp24703 = s6 ? tmp24556 : tmp24704;
  assign tmp24702 = s7 ? tmp24494 : tmp24703;
  assign tmp24701 = s8 ? tmp24702 : tmp24494;
  assign tmp24718 = s2 ? tmp24514 : tmp24498;
  assign tmp24717 = s3 ? tmp24718 : tmp24536;
  assign tmp24716 = s4 ? tmp24573 : tmp24717;
  assign tmp24715 = s5 ? tmp24563 : tmp24716;
  assign tmp24714 = s6 ? tmp24556 : tmp24715;
  assign tmp24723 = s2 ? tmp24514 : tmp24588;
  assign tmp24722 = s3 ? tmp24723 : tmp24536;
  assign tmp24721 = s4 ? tmp24695 : tmp24722;
  assign tmp24720 = s5 ? tmp24685 : tmp24721;
  assign tmp24719 = s6 ? tmp24683 : tmp24720;
  assign tmp24713 = s7 ? tmp24714 : tmp24719;
  assign tmp24727 = s4 ? tmp24649 : tmp24722;
  assign tmp24726 = s5 ? tmp24638 : tmp24727;
  assign tmp24725 = s6 ? tmp24632 : tmp24726;
  assign tmp24730 = s4 ? tmp24706 : tmp24717;
  assign tmp24729 = s5 ? tmp24563 : tmp24730;
  assign tmp24728 = s6 ? tmp24556 : tmp24729;
  assign tmp24724 = s7 ? tmp24725 : tmp24728;
  assign tmp24712 = s8 ? tmp24713 : tmp24724;
  assign tmp24700 = s9 ? tmp24701 : tmp24712;
  assign tmp24490 = s10 ? tmp24491 : tmp24700;
  assign tmp24734 = s7 ? tmp24555 : tmp24682;
  assign tmp24735 = s7 ? tmp24631 : tmp24703;
  assign tmp24733 = s8 ? tmp24734 : tmp24735;
  assign tmp24732 = s9 ? tmp24701 : tmp24733;
  assign tmp24731 = s10 ? tmp24491 : tmp24732;
  assign tmp24489 = s11 ? tmp24490 : tmp24731;
  assign tmp24744 = s1 ? tmp24536 : tmp24535;
  assign tmp24747 = s0 ? tmp24536 : tmp23982;
  assign tmp24746 = s1 ? tmp24747 : tmp24536;
  assign tmp24745 = s2 ? tmp24536 : tmp24746;
  assign tmp24743 = s3 ? tmp24744 : tmp24745;
  assign tmp24750 = s1 ? tmp24747 : tmp23982;
  assign tmp24749 = s2 ? tmp24746 : tmp24750;
  assign tmp24753 = s0 ? tmp23982 : tmp24514;
  assign tmp24752 = s1 ? tmp23982 : tmp24753;
  assign tmp24751 = s2 ? tmp24752 : tmp24536;
  assign tmp24748 = s3 ? tmp24749 : tmp24751;
  assign tmp24742 = s4 ? tmp24743 : tmp24748;
  assign tmp24758 = s1 ? tmp24747 : tmp24535;
  assign tmp24759 = s1 ? tmp24535 : tmp24747;
  assign tmp24757 = s2 ? tmp24758 : tmp24759;
  assign tmp24760 = s2 ? tmp24535 : tmp24579;
  assign tmp24756 = s3 ? tmp24757 : tmp24760;
  assign tmp24763 = s1 ? tmp24549 : tmp23982;
  assign tmp24764 = s1 ? tmp23982 : tmp24747;
  assign tmp24762 = s2 ? tmp24763 : tmp24764;
  assign tmp24765 = s2 ? tmp24744 : tmp24514;
  assign tmp24761 = s3 ? tmp24762 : tmp24765;
  assign tmp24755 = s4 ? tmp24756 : tmp24761;
  assign tmp24768 = s2 ? tmp24546 : tmp24536;
  assign tmp24767 = s3 ? tmp24768 : tmp24545;
  assign tmp24771 = s1 ? tmp24549 : tmp24536;
  assign tmp24770 = s2 ? tmp24536 : tmp24771;
  assign tmp24769 = s3 ? tmp24770 : tmp24553;
  assign tmp24766 = s4 ? tmp24767 : tmp24769;
  assign tmp24754 = s5 ? tmp24755 : tmp24766;
  assign tmp24741 = s6 ? tmp24742 : tmp24754;
  assign tmp24776 = s1 ? tmp23982 : tmp24514;
  assign tmp24775 = s2 ? tmp24776 : tmp24536;
  assign tmp24774 = s3 ? tmp24749 : tmp24775;
  assign tmp24773 = s4 ? tmp24743 : tmp24774;
  assign tmp24781 = s1 ? tmp24536 : tmp24747;
  assign tmp24780 = s2 ? tmp24746 : tmp24781;
  assign tmp24782 = s2 ? tmp24536 : tmp24579;
  assign tmp24779 = s3 ? tmp24780 : tmp24782;
  assign tmp24784 = s2 ? tmp24763 : tmp24536;
  assign tmp24785 = s2 ? tmp24536 : tmp24514;
  assign tmp24783 = s3 ? tmp24784 : tmp24785;
  assign tmp24778 = s4 ? tmp24779 : tmp24783;
  assign tmp24787 = s3 ? tmp24768 : tmp24576;
  assign tmp24789 = s2 ? tmp24536 : tmp24527;
  assign tmp24788 = s3 ? tmp24789 : tmp24536;
  assign tmp24786 = s4 ? tmp24787 : tmp24788;
  assign tmp24777 = s5 ? tmp24778 : tmp24786;
  assign tmp24772 = s6 ? tmp24773 : tmp24777;
  assign tmp24740 = s7 ? tmp24741 : tmp24772;
  assign tmp24795 = s1 ? tmp24547 : tmp24536;
  assign tmp24794 = s2 ? tmp24536 : tmp24795;
  assign tmp24793 = s3 ? tmp24744 : tmp24794;
  assign tmp24792 = s4 ? tmp24793 : tmp24748;
  assign tmp24800 = s1 ? tmp24535 : tmp24547;
  assign tmp24799 = s2 ? tmp24758 : tmp24800;
  assign tmp24801 = s2 ? tmp24549 : tmp24579;
  assign tmp24798 = s3 ? tmp24799 : tmp24801;
  assign tmp24797 = s4 ? tmp24798 : tmp24761;
  assign tmp24804 = s2 ? tmp24628 : tmp24771;
  assign tmp24803 = s3 ? tmp24804 : tmp24553;
  assign tmp24802 = s4 ? tmp24767 : tmp24803;
  assign tmp24796 = s5 ? tmp24797 : tmp24802;
  assign tmp24791 = s6 ? tmp24792 : tmp24796;
  assign tmp24806 = s4 ? tmp24793 : tmp24774;
  assign tmp24811 = s1 ? tmp24536 : tmp24547;
  assign tmp24810 = s2 ? tmp24746 : tmp24811;
  assign tmp24809 = s3 ? tmp24810 : tmp24782;
  assign tmp24808 = s4 ? tmp24809 : tmp24783;
  assign tmp24815 = s1 ? tmp24536 : tmp24527;
  assign tmp24814 = s2 ? tmp24514 : tmp24815;
  assign tmp24813 = s3 ? tmp24814 : tmp24536;
  assign tmp24812 = s4 ? tmp24787 : tmp24813;
  assign tmp24807 = s5 ? tmp24808 : tmp24812;
  assign tmp24805 = s6 ? tmp24806 : tmp24807;
  assign tmp24790 = s7 ? tmp24791 : tmp24805;
  assign tmp24739 = s8 ? tmp24740 : tmp24790;
  assign tmp24823 = s1 ? tmp24535 : tmp24536;
  assign tmp24822 = s2 ? tmp24758 : tmp24823;
  assign tmp24821 = s3 ? tmp24822 : tmp24782;
  assign tmp24820 = s4 ? tmp24821 : tmp24761;
  assign tmp24819 = s5 ? tmp24820 : tmp24766;
  assign tmp24818 = s6 ? tmp24742 : tmp24819;
  assign tmp24828 = s2 ? tmp24746 : tmp24536;
  assign tmp24827 = s3 ? tmp24828 : tmp24782;
  assign tmp24826 = s4 ? tmp24827 : tmp24783;
  assign tmp24830 = s3 ? tmp24768 : tmp24696;
  assign tmp24829 = s4 ? tmp24830 : tmp24536;
  assign tmp24825 = s5 ? tmp24826 : tmp24829;
  assign tmp24824 = s6 ? tmp24773 : tmp24825;
  assign tmp24817 = s7 ? tmp24818 : tmp24824;
  assign tmp24816 = s8 ? tmp24790 : tmp24817;
  assign tmp24738 = s9 ? tmp24739 : tmp24816;
  assign tmp24835 = s5 ? tmp24826 : tmp24786;
  assign tmp24834 = s6 ? tmp24773 : tmp24835;
  assign tmp24833 = s7 ? tmp24818 : tmp24834;
  assign tmp24832 = s8 ? tmp24833 : tmp24818;
  assign tmp24842 = s2 ? tmp24514 : tmp24536;
  assign tmp24841 = s3 ? tmp24842 : tmp24536;
  assign tmp24840 = s4 ? tmp24787 : tmp24841;
  assign tmp24839 = s5 ? tmp24778 : tmp24840;
  assign tmp24838 = s6 ? tmp24773 : tmp24839;
  assign tmp24845 = s4 ? tmp24830 : tmp24841;
  assign tmp24844 = s5 ? tmp24778 : tmp24845;
  assign tmp24843 = s6 ? tmp24773 : tmp24844;
  assign tmp24837 = s7 ? tmp24838 : tmp24843;
  assign tmp24848 = s5 ? tmp24808 : tmp24840;
  assign tmp24847 = s6 ? tmp24806 : tmp24848;
  assign tmp24850 = s5 ? tmp24826 : tmp24840;
  assign tmp24849 = s6 ? tmp24773 : tmp24850;
  assign tmp24846 = s7 ? tmp24847 : tmp24849;
  assign tmp24836 = s8 ? tmp24837 : tmp24846;
  assign tmp24831 = s9 ? tmp24832 : tmp24836;
  assign tmp24737 = s10 ? tmp24738 : tmp24831;
  assign tmp24856 = s5 ? tmp24778 : tmp24829;
  assign tmp24855 = s6 ? tmp24773 : tmp24856;
  assign tmp24854 = s7 ? tmp24772 : tmp24855;
  assign tmp24857 = s7 ? tmp24805 : tmp24834;
  assign tmp24853 = s8 ? tmp24854 : tmp24857;
  assign tmp24852 = s9 ? tmp24832 : tmp24853;
  assign tmp24851 = s10 ? tmp24738 : tmp24852;
  assign tmp24736 = s11 ? tmp24737 : tmp24851;
  assign tmp24488 = s12 ? tmp24489 : tmp24736;
  assign tmp24341 = s13 ? tmp24342 : tmp24488;
  assign tmp23954 = s14 ? tmp23955 : tmp24341;
  assign tmp24869 = l3 ? tmp23968 : 1;
  assign tmp24868 = l1 ? tmp24869 : 1;
  assign tmp24871 = l2 ? 1 : tmp24869;
  assign tmp24870 = l1 ? tmp24871 : 1;
  assign tmp24867 = s1 ? tmp24868 : tmp24870;
  assign tmp24875 = l2 ? tmp24869 : 1;
  assign tmp24874 = l1 ? tmp24869 : tmp24875;
  assign tmp24873 = s0 ? tmp24870 : tmp24874;
  assign tmp24876 = s1 ? tmp24870 : tmp24874;
  assign tmp24872 = s2 ? tmp24873 : tmp24876;
  assign tmp24866 = s3 ? tmp24867 : tmp24872;
  assign tmp24880 = s0 ? tmp24868 : tmp24870;
  assign tmp24879 = s1 ? tmp24880 : tmp24870;
  assign tmp24878 = s2 ? tmp24876 : tmp24879;
  assign tmp24882 = s1 ? tmp24870 : tmp24873;
  assign tmp24881 = s2 ? tmp24882 : tmp24874;
  assign tmp24877 = s3 ? tmp24878 : tmp24881;
  assign tmp24865 = s4 ? tmp24866 : tmp24877;
  assign tmp24888 = s0 ? tmp24874 : tmp24870;
  assign tmp24887 = s1 ? tmp24870 : tmp24888;
  assign tmp24886 = s2 ? tmp24870 : tmp24887;
  assign tmp24885 = s3 ? tmp24886 : tmp24881;
  assign tmp24891 = s1 ? tmp24874 : tmp24870;
  assign tmp24890 = s2 ? tmp24891 : tmp24870;
  assign tmp24894 = s0 ? tmp24870 : tmp24868;
  assign tmp24893 = s1 ? tmp24894 : tmp24873;
  assign tmp24892 = s2 ? tmp24893 : tmp24874;
  assign tmp24889 = s3 ? tmp24890 : tmp24892;
  assign tmp24884 = s4 ? tmp24885 : tmp24889;
  assign tmp24898 = s1 ? tmp24874 : tmp24888;
  assign tmp24897 = s2 ? tmp24898 : tmp24870;
  assign tmp24902 = l1 ? tmp24871 : tmp24875;
  assign tmp24901 = s0 ? tmp24870 : tmp24902;
  assign tmp24900 = s1 ? tmp24870 : tmp24901;
  assign tmp24904 = s0 ? tmp24902 : tmp24868;
  assign tmp24903 = s1 ? tmp24904 : tmp24880;
  assign tmp24899 = s2 ? tmp24900 : tmp24903;
  assign tmp24896 = s3 ? tmp24897 : tmp24899;
  assign tmp24907 = s1 ? tmp24888 : tmp24870;
  assign tmp24906 = s2 ? tmp24882 : tmp24907;
  assign tmp24909 = s1 ? tmp24902 : tmp24904;
  assign tmp24908 = s2 ? tmp24909 : tmp24879;
  assign tmp24905 = s3 ? tmp24906 : tmp24908;
  assign tmp24895 = s4 ? tmp24896 : tmp24905;
  assign tmp24883 = s5 ? tmp24884 : tmp24895;
  assign tmp24864 = s6 ? tmp24865 : tmp24883;
  assign tmp24913 = s2 ? tmp24876 : tmp24874;
  assign tmp24912 = s3 ? tmp24878 : tmp24913;
  assign tmp24911 = s4 ? tmp24866 : tmp24912;
  assign tmp24916 = s3 ? tmp24886 : tmp24913;
  assign tmp24919 = s1 ? tmp24894 : tmp24874;
  assign tmp24918 = s2 ? tmp24919 : tmp24874;
  assign tmp24917 = s3 ? tmp24890 : tmp24918;
  assign tmp24915 = s4 ? tmp24916 : tmp24917;
  assign tmp24923 = s1 ? tmp24870 : tmp24902;
  assign tmp24922 = s2 ? tmp24923 : tmp24867;
  assign tmp24921 = s3 ? tmp24897 : tmp24922;
  assign tmp24925 = s2 ? tmp24876 : tmp24888;
  assign tmp24926 = s1 ? tmp24902 : tmp24868;
  assign tmp24924 = s3 ? tmp24925 : tmp24926;
  assign tmp24920 = s4 ? tmp24921 : tmp24924;
  assign tmp24914 = s5 ? tmp24915 : tmp24920;
  assign tmp24910 = s6 ? tmp24911 : tmp24914;
  assign tmp24863 = s7 ? tmp24864 : tmp24910;
  assign tmp24928 = s8 ? tmp24863 : tmp24864;
  assign tmp24933 = s2 ? tmp24876 : tmp24870;
  assign tmp24932 = s3 ? tmp24933 : tmp24926;
  assign tmp24931 = s4 ? tmp24921 : tmp24932;
  assign tmp24930 = s5 ? tmp24915 : tmp24931;
  assign tmp24929 = s6 ? tmp24911 : tmp24930;
  assign tmp24927 = s9 ? tmp24928 : tmp24929;
  assign tmp24862 = s10 ? tmp24863 : tmp24927;
  assign tmp24935 = s9 ? tmp24928 : tmp24910;
  assign tmp24934 = s10 ? tmp24863 : tmp24935;
  assign tmp24861 = s11 ? tmp24862 : tmp24934;
  assign tmp24942 = l1 ? tmp24875 : tmp24871;
  assign tmp24943 = l1 ? 1 : tmp24871;
  assign tmp24941 = s1 ? tmp24942 : tmp24943;
  assign tmp24946 = l1 ? tmp24875 : tmp24869;
  assign tmp24945 = s0 ? tmp24942 : tmp24946;
  assign tmp24948 = s0 ? tmp24946 : tmp24942;
  assign tmp24947 = s1 ? tmp24942 : tmp24948;
  assign tmp24944 = s2 ? tmp24945 : tmp24947;
  assign tmp24940 = s3 ? tmp24941 : tmp24944;
  assign tmp24951 = s1 ? tmp24942 : tmp24945;
  assign tmp24950 = s2 ? tmp24951 : tmp24942;
  assign tmp24952 = s2 ? tmp24951 : tmp24946;
  assign tmp24949 = s3 ? tmp24950 : tmp24952;
  assign tmp24939 = s4 ? tmp24940 : tmp24949;
  assign tmp24958 = s0 ? tmp24946 : tmp24875;
  assign tmp24957 = s1 ? tmp24943 : tmp24958;
  assign tmp24956 = s2 ? tmp24943 : tmp24957;
  assign tmp24961 = s0 ? tmp24875 : tmp24946;
  assign tmp24960 = s1 ? tmp24942 : tmp24961;
  assign tmp24959 = s2 ? tmp24960 : tmp24946;
  assign tmp24955 = s3 ? tmp24956 : tmp24959;
  assign tmp24964 = s1 ? tmp24948 : tmp24942;
  assign tmp24963 = s2 ? tmp24964 : tmp24942;
  assign tmp24962 = s3 ? tmp24963 : tmp24952;
  assign tmp24954 = s4 ? tmp24955 : tmp24962;
  assign tmp24969 = s0 ? tmp24875 : tmp24942;
  assign tmp24968 = s1 ? tmp24946 : tmp24969;
  assign tmp24967 = s2 ? tmp24968 : tmp24942;
  assign tmp24973 = l1 ? 1 : tmp24869;
  assign tmp24972 = s0 ? tmp24943 : tmp24973;
  assign tmp24971 = s1 ? tmp24943 : tmp24972;
  assign tmp24975 = s0 ? tmp24973 : tmp24942;
  assign tmp24974 = s1 ? tmp24975 : tmp24942;
  assign tmp24970 = s2 ? tmp24971 : tmp24974;
  assign tmp24966 = s3 ? tmp24967 : tmp24970;
  assign tmp24979 = s0 ? tmp24943 : tmp24946;
  assign tmp24978 = s1 ? tmp24943 : tmp24979;
  assign tmp24981 = s0 ? tmp24875 : tmp24943;
  assign tmp24980 = s1 ? tmp24981 : tmp24943;
  assign tmp24977 = s2 ? tmp24978 : tmp24980;
  assign tmp24983 = s1 ? tmp24972 : tmp24975;
  assign tmp24985 = s0 ? tmp24942 : tmp24943;
  assign tmp24984 = s1 ? tmp24985 : tmp24943;
  assign tmp24982 = s2 ? tmp24983 : tmp24984;
  assign tmp24976 = s3 ? tmp24977 : tmp24982;
  assign tmp24965 = s4 ? tmp24966 : tmp24976;
  assign tmp24953 = s5 ? tmp24954 : tmp24965;
  assign tmp24938 = s6 ? tmp24939 : tmp24953;
  assign tmp24990 = s1 ? tmp24942 : tmp24946;
  assign tmp24989 = s2 ? tmp24990 : tmp24946;
  assign tmp24988 = s3 ? tmp24950 : tmp24989;
  assign tmp24987 = s4 ? tmp24940 : tmp24988;
  assign tmp24993 = s3 ? tmp24956 : tmp24989;
  assign tmp24994 = s3 ? tmp24963 : tmp24989;
  assign tmp24992 = s4 ? tmp24993 : tmp24994;
  assign tmp24998 = s1 ? tmp24946 : tmp24942;
  assign tmp24997 = s2 ? tmp24998 : tmp24942;
  assign tmp25000 = s1 ? tmp24943 : tmp24973;
  assign tmp24999 = s2 ? tmp25000 : tmp24942;
  assign tmp24996 = s3 ? tmp24997 : tmp24999;
  assign tmp25003 = s1 ? tmp24943 : tmp24946;
  assign tmp25002 = s2 ? tmp25003 : tmp24943;
  assign tmp25004 = s1 ? tmp24973 : tmp24942;
  assign tmp25001 = s3 ? tmp25002 : tmp25004;
  assign tmp24995 = s4 ? tmp24996 : tmp25001;
  assign tmp24991 = s5 ? tmp24992 : tmp24995;
  assign tmp24986 = s6 ? tmp24987 : tmp24991;
  assign tmp24937 = s7 ? tmp24938 : tmp24986;
  assign tmp25006 = s8 ? tmp24937 : tmp24938;
  assign tmp25005 = s9 ? tmp25006 : tmp24986;
  assign tmp24936 = s10 ? tmp24937 : tmp25005;
  assign tmp24860 = s12 ? tmp24861 : tmp24936;
  assign tmp25018 = l2 ? tmp24401 : tmp23968;
  assign tmp25017 = l1 ? tmp24869 : tmp25018;
  assign tmp25020 = l1 ? 1 : tmp24401;
  assign tmp25021 = l1 ? tmp24871 : tmp24401;
  assign tmp25019 = s0 ? tmp25020 : tmp25021;
  assign tmp25016 = s1 ? tmp25017 : tmp25019;
  assign tmp25024 = s0 ? tmp24410 : tmp25017;
  assign tmp25026 = l1 ? tmp24871 : tmp24400;
  assign tmp25025 = s0 ? tmp25026 : tmp25017;
  assign tmp25023 = s1 ? tmp25024 : tmp25025;
  assign tmp25028 = s0 ? tmp25026 : tmp24410;
  assign tmp25027 = s1 ? tmp25028 : tmp25017;
  assign tmp25022 = s2 ? tmp25023 : tmp25027;
  assign tmp25015 = s3 ? tmp25016 : tmp25022;
  assign tmp25032 = s0 ? tmp25020 : tmp24410;
  assign tmp25031 = s1 ? tmp25032 : tmp25017;
  assign tmp25034 = s0 ? tmp25017 : tmp24410;
  assign tmp25033 = s1 ? tmp25034 : tmp24410;
  assign tmp25030 = s2 ? tmp25031 : tmp25033;
  assign tmp25036 = s1 ? tmp24410 : tmp25024;
  assign tmp25035 = s2 ? tmp25036 : tmp25017;
  assign tmp25029 = s3 ? tmp25030 : tmp25035;
  assign tmp25014 = s4 ? tmp25015 : tmp25029;
  assign tmp25042 = s0 ? tmp25021 : tmp25020;
  assign tmp25041 = s1 ? tmp25042 : tmp24410;
  assign tmp25043 = s1 ? tmp25019 : tmp25034;
  assign tmp25040 = s2 ? tmp25041 : tmp25043;
  assign tmp25046 = s0 ? tmp24410 : tmp25026;
  assign tmp25045 = s1 ? tmp25046 : tmp25024;
  assign tmp25050 = l2 ? 1 : tmp23968;
  assign tmp25049 = l1 ? tmp24869 : tmp25050;
  assign tmp25048 = s0 ? tmp25017 : tmp25049;
  assign tmp25047 = s1 ? tmp25048 : tmp25017;
  assign tmp25044 = s2 ? tmp25045 : tmp25047;
  assign tmp25039 = s3 ? tmp25040 : tmp25044;
  assign tmp25053 = s1 ? tmp25017 : tmp24410;
  assign tmp25054 = s1 ? tmp24410 : tmp25032;
  assign tmp25052 = s2 ? tmp25053 : tmp25054;
  assign tmp25056 = s0 ? tmp25020 : tmp25017;
  assign tmp25058 = l1 ? tmp24875 : tmp25050;
  assign tmp25059 = s0 ? tmp25017 : tmp25058;
  assign tmp25057 = s1 ? tmp25058 : tmp25059;
  assign tmp25055 = s2 ? tmp25056 : tmp25057;
  assign tmp25051 = s3 ? tmp25052 : tmp25055;
  assign tmp25038 = s4 ? tmp25039 : tmp25051;
  assign tmp25065 = l1 ? tmp24869 : tmp24401;
  assign tmp25064 = s0 ? tmp25017 : tmp25065;
  assign tmp25066 = s0 ? tmp24868 : tmp25026;
  assign tmp25063 = s1 ? tmp25064 : tmp25066;
  assign tmp25067 = s1 ? tmp25028 : tmp24410;
  assign tmp25062 = s2 ? tmp25063 : tmp25067;
  assign tmp25072 = l2 ? 1 : tmp24401;
  assign tmp25071 = l1 ? 1 : tmp25072;
  assign tmp25073 = l1 ? 1 : tmp25050;
  assign tmp25070 = s0 ? tmp25071 : tmp25073;
  assign tmp25074 = s0 ? tmp25073 : tmp24871;
  assign tmp25069 = s1 ? tmp25070 : tmp25074;
  assign tmp25077 = l1 ? tmp24871 : tmp25050;
  assign tmp25076 = s0 ? tmp25077 : tmp25017;
  assign tmp25078 = s0 ? tmp25017 : tmp25020;
  assign tmp25075 = s1 ? tmp25076 : tmp25078;
  assign tmp25068 = s2 ? tmp25069 : tmp25075;
  assign tmp25061 = s3 ? tmp25062 : tmp25068;
  assign tmp25083 = l1 ? tmp24871 : tmp25072;
  assign tmp25082 = s0 ? tmp25020 : tmp25083;
  assign tmp25084 = s0 ? tmp25083 : tmp25017;
  assign tmp25081 = s1 ? tmp25082 : tmp25084;
  assign tmp25086 = s0 ? tmp24868 : tmp25021;
  assign tmp25085 = s1 ? tmp25086 : tmp24410;
  assign tmp25080 = s2 ? tmp25081 : tmp25085;
  assign tmp25089 = s0 ? tmp25026 : tmp25077;
  assign tmp25088 = s1 ? tmp25089 : tmp25076;
  assign tmp25091 = s0 ? tmp25073 : tmp25083;
  assign tmp25090 = s1 ? tmp25078 : tmp25091;
  assign tmp25087 = s2 ? tmp25088 : tmp25090;
  assign tmp25079 = s3 ? tmp25080 : tmp25087;
  assign tmp25060 = s4 ? tmp25061 : tmp25079;
  assign tmp25037 = s5 ? tmp25038 : tmp25060;
  assign tmp25013 = s6 ? tmp25014 : tmp25037;
  assign tmp25096 = s1 ? tmp24410 : tmp25017;
  assign tmp25095 = s2 ? tmp25096 : tmp25017;
  assign tmp25094 = s3 ? tmp25030 : tmp25095;
  assign tmp25093 = s4 ? tmp25015 : tmp25094;
  assign tmp25101 = s1 ? tmp25021 : tmp25034;
  assign tmp25100 = s2 ? tmp25041 : tmp25101;
  assign tmp25103 = s1 ? tmp25026 : tmp25017;
  assign tmp25102 = s2 ? tmp25103 : tmp25047;
  assign tmp25099 = s3 ? tmp25100 : tmp25102;
  assign tmp25105 = s2 ? tmp25053 : tmp25020;
  assign tmp25107 = s1 ? tmp25056 : tmp25017;
  assign tmp25108 = s1 ? tmp25058 : tmp25017;
  assign tmp25106 = s2 ? tmp25107 : tmp25108;
  assign tmp25104 = s3 ? tmp25105 : tmp25106;
  assign tmp25098 = s4 ? tmp25099 : tmp25104;
  assign tmp25112 = s1 ? tmp25064 : tmp25026;
  assign tmp25111 = s2 ? tmp25112 : tmp24410;
  assign tmp25114 = s1 ? tmp25073 : tmp24871;
  assign tmp25115 = s1 ? tmp25017 : tmp25078;
  assign tmp25113 = s2 ? tmp25114 : tmp25115;
  assign tmp25110 = s3 ? tmp25111 : tmp25113;
  assign tmp25118 = s1 ? tmp25083 : tmp25017;
  assign tmp25117 = s2 ? tmp25118 : tmp25021;
  assign tmp25120 = s1 ? tmp25077 : tmp25017;
  assign tmp25119 = s2 ? tmp25120 : tmp25017;
  assign tmp25116 = s3 ? tmp25117 : tmp25119;
  assign tmp25109 = s4 ? tmp25110 : tmp25116;
  assign tmp25097 = s5 ? tmp25098 : tmp25109;
  assign tmp25092 = s6 ? tmp25093 : tmp25097;
  assign tmp25012 = s7 ? tmp25013 : tmp25092;
  assign tmp25126 = s1 ? tmp25020 : tmp25017;
  assign tmp25125 = s2 ? tmp25126 : tmp25033;
  assign tmp25124 = s3 ? tmp25125 : tmp25035;
  assign tmp25123 = s4 ? tmp25015 : tmp25124;
  assign tmp25131 = s1 ? tmp24410 : tmp25020;
  assign tmp25130 = s2 ? tmp25053 : tmp25131;
  assign tmp25129 = s3 ? tmp25130 : tmp25055;
  assign tmp25128 = s4 ? tmp25039 : tmp25129;
  assign tmp25127 = s5 ? tmp25128 : tmp25060;
  assign tmp25122 = s6 ? tmp25123 : tmp25127;
  assign tmp25134 = s3 ? tmp25125 : tmp25095;
  assign tmp25133 = s4 ? tmp25015 : tmp25134;
  assign tmp25132 = s6 ? tmp25133 : tmp25097;
  assign tmp25121 = s7 ? tmp25122 : tmp25132;
  assign tmp25011 = s8 ? tmp25012 : tmp25121;
  assign tmp25142 = s1 ? tmp25086 : tmp25020;
  assign tmp25141 = s2 ? tmp25081 : tmp25142;
  assign tmp25140 = s3 ? tmp25141 : tmp25087;
  assign tmp25139 = s4 ? tmp25061 : tmp25140;
  assign tmp25138 = s5 ? tmp25128 : tmp25139;
  assign tmp25137 = s6 ? tmp25123 : tmp25138;
  assign tmp25148 = s1 ? tmp25020 : tmp24410;
  assign tmp25147 = s2 ? tmp25112 : tmp25148;
  assign tmp25146 = s3 ? tmp25147 : tmp25113;
  assign tmp25145 = s4 ? tmp25146 : tmp25116;
  assign tmp25144 = s5 ? tmp25098 : tmp25145;
  assign tmp25143 = s6 ? tmp25133 : tmp25144;
  assign tmp25136 = s7 ? tmp25137 : tmp25143;
  assign tmp25135 = s8 ? tmp25121 : tmp25136;
  assign tmp25010 = s9 ? tmp25011 : tmp25135;
  assign tmp25150 = s8 ? tmp25136 : tmp25137;
  assign tmp25156 = s3 ? tmp25117 : tmp25120;
  assign tmp25155 = s4 ? tmp25110 : tmp25156;
  assign tmp25154 = s5 ? tmp25098 : tmp25155;
  assign tmp25153 = s6 ? tmp25093 : tmp25154;
  assign tmp25159 = s4 ? tmp25146 : tmp25156;
  assign tmp25158 = s5 ? tmp25098 : tmp25159;
  assign tmp25157 = s6 ? tmp25133 : tmp25158;
  assign tmp25152 = s7 ? tmp25153 : tmp25157;
  assign tmp25161 = s6 ? tmp25133 : tmp25154;
  assign tmp25160 = s7 ? tmp25161 : tmp25157;
  assign tmp25151 = s8 ? tmp25152 : tmp25160;
  assign tmp25149 = s9 ? tmp25150 : tmp25151;
  assign tmp25009 = s10 ? tmp25010 : tmp25149;
  assign tmp25165 = s7 ? tmp25092 : tmp25143;
  assign tmp25166 = s7 ? tmp25132 : tmp25143;
  assign tmp25164 = s8 ? tmp25165 : tmp25166;
  assign tmp25163 = s9 ? tmp25150 : tmp25164;
  assign tmp25162 = s10 ? tmp25010 : tmp25163;
  assign tmp25008 = s11 ? tmp25009 : tmp25162;
  assign tmp25177 = l1 ? tmp25050 : 1;
  assign tmp25176 = s0 ? tmp24870 : tmp25177;
  assign tmp25175 = s1 ? tmp24871 : tmp25176;
  assign tmp25180 = l1 ? tmp25050 : tmp24869;
  assign tmp25179 = s0 ? tmp24870 : tmp25180;
  assign tmp25183 = l1 ? tmp25050 : tmp24871;
  assign tmp25182 = s0 ? tmp25180 : tmp25183;
  assign tmp25181 = s1 ? tmp24870 : tmp25182;
  assign tmp25178 = s2 ? tmp25179 : tmp25181;
  assign tmp25174 = s3 ? tmp25175 : tmp25178;
  assign tmp25187 = s0 ? tmp25183 : tmp25180;
  assign tmp25186 = s1 ? tmp24870 : tmp25187;
  assign tmp25189 = s0 ? tmp24871 : tmp24870;
  assign tmp25188 = s1 ? tmp25189 : tmp24870;
  assign tmp25185 = s2 ? tmp25186 : tmp25188;
  assign tmp25192 = s0 ? tmp25177 : tmp25180;
  assign tmp25191 = s1 ? tmp24870 : tmp25192;
  assign tmp25190 = s2 ? tmp25191 : tmp25180;
  assign tmp25184 = s3 ? tmp25185 : tmp25190;
  assign tmp25173 = s4 ? tmp25174 : tmp25184;
  assign tmp25197 = s1 ? tmp25177 : tmp24870;
  assign tmp25199 = s0 ? tmp25180 : tmp24870;
  assign tmp25198 = s1 ? tmp25177 : tmp25199;
  assign tmp25196 = s2 ? tmp25197 : tmp25198;
  assign tmp25201 = s1 ? tmp24870 : tmp25179;
  assign tmp25200 = s2 ? tmp25201 : tmp25180;
  assign tmp25195 = s3 ? tmp25196 : tmp25200;
  assign tmp25204 = s1 ? tmp25182 : tmp24870;
  assign tmp25203 = s2 ? tmp25204 : tmp24870;
  assign tmp25207 = s0 ? tmp24870 : tmp24871;
  assign tmp25206 = s1 ? tmp25207 : tmp25179;
  assign tmp25209 = s0 ? tmp25180 : tmp24973;
  assign tmp25208 = s1 ? tmp24973 : tmp25209;
  assign tmp25205 = s2 ? tmp25206 : tmp25208;
  assign tmp25202 = s3 ? tmp25203 : tmp25205;
  assign tmp25194 = s4 ? tmp25195 : tmp25202;
  assign tmp25215 = l1 ? tmp25050 : tmp24875;
  assign tmp25214 = s0 ? tmp25215 : tmp25183;
  assign tmp25213 = s1 ? tmp25180 : tmp25214;
  assign tmp25212 = s2 ? tmp25213 : tmp24870;
  assign tmp25219 = l1 ? tmp25072 : 1;
  assign tmp25220 = l1 ? tmp25072 : tmp24871;
  assign tmp25218 = s0 ? tmp25219 : tmp25220;
  assign tmp25221 = s0 ? tmp25220 : tmp25180;
  assign tmp25217 = s1 ? tmp25218 : tmp25221;
  assign tmp25222 = s1 ? tmp25182 : tmp25189;
  assign tmp25216 = s2 ? tmp25217 : tmp25222;
  assign tmp25211 = s3 ? tmp25212 : tmp25216;
  assign tmp25225 = s1 ? tmp25176 : tmp25187;
  assign tmp25227 = s0 ? tmp24902 : tmp25177;
  assign tmp25226 = s1 ? tmp25227 : tmp24870;
  assign tmp25224 = s2 ? tmp25225 : tmp25226;
  assign tmp25229 = s1 ? tmp25179 : tmp25182;
  assign tmp25231 = s0 ? tmp25220 : tmp25177;
  assign tmp25230 = s1 ? tmp25189 : tmp25231;
  assign tmp25228 = s2 ? tmp25229 : tmp25230;
  assign tmp25223 = s3 ? tmp25224 : tmp25228;
  assign tmp25210 = s4 ? tmp25211 : tmp25223;
  assign tmp25193 = s5 ? tmp25194 : tmp25210;
  assign tmp25172 = s6 ? tmp25173 : tmp25193;
  assign tmp25236 = s1 ? tmp24870 : tmp25180;
  assign tmp25235 = s2 ? tmp25236 : tmp25180;
  assign tmp25234 = s3 ? tmp25185 : tmp25235;
  assign tmp25233 = s4 ? tmp25174 : tmp25234;
  assign tmp25239 = s3 ? tmp25196 : tmp25235;
  assign tmp25242 = s1 ? tmp25207 : tmp25180;
  assign tmp25243 = s1 ? tmp24973 : tmp25180;
  assign tmp25241 = s2 ? tmp25242 : tmp25243;
  assign tmp25240 = s3 ? tmp25203 : tmp25241;
  assign tmp25238 = s4 ? tmp25239 : tmp25240;
  assign tmp25247 = s1 ? tmp25180 : tmp24870;
  assign tmp25246 = s2 ? tmp25247 : tmp24870;
  assign tmp25249 = s1 ? tmp25220 : tmp25180;
  assign tmp25248 = s2 ? tmp25249 : tmp25204;
  assign tmp25245 = s3 ? tmp25246 : tmp25248;
  assign tmp25252 = s1 ? tmp25183 : tmp25180;
  assign tmp25251 = s2 ? tmp25252 : tmp25177;
  assign tmp25253 = s1 ? tmp25180 : tmp25182;
  assign tmp25250 = s3 ? tmp25251 : tmp25253;
  assign tmp25244 = s4 ? tmp25245 : tmp25250;
  assign tmp25237 = s5 ? tmp25238 : tmp25244;
  assign tmp25232 = s6 ? tmp25233 : tmp25237;
  assign tmp25171 = s7 ? tmp25172 : tmp25232;
  assign tmp25257 = s3 ? tmp25185 : tmp25200;
  assign tmp25256 = s4 ? tmp25174 : tmp25257;
  assign tmp25255 = s6 ? tmp25256 : tmp25193;
  assign tmp25254 = s7 ? tmp25255 : tmp25232;
  assign tmp25170 = s8 ? tmp25171 : tmp25254;
  assign tmp25169 = s9 ? tmp25170 : tmp25254;
  assign tmp25259 = s8 ? tmp25254 : tmp25255;
  assign tmp25264 = s1 ? tmp25180 : tmp25183;
  assign tmp25263 = s3 ? tmp25251 : tmp25264;
  assign tmp25262 = s4 ? tmp25245 : tmp25263;
  assign tmp25261 = s5 ? tmp25238 : tmp25262;
  assign tmp25260 = s6 ? tmp25233 : tmp25261;
  assign tmp25258 = s9 ? tmp25259 : tmp25260;
  assign tmp25168 = s10 ? tmp25169 : tmp25258;
  assign tmp25266 = s9 ? tmp25259 : tmp25232;
  assign tmp25265 = s10 ? tmp25169 : tmp25266;
  assign tmp25167 = s11 ? tmp25168 : tmp25265;
  assign tmp25007 = s12 ? tmp25008 : tmp25167;
  assign tmp24859 = s13 ? tmp24860 : tmp25007;
  assign tmp25280 = l3 ? 1 : 0;
  assign tmp25279 = l2 ? tmp24401 : tmp25280;
  assign tmp25278 = l1 ? tmp24499 : tmp25279;
  assign tmp25281 = s0 ? tmp24399 : tmp25278;
  assign tmp25277 = s1 ? tmp25278 : tmp25281;
  assign tmp25286 = l2 ? 1 : tmp25280;
  assign tmp25285 = l1 ? tmp24499 : tmp25286;
  assign tmp25284 = s0 ? tmp25285 : tmp25278;
  assign tmp25283 = s1 ? tmp25284 : tmp25278;
  assign tmp25288 = s0 ? tmp24499 : tmp23982;
  assign tmp25287 = s1 ? tmp25288 : tmp25278;
  assign tmp25282 = s2 ? tmp25283 : tmp25287;
  assign tmp25276 = s3 ? tmp25277 : tmp25282;
  assign tmp25292 = s0 ? tmp25278 : tmp23982;
  assign tmp25291 = s1 ? tmp25292 : tmp25278;
  assign tmp25293 = s1 ? tmp25292 : tmp24404;
  assign tmp25290 = s2 ? tmp25291 : tmp25293;
  assign tmp25296 = s0 ? tmp23982 : tmp25020;
  assign tmp25295 = s1 ? tmp24399 : tmp25296;
  assign tmp25299 = l1 ? tmp24499 : tmp24401;
  assign tmp25298 = s0 ? tmp25299 : tmp25278;
  assign tmp25297 = s1 ? tmp25278 : tmp25298;
  assign tmp25294 = s2 ? tmp25295 : tmp25297;
  assign tmp25289 = s3 ? tmp25290 : tmp25294;
  assign tmp25275 = s4 ? tmp25276 : tmp25289;
  assign tmp25304 = s1 ? tmp25292 : tmp24535;
  assign tmp25306 = s0 ? tmp23982 : tmp25278;
  assign tmp25307 = s0 ? tmp25278 : tmp23983;
  assign tmp25305 = s1 ? tmp25306 : tmp25307;
  assign tmp25303 = s2 ? tmp25304 : tmp25305;
  assign tmp25309 = s0 ? tmp23983 : tmp25278;
  assign tmp25311 = s0 ? tmp25299 : tmp25071;
  assign tmp25310 = s1 ? tmp25311 : tmp25278;
  assign tmp25308 = s2 ? tmp25309 : tmp25310;
  assign tmp25302 = s3 ? tmp25303 : tmp25308;
  assign tmp25315 = s0 ? tmp25020 : tmp25278;
  assign tmp25317 = l1 ? tmp23983 : tmp25072;
  assign tmp25316 = s0 ? tmp25317 : tmp24399;
  assign tmp25314 = s1 ? tmp25315 : tmp25316;
  assign tmp25318 = s1 ? tmp25316 : tmp25292;
  assign tmp25313 = s2 ? tmp25314 : tmp25318;
  assign tmp25319 = s2 ? tmp25277 : tmp25020;
  assign tmp25312 = s3 ? tmp25313 : tmp25319;
  assign tmp25301 = s4 ? tmp25302 : tmp25312;
  assign tmp25324 = s0 ? tmp25278 : tmp25020;
  assign tmp25325 = s0 ? tmp24410 : tmp24400;
  assign tmp25323 = s1 ? tmp25324 : tmp25325;
  assign tmp25327 = s0 ? tmp24400 : tmp24536;
  assign tmp25326 = s1 ? tmp25327 : tmp24536;
  assign tmp25322 = s2 ? tmp25323 : tmp25326;
  assign tmp25330 = s0 ? tmp24536 : tmp25071;
  assign tmp25329 = s1 ? tmp25330 : tmp25071;
  assign tmp25332 = s0 ? tmp25071 : tmp25020;
  assign tmp25331 = s1 ? tmp25332 : tmp25315;
  assign tmp25328 = s2 ? tmp25329 : tmp25331;
  assign tmp25321 = s3 ? tmp25322 : tmp25328;
  assign tmp25337 = l1 ? tmp24400 : tmp25072;
  assign tmp25336 = s0 ? tmp25278 : tmp25337;
  assign tmp25338 = s0 ? tmp25337 : tmp25299;
  assign tmp25335 = s1 ? tmp25336 : tmp25338;
  assign tmp25339 = s1 ? tmp25315 : tmp24536;
  assign tmp25334 = s2 ? tmp25335 : tmp25339;
  assign tmp25342 = s0 ? tmp24400 : tmp25337;
  assign tmp25343 = s0 ? tmp25071 : tmp25278;
  assign tmp25341 = s1 ? tmp25342 : tmp25343;
  assign tmp25345 = s0 ? tmp25071 : tmp25337;
  assign tmp25344 = s1 ? tmp25315 : tmp25345;
  assign tmp25340 = s2 ? tmp25341 : tmp25344;
  assign tmp25333 = s3 ? tmp25334 : tmp25340;
  assign tmp25320 = s4 ? tmp25321 : tmp25333;
  assign tmp25300 = s5 ? tmp25301 : tmp25320;
  assign tmp25274 = s6 ? tmp25275 : tmp25300;
  assign tmp25350 = s1 ? tmp25292 : tmp24399;
  assign tmp25349 = s2 ? tmp25291 : tmp25350;
  assign tmp25353 = l1 ? tmp23983 : tmp24401;
  assign tmp25352 = s1 ? tmp25353 : tmp25020;
  assign tmp25351 = s2 ? tmp25352 : tmp25297;
  assign tmp25348 = s3 ? tmp25349 : tmp25351;
  assign tmp25347 = s4 ? tmp25276 : tmp25348;
  assign tmp25358 = s1 ? tmp25292 : tmp24536;
  assign tmp25359 = s1 ? tmp25278 : tmp25307;
  assign tmp25357 = s2 ? tmp25358 : tmp25359;
  assign tmp25360 = s2 ? tmp25278 : tmp25310;
  assign tmp25356 = s3 ? tmp25357 : tmp25360;
  assign tmp25363 = s1 ? tmp24399 : tmp25278;
  assign tmp25362 = s2 ? tmp25314 : tmp25363;
  assign tmp25361 = s3 ? tmp25362 : tmp25319;
  assign tmp25355 = s4 ? tmp25356 : tmp25361;
  assign tmp25367 = s1 ? tmp25324 : tmp24400;
  assign tmp25366 = s2 ? tmp25367 : tmp24536;
  assign tmp25370 = s0 ? tmp24527 : tmp25071;
  assign tmp25369 = s1 ? tmp25370 : tmp25071;
  assign tmp25371 = s1 ? tmp25020 : tmp25278;
  assign tmp25368 = s2 ? tmp25369 : tmp25371;
  assign tmp25365 = s3 ? tmp25366 : tmp25368;
  assign tmp25374 = s1 ? tmp25336 : tmp25299;
  assign tmp25375 = s1 ? tmp25278 : tmp25285;
  assign tmp25373 = s2 ? tmp25374 : tmp25375;
  assign tmp25377 = s1 ? tmp25337 : tmp25278;
  assign tmp25376 = s2 ? tmp25377 : tmp25278;
  assign tmp25372 = s3 ? tmp25373 : tmp25376;
  assign tmp25364 = s4 ? tmp25365 : tmp25372;
  assign tmp25354 = s5 ? tmp25355 : tmp25364;
  assign tmp25346 = s6 ? tmp25347 : tmp25354;
  assign tmp25273 = s7 ? tmp25274 : tmp25346;
  assign tmp25385 = l1 ? tmp24499 : tmp24400;
  assign tmp25384 = s0 ? tmp25385 : tmp24514;
  assign tmp25383 = s1 ? tmp25384 : tmp25278;
  assign tmp25382 = s2 ? tmp25278 : tmp25383;
  assign tmp25381 = s3 ? tmp25277 : tmp25382;
  assign tmp25380 = s4 ? tmp25381 : tmp25289;
  assign tmp25391 = s0 ? tmp25278 : tmp24514;
  assign tmp25390 = s1 ? tmp25306 : tmp25391;
  assign tmp25389 = s2 ? tmp25304 : tmp25390;
  assign tmp25393 = s0 ? tmp24514 : tmp25278;
  assign tmp25396 = l1 ? tmp24400 : tmp24401;
  assign tmp25395 = s0 ? tmp25396 : tmp25071;
  assign tmp25394 = s1 ? tmp25395 : tmp25278;
  assign tmp25392 = s2 ? tmp25393 : tmp25394;
  assign tmp25388 = s3 ? tmp25389 : tmp25392;
  assign tmp25399 = s1 ? tmp25315 : tmp24419;
  assign tmp25400 = s1 ? tmp24419 : tmp25292;
  assign tmp25398 = s2 ? tmp25399 : tmp25400;
  assign tmp25397 = s3 ? tmp25398 : tmp25319;
  assign tmp25387 = s4 ? tmp25388 : tmp25397;
  assign tmp25405 = s0 ? tmp25337 : tmp25396;
  assign tmp25404 = s1 ? tmp25336 : tmp25405;
  assign tmp25403 = s2 ? tmp25404 : tmp25339;
  assign tmp25402 = s3 ? tmp25403 : tmp25340;
  assign tmp25401 = s4 ? tmp25321 : tmp25402;
  assign tmp25386 = s5 ? tmp25387 : tmp25401;
  assign tmp25379 = s6 ? tmp25380 : tmp25386;
  assign tmp25410 = s1 ? tmp24399 : tmp25020;
  assign tmp25409 = s2 ? tmp25410 : tmp25297;
  assign tmp25408 = s3 ? tmp25349 : tmp25409;
  assign tmp25407 = s4 ? tmp25381 : tmp25408;
  assign tmp25415 = s1 ? tmp25278 : tmp25391;
  assign tmp25414 = s2 ? tmp25358 : tmp25415;
  assign tmp25416 = s2 ? tmp25278 : tmp25394;
  assign tmp25413 = s3 ? tmp25414 : tmp25416;
  assign tmp25418 = s2 ? tmp25399 : tmp25278;
  assign tmp25419 = s2 ? tmp25278 : tmp25020;
  assign tmp25417 = s3 ? tmp25418 : tmp25419;
  assign tmp25412 = s4 ? tmp25413 : tmp25417;
  assign tmp25423 = s1 ? tmp25336 : tmp25396;
  assign tmp25422 = s2 ? tmp25423 : tmp25375;
  assign tmp25421 = s3 ? tmp25422 : tmp25376;
  assign tmp25420 = s4 ? tmp25365 : tmp25421;
  assign tmp25411 = s5 ? tmp25412 : tmp25420;
  assign tmp25406 = s6 ? tmp25407 : tmp25411;
  assign tmp25378 = s7 ? tmp25379 : tmp25406;
  assign tmp25272 = s8 ? tmp25273 : tmp25378;
  assign tmp25430 = s0 ? tmp24399 : tmp25299;
  assign tmp25429 = s1 ? tmp25299 : tmp25430;
  assign tmp25433 = s0 ? tmp25299 : tmp23982;
  assign tmp25432 = s1 ? tmp25433 : tmp25299;
  assign tmp25431 = s2 ? tmp25299 : tmp25432;
  assign tmp25428 = s3 ? tmp25429 : tmp25431;
  assign tmp25436 = s1 ? tmp25433 : tmp24404;
  assign tmp25435 = s2 ? tmp25432 : tmp25436;
  assign tmp25437 = s2 ? tmp25295 : tmp25299;
  assign tmp25434 = s3 ? tmp25435 : tmp25437;
  assign tmp25427 = s4 ? tmp25428 : tmp25434;
  assign tmp25442 = s1 ? tmp25433 : tmp24535;
  assign tmp25444 = s0 ? tmp23982 : tmp25299;
  assign tmp25445 = s0 ? tmp25299 : tmp24499;
  assign tmp25443 = s1 ? tmp25444 : tmp25445;
  assign tmp25441 = s2 ? tmp25442 : tmp25443;
  assign tmp25447 = s0 ? tmp24499 : tmp25299;
  assign tmp25448 = s1 ? tmp25311 : tmp25299;
  assign tmp25446 = s2 ? tmp25447 : tmp25448;
  assign tmp25440 = s3 ? tmp25441 : tmp25446;
  assign tmp25452 = s0 ? tmp25020 : tmp25299;
  assign tmp25451 = s1 ? tmp25452 : tmp25316;
  assign tmp25453 = s1 ? tmp25316 : tmp25433;
  assign tmp25450 = s2 ? tmp25451 : tmp25453;
  assign tmp25454 = s2 ? tmp25429 : tmp25020;
  assign tmp25449 = s3 ? tmp25450 : tmp25454;
  assign tmp25439 = s4 ? tmp25440 : tmp25449;
  assign tmp25459 = s0 ? tmp25299 : tmp25020;
  assign tmp25458 = s1 ? tmp25459 : tmp25325;
  assign tmp25457 = s2 ? tmp25458 : tmp25326;
  assign tmp25461 = s1 ? tmp25332 : tmp25452;
  assign tmp25460 = s2 ? tmp25329 : tmp25461;
  assign tmp25456 = s3 ? tmp25457 : tmp25460;
  assign tmp25465 = s0 ? tmp25299 : tmp25337;
  assign tmp25464 = s1 ? tmp25465 : tmp25338;
  assign tmp25466 = s1 ? tmp25452 : tmp24536;
  assign tmp25463 = s2 ? tmp25464 : tmp25466;
  assign tmp25469 = s0 ? tmp25071 : tmp25299;
  assign tmp25468 = s1 ? tmp25342 : tmp25469;
  assign tmp25470 = s1 ? tmp25452 : tmp25345;
  assign tmp25467 = s2 ? tmp25468 : tmp25470;
  assign tmp25462 = s3 ? tmp25463 : tmp25467;
  assign tmp25455 = s4 ? tmp25456 : tmp25462;
  assign tmp25438 = s5 ? tmp25439 : tmp25455;
  assign tmp25426 = s6 ? tmp25427 : tmp25438;
  assign tmp25475 = s1 ? tmp25433 : tmp24399;
  assign tmp25474 = s2 ? tmp25432 : tmp25475;
  assign tmp25476 = s2 ? tmp25352 : tmp25299;
  assign tmp25473 = s3 ? tmp25474 : tmp25476;
  assign tmp25472 = s4 ? tmp25428 : tmp25473;
  assign tmp25481 = s1 ? tmp25433 : tmp24536;
  assign tmp25482 = s1 ? tmp25299 : tmp25445;
  assign tmp25480 = s2 ? tmp25481 : tmp25482;
  assign tmp25483 = s2 ? tmp25299 : tmp25448;
  assign tmp25479 = s3 ? tmp25480 : tmp25483;
  assign tmp25485 = s2 ? tmp25451 : tmp25299;
  assign tmp25486 = s2 ? tmp25299 : tmp25020;
  assign tmp25484 = s3 ? tmp25485 : tmp25486;
  assign tmp25478 = s4 ? tmp25479 : tmp25484;
  assign tmp25490 = s1 ? tmp25459 : tmp24400;
  assign tmp25489 = s2 ? tmp25490 : tmp24536;
  assign tmp25492 = s1 ? tmp25020 : tmp25299;
  assign tmp25491 = s2 ? tmp25329 : tmp25492;
  assign tmp25488 = s3 ? tmp25489 : tmp25491;
  assign tmp25495 = s1 ? tmp25465 : tmp25299;
  assign tmp25494 = s2 ? tmp25495 : tmp25299;
  assign tmp25497 = s1 ? tmp25337 : tmp25299;
  assign tmp25496 = s2 ? tmp25497 : tmp25299;
  assign tmp25493 = s3 ? tmp25494 : tmp25496;
  assign tmp25487 = s4 ? tmp25488 : tmp25493;
  assign tmp25477 = s5 ? tmp25478 : tmp25487;
  assign tmp25471 = s6 ? tmp25472 : tmp25477;
  assign tmp25425 = s7 ? tmp25426 : tmp25471;
  assign tmp25424 = s8 ? tmp25378 : tmp25425;
  assign tmp25271 = s9 ? tmp25272 : tmp25424;
  assign tmp25507 = s0 ? tmp25278 : tmp24499;
  assign tmp25506 = s1 ? tmp25306 : tmp25507;
  assign tmp25505 = s2 ? tmp25304 : tmp25506;
  assign tmp25509 = s0 ? tmp24499 : tmp25278;
  assign tmp25508 = s2 ? tmp25509 : tmp25310;
  assign tmp25504 = s3 ? tmp25505 : tmp25508;
  assign tmp25503 = s4 ? tmp25504 : tmp25312;
  assign tmp25502 = s5 ? tmp25503 : tmp25320;
  assign tmp25501 = s6 ? tmp25275 : tmp25502;
  assign tmp25515 = s1 ? tmp25278 : tmp25507;
  assign tmp25514 = s2 ? tmp25358 : tmp25515;
  assign tmp25513 = s3 ? tmp25514 : tmp25360;
  assign tmp25517 = s2 ? tmp25314 : tmp25278;
  assign tmp25516 = s3 ? tmp25517 : tmp25419;
  assign tmp25512 = s4 ? tmp25513 : tmp25516;
  assign tmp25511 = s5 ? tmp25512 : tmp25364;
  assign tmp25510 = s6 ? tmp25347 : tmp25511;
  assign tmp25500 = s7 ? tmp25501 : tmp25510;
  assign tmp25499 = s8 ? tmp25500 : tmp25501;
  assign tmp25523 = s3 ? tmp25362 : tmp25419;
  assign tmp25522 = s4 ? tmp25356 : tmp25523;
  assign tmp25526 = s2 ? tmp25374 : tmp25278;
  assign tmp25525 = s3 ? tmp25526 : tmp25377;
  assign tmp25524 = s4 ? tmp25365 : tmp25525;
  assign tmp25521 = s5 ? tmp25522 : tmp25524;
  assign tmp25520 = s6 ? tmp25347 : tmp25521;
  assign tmp25530 = s3 ? tmp25494 : tmp25497;
  assign tmp25529 = s4 ? tmp25488 : tmp25530;
  assign tmp25528 = s5 ? tmp25478 : tmp25529;
  assign tmp25527 = s6 ? tmp25472 : tmp25528;
  assign tmp25519 = s7 ? tmp25520 : tmp25527;
  assign tmp25536 = s2 ? tmp25423 : tmp25278;
  assign tmp25535 = s3 ? tmp25536 : tmp25377;
  assign tmp25534 = s4 ? tmp25365 : tmp25535;
  assign tmp25533 = s5 ? tmp25412 : tmp25534;
  assign tmp25532 = s6 ? tmp25407 : tmp25533;
  assign tmp25538 = s5 ? tmp25512 : tmp25524;
  assign tmp25537 = s6 ? tmp25347 : tmp25538;
  assign tmp25531 = s7 ? tmp25532 : tmp25537;
  assign tmp25518 = s8 ? tmp25519 : tmp25531;
  assign tmp25498 = s9 ? tmp25499 : tmp25518;
  assign tmp25270 = s10 ? tmp25271 : tmp25498;
  assign tmp25542 = s7 ? tmp25346 : tmp25471;
  assign tmp25543 = s7 ? tmp25406 : tmp25510;
  assign tmp25541 = s8 ? tmp25542 : tmp25543;
  assign tmp25540 = s9 ? tmp25499 : tmp25541;
  assign tmp25539 = s10 ? tmp25271 : tmp25540;
  assign tmp25269 = s11 ? tmp25270 : tmp25539;
  assign tmp25554 = l2 ? tmp24401 : tmp24869;
  assign tmp25553 = l1 ? tmp25554 : tmp24400;
  assign tmp25555 = s0 ? tmp24410 : tmp25553;
  assign tmp25552 = s1 ? tmp25553 : tmp25555;
  assign tmp25558 = s0 ? tmp24514 : tmp25553;
  assign tmp25557 = s1 ? tmp25558 : tmp25553;
  assign tmp25560 = s0 ? tmp25553 : tmp24410;
  assign tmp25559 = s1 ? tmp25560 : tmp25553;
  assign tmp25556 = s2 ? tmp25557 : tmp25559;
  assign tmp25551 = s3 ? tmp25552 : tmp25556;
  assign tmp25564 = s0 ? tmp24400 : 1;
  assign tmp25563 = s1 ? tmp25564 : tmp25553;
  assign tmp25565 = s1 ? tmp25560 : tmp24410;
  assign tmp25562 = s2 ? tmp25563 : tmp25565;
  assign tmp25567 = s1 ? tmp24410 : tmp25046;
  assign tmp25566 = s2 ? tmp25567 : tmp25553;
  assign tmp25561 = s3 ? tmp25562 : tmp25566;
  assign tmp25550 = s4 ? tmp25551 : tmp25561;
  assign tmp25573 = s0 ? tmp25553 : tmp24514;
  assign tmp25572 = s1 ? tmp25573 : tmp24514;
  assign tmp25574 = s1 ? tmp25558 : tmp25560;
  assign tmp25571 = s2 ? tmp25572 : tmp25574;
  assign tmp25577 = s0 ? tmp25553 : tmp24870;
  assign tmp25576 = s1 ? tmp25577 : tmp25553;
  assign tmp25575 = s2 ? tmp25555 : tmp25576;
  assign tmp25570 = s3 ? tmp25571 : tmp25575;
  assign tmp25581 = s0 ? tmp25026 : tmp25553;
  assign tmp25582 = s0 ? 1 : tmp24410;
  assign tmp25580 = s1 ? tmp25581 : tmp25582;
  assign tmp25583 = s1 ? tmp25582 : tmp25564;
  assign tmp25579 = s2 ? tmp25580 : tmp25583;
  assign tmp25586 = s0 ? tmp25026 : tmp24870;
  assign tmp25585 = s1 ? tmp24870 : tmp25586;
  assign tmp25584 = s2 ? tmp25552 : tmp25585;
  assign tmp25578 = s3 ? tmp25579 : tmp25584;
  assign tmp25569 = s4 ? tmp25570 : tmp25578;
  assign tmp25591 = s0 ? tmp24870 : tmp25553;
  assign tmp25590 = s1 ? tmp25577 : tmp25591;
  assign tmp25589 = s2 ? tmp25590 : tmp25572;
  assign tmp25594 = s0 ? tmp24514 : tmp24870;
  assign tmp25593 = s1 ? tmp25594 : tmp24870;
  assign tmp25596 = s0 ? tmp25026 : tmp24400;
  assign tmp25595 = s1 ? tmp25026 : tmp25596;
  assign tmp25592 = s2 ? tmp25593 : tmp25595;
  assign tmp25588 = s3 ? tmp25589 : tmp25592;
  assign tmp25601 = l1 ? tmp25554 : 1;
  assign tmp25600 = s0 ? tmp24400 : tmp25601;
  assign tmp25599 = s1 ? tmp25600 : tmp25553;
  assign tmp25602 = s1 ? tmp25591 : tmp24514;
  assign tmp25598 = s2 ? tmp25599 : tmp25602;
  assign tmp25604 = s1 ? tmp25553 : tmp25591;
  assign tmp25606 = s0 ? tmp24870 : tmp25601;
  assign tmp25605 = s1 ? tmp25596 : tmp25606;
  assign tmp25603 = s2 ? tmp25604 : tmp25605;
  assign tmp25597 = s3 ? tmp25598 : tmp25603;
  assign tmp25587 = s4 ? tmp25588 : tmp25597;
  assign tmp25568 = s5 ? tmp25569 : tmp25587;
  assign tmp25549 = s6 ? tmp25550 : tmp25568;
  assign tmp25611 = s1 ? tmp24410 : tmp25026;
  assign tmp25610 = s2 ? tmp25611 : tmp25553;
  assign tmp25609 = s3 ? tmp25562 : tmp25610;
  assign tmp25608 = s4 ? tmp25551 : tmp25609;
  assign tmp25616 = s1 ? tmp25553 : tmp25560;
  assign tmp25615 = s2 ? tmp25572 : tmp25616;
  assign tmp25617 = s2 ? tmp25553 : tmp25576;
  assign tmp25614 = s3 ? tmp25615 : tmp25617;
  assign tmp25619 = s2 ? tmp25580 : tmp24400;
  assign tmp25621 = s1 ? tmp24870 : tmp25026;
  assign tmp25620 = s2 ? tmp25553 : tmp25621;
  assign tmp25618 = s3 ? tmp25619 : tmp25620;
  assign tmp25613 = s4 ? tmp25614 : tmp25618;
  assign tmp25624 = s2 ? tmp25576 : tmp25572;
  assign tmp25626 = s1 ? tmp25026 : tmp24400;
  assign tmp25625 = s2 ? tmp24870 : tmp25626;
  assign tmp25623 = s3 ? tmp25624 : tmp25625;
  assign tmp25622 = s4 ? tmp25623 : tmp25553;
  assign tmp25612 = s5 ? tmp25613 : tmp25622;
  assign tmp25607 = s6 ? tmp25608 : tmp25612;
  assign tmp25548 = s7 ? tmp25549 : tmp25607;
  assign tmp25632 = s1 ? tmp25573 : tmp25553;
  assign tmp25631 = s2 ? tmp25557 : tmp25632;
  assign tmp25630 = s3 ? tmp25552 : tmp25631;
  assign tmp25636 = s0 ? tmp24400 : tmp24514;
  assign tmp25635 = s1 ? tmp25636 : tmp25553;
  assign tmp25634 = s2 ? tmp25635 : tmp25565;
  assign tmp25633 = s3 ? tmp25634 : tmp25566;
  assign tmp25629 = s4 ? tmp25630 : tmp25633;
  assign tmp25641 = s1 ? tmp25558 : tmp25573;
  assign tmp25640 = s2 ? tmp25572 : tmp25641;
  assign tmp25642 = s2 ? tmp25558 : tmp25576;
  assign tmp25639 = s3 ? tmp25640 : tmp25642;
  assign tmp25646 = s0 ? tmp24514 : tmp24410;
  assign tmp25645 = s1 ? tmp25581 : tmp25646;
  assign tmp25647 = s1 ? tmp25646 : tmp25636;
  assign tmp25644 = s2 ? tmp25645 : tmp25647;
  assign tmp25643 = s3 ? tmp25644 : tmp25584;
  assign tmp25638 = s4 ? tmp25639 : tmp25643;
  assign tmp25652 = s0 ? tmp25601 : tmp25553;
  assign tmp25651 = s1 ? tmp25600 : tmp25652;
  assign tmp25650 = s2 ? tmp25651 : tmp25602;
  assign tmp25655 = s0 ? tmp25553 : tmp25601;
  assign tmp25654 = s1 ? tmp25655 : tmp25591;
  assign tmp25653 = s2 ? tmp25654 : tmp25605;
  assign tmp25649 = s3 ? tmp25650 : tmp25653;
  assign tmp25648 = s4 ? tmp25588 : tmp25649;
  assign tmp25637 = s5 ? tmp25638 : tmp25648;
  assign tmp25628 = s6 ? tmp25629 : tmp25637;
  assign tmp25658 = s3 ? tmp25634 : tmp25610;
  assign tmp25657 = s4 ? tmp25630 : tmp25658;
  assign tmp25663 = s1 ? tmp25553 : tmp25573;
  assign tmp25662 = s2 ? tmp25572 : tmp25663;
  assign tmp25661 = s3 ? tmp25662 : tmp25617;
  assign tmp25665 = s2 ? tmp25645 : tmp24400;
  assign tmp25664 = s3 ? tmp25665 : tmp25620;
  assign tmp25660 = s4 ? tmp25661 : tmp25664;
  assign tmp25668 = s2 ? tmp25576 : tmp24514;
  assign tmp25667 = s3 ? tmp25668 : tmp25625;
  assign tmp25671 = s1 ? tmp25601 : tmp25553;
  assign tmp25670 = s2 ? tmp25671 : tmp25553;
  assign tmp25669 = s3 ? tmp25670 : tmp25671;
  assign tmp25666 = s4 ? tmp25667 : tmp25669;
  assign tmp25659 = s5 ? tmp25660 : tmp25666;
  assign tmp25656 = s6 ? tmp25657 : tmp25659;
  assign tmp25627 = s7 ? tmp25628 : tmp25656;
  assign tmp25547 = s8 ? tmp25548 : tmp25627;
  assign tmp25679 = s0 ? tmp25553 : tmp24400;
  assign tmp25678 = s1 ? tmp25679 : tmp25553;
  assign tmp25677 = s2 ? tmp25557 : tmp25678;
  assign tmp25676 = s3 ? tmp25552 : tmp25677;
  assign tmp25675 = s4 ? tmp25676 : tmp25633;
  assign tmp25684 = s1 ? tmp25558 : tmp25679;
  assign tmp25683 = s2 ? tmp25572 : tmp25684;
  assign tmp25686 = s0 ? tmp24400 : tmp25553;
  assign tmp25685 = s2 ? tmp25686 : tmp25576;
  assign tmp25682 = s3 ? tmp25683 : tmp25685;
  assign tmp25681 = s4 ? tmp25682 : tmp25643;
  assign tmp25680 = s5 ? tmp25681 : tmp25587;
  assign tmp25674 = s6 ? tmp25675 : tmp25680;
  assign tmp25688 = s4 ? tmp25676 : tmp25658;
  assign tmp25693 = s1 ? tmp25553 : tmp25679;
  assign tmp25692 = s2 ? tmp25572 : tmp25693;
  assign tmp25691 = s3 ? tmp25692 : tmp25617;
  assign tmp25690 = s4 ? tmp25691 : tmp25664;
  assign tmp25694 = s4 ? tmp25667 : tmp25553;
  assign tmp25689 = s5 ? tmp25690 : tmp25694;
  assign tmp25687 = s6 ? tmp25688 : tmp25689;
  assign tmp25673 = s7 ? tmp25674 : tmp25687;
  assign tmp25672 = s8 ? tmp25627 : tmp25673;
  assign tmp25546 = s9 ? tmp25547 : tmp25672;
  assign tmp25701 = s3 ? tmp25553 : tmp25671;
  assign tmp25700 = s4 ? tmp25667 : tmp25701;
  assign tmp25699 = s5 ? tmp25690 : tmp25700;
  assign tmp25698 = s6 ? tmp25688 : tmp25699;
  assign tmp25697 = s7 ? tmp25674 : tmp25698;
  assign tmp25696 = s8 ? tmp25697 : tmp25674;
  assign tmp25706 = s4 ? tmp25623 : tmp25701;
  assign tmp25705 = s5 ? tmp25613 : tmp25706;
  assign tmp25704 = s6 ? tmp25608 : tmp25705;
  assign tmp25703 = s7 ? tmp25704 : tmp25687;
  assign tmp25707 = s7 ? tmp25656 : tmp25698;
  assign tmp25702 = s8 ? tmp25703 : tmp25707;
  assign tmp25695 = s9 ? tmp25696 : tmp25702;
  assign tmp25545 = s10 ? tmp25546 : tmp25695;
  assign tmp25711 = s7 ? tmp25607 : tmp25687;
  assign tmp25710 = s8 ? tmp25711 : tmp25707;
  assign tmp25709 = s9 ? tmp25696 : tmp25710;
  assign tmp25708 = s10 ? tmp25546 : tmp25709;
  assign tmp25544 = s11 ? tmp25545 : tmp25708;
  assign tmp25268 = s12 ? tmp25269 : tmp25544;
  assign tmp25719 = s0 ? tmp25071 : tmp25072;
  assign tmp25718 = s1 ? tmp25073 : tmp25719;
  assign tmp25722 = l1 ? tmp25072 : tmp25050;
  assign tmp25721 = s0 ? tmp25071 : tmp25722;
  assign tmp25723 = s1 ? tmp25071 : tmp25722;
  assign tmp25720 = s2 ? tmp25721 : tmp25723;
  assign tmp25717 = s3 ? tmp25718 : tmp25720;
  assign tmp25727 = s0 ? tmp25073 : tmp25071;
  assign tmp25726 = s1 ? tmp25727 : tmp25071;
  assign tmp25725 = s2 ? tmp25723 : tmp25726;
  assign tmp25729 = s1 ? tmp25071 : tmp25721;
  assign tmp25728 = s2 ? tmp25729 : tmp25722;
  assign tmp25724 = s3 ? tmp25725 : tmp25728;
  assign tmp25716 = s4 ? tmp25717 : tmp25724;
  assign tmp25735 = s0 ? tmp25072 : tmp25071;
  assign tmp25734 = s1 ? tmp25735 : tmp25071;
  assign tmp25737 = s0 ? tmp25722 : tmp25071;
  assign tmp25736 = s1 ? tmp25719 : tmp25737;
  assign tmp25733 = s2 ? tmp25734 : tmp25736;
  assign tmp25732 = s3 ? tmp25733 : tmp25728;
  assign tmp25741 = s0 ? tmp25073 : tmp25722;
  assign tmp25740 = s1 ? tmp25741 : tmp25071;
  assign tmp25739 = s2 ? tmp25740 : tmp25071;
  assign tmp25743 = s1 ? tmp25070 : tmp25721;
  assign tmp25745 = s0 ? tmp25722 : tmp25073;
  assign tmp25744 = s1 ? tmp25073 : tmp25745;
  assign tmp25742 = s2 ? tmp25743 : tmp25744;
  assign tmp25738 = s3 ? tmp25739 : tmp25742;
  assign tmp25731 = s4 ? tmp25732 : tmp25738;
  assign tmp25750 = s0 ? tmp25722 : tmp24943;
  assign tmp25751 = s0 ? tmp24943 : tmp25071;
  assign tmp25749 = s1 ? tmp25750 : tmp25751;
  assign tmp25748 = s2 ? tmp25749 : tmp25071;
  assign tmp25753 = s1 ? tmp25721 : tmp25722;
  assign tmp25754 = s1 ? tmp25745 : tmp25727;
  assign tmp25752 = s2 ? tmp25753 : tmp25754;
  assign tmp25747 = s3 ? tmp25748 : tmp25752;
  assign tmp25758 = s0 ? tmp25072 : tmp25722;
  assign tmp25757 = s1 ? tmp25719 : tmp25758;
  assign tmp25760 = s0 ? tmp24943 : tmp25072;
  assign tmp25759 = s1 ? tmp25760 : tmp25071;
  assign tmp25756 = s2 ? tmp25757 : tmp25759;
  assign tmp25763 = s0 ? tmp25722 : tmp25072;
  assign tmp25762 = s1 ? tmp25727 : tmp25763;
  assign tmp25761 = s2 ? tmp25753 : tmp25762;
  assign tmp25755 = s3 ? tmp25756 : tmp25761;
  assign tmp25746 = s4 ? tmp25747 : tmp25755;
  assign tmp25730 = s5 ? tmp25731 : tmp25746;
  assign tmp25715 = s6 ? tmp25716 : tmp25730;
  assign tmp25767 = s2 ? tmp25723 : tmp25722;
  assign tmp25766 = s3 ? tmp25725 : tmp25767;
  assign tmp25765 = s4 ? tmp25717 : tmp25766;
  assign tmp25772 = s1 ? tmp25072 : tmp25737;
  assign tmp25771 = s2 ? tmp25734 : tmp25772;
  assign tmp25770 = s3 ? tmp25771 : tmp25767;
  assign tmp25775 = s1 ? tmp25070 : tmp25722;
  assign tmp25776 = s1 ? tmp25073 : tmp25722;
  assign tmp25774 = s2 ? tmp25775 : tmp25776;
  assign tmp25773 = s3 ? tmp25739 : tmp25774;
  assign tmp25769 = s4 ? tmp25770 : tmp25773;
  assign tmp25780 = s1 ? tmp25750 : tmp25071;
  assign tmp25779 = s2 ? tmp25780 : tmp25071;
  assign tmp25782 = s1 ? tmp25073 : tmp25071;
  assign tmp25781 = s2 ? tmp25722 : tmp25782;
  assign tmp25778 = s3 ? tmp25779 : tmp25781;
  assign tmp25785 = s1 ? tmp25072 : tmp25722;
  assign tmp25784 = s2 ? tmp25785 : tmp25072;
  assign tmp25783 = s3 ? tmp25784 : tmp25722;
  assign tmp25777 = s4 ? tmp25778 : tmp25783;
  assign tmp25768 = s5 ? tmp25769 : tmp25777;
  assign tmp25764 = s6 ? tmp25765 : tmp25768;
  assign tmp25714 = s7 ? tmp25715 : tmp25764;
  assign tmp25787 = s8 ? tmp25714 : tmp25715;
  assign tmp25786 = s9 ? tmp25787 : tmp25764;
  assign tmp25713 = s10 ? tmp25714 : tmp25786;
  assign tmp25796 = l1 ? tmp25018 : tmp25072;
  assign tmp25797 = s0 ? tmp24514 : tmp25796;
  assign tmp25795 = s1 ? tmp25796 : tmp25797;
  assign tmp25801 = l1 ? tmp24401 : 1;
  assign tmp25800 = s0 ? tmp25801 : tmp25796;
  assign tmp25803 = l1 ? tmp25018 : 1;
  assign tmp25802 = s0 ? tmp25803 : tmp25796;
  assign tmp25799 = s1 ? tmp25800 : tmp25802;
  assign tmp25804 = s1 ? tmp25601 : tmp25796;
  assign tmp25798 = s2 ? tmp25799 : tmp25804;
  assign tmp25794 = s3 ? tmp25795 : tmp25798;
  assign tmp25808 = s0 ? tmp25337 : tmp24514;
  assign tmp25807 = s1 ? tmp25808 : tmp25796;
  assign tmp25811 = l1 ? tmp25554 : tmp25072;
  assign tmp25810 = s0 ? tmp25811 : tmp25337;
  assign tmp25809 = s1 ? tmp25810 : tmp24514;
  assign tmp25806 = s2 ? tmp25807 : tmp25809;
  assign tmp25815 = l1 ? tmp25050 : tmp25072;
  assign tmp25814 = s0 ? tmp25337 : tmp25815;
  assign tmp25813 = s1 ? tmp24514 : tmp25814;
  assign tmp25812 = s2 ? tmp25813 : tmp25796;
  assign tmp25805 = s3 ? tmp25806 : tmp25812;
  assign tmp25793 = s4 ? tmp25794 : tmp25805;
  assign tmp25821 = s0 ? tmp25796 : tmp24514;
  assign tmp25820 = s1 ? tmp25821 : tmp24514;
  assign tmp25823 = s0 ? tmp25796 : tmp25601;
  assign tmp25822 = s1 ? tmp25797 : tmp25823;
  assign tmp25819 = s2 ? tmp25820 : tmp25822;
  assign tmp25826 = s0 ? tmp25601 : tmp25803;
  assign tmp25827 = s0 ? tmp25601 : tmp25796;
  assign tmp25825 = s1 ? tmp25826 : tmp25827;
  assign tmp25829 = s0 ? tmp25796 : tmp25177;
  assign tmp25828 = s1 ? tmp25829 : tmp25796;
  assign tmp25824 = s2 ? tmp25825 : tmp25828;
  assign tmp25818 = s3 ? tmp25819 : tmp25824;
  assign tmp25833 = s0 ? tmp25815 : tmp25796;
  assign tmp25832 = s1 ? tmp25833 : tmp24514;
  assign tmp25834 = s1 ? tmp24514 : tmp25808;
  assign tmp25831 = s2 ? tmp25832 : tmp25834;
  assign tmp25838 = l1 ? tmp24401 : tmp25072;
  assign tmp25837 = s0 ? tmp25838 : tmp25796;
  assign tmp25836 = s1 ? tmp25837 : tmp25797;
  assign tmp25840 = s0 ? tmp25815 : tmp24870;
  assign tmp25839 = s1 ? tmp24870 : tmp25840;
  assign tmp25835 = s2 ? tmp25836 : tmp25839;
  assign tmp25830 = s3 ? tmp25831 : tmp25835;
  assign tmp25817 = s4 ? tmp25818 : tmp25830;
  assign tmp25845 = s0 ? tmp25177 : tmp25803;
  assign tmp25844 = s1 ? tmp25829 : tmp25845;
  assign tmp25847 = s0 ? tmp25601 : tmp24514;
  assign tmp25846 = s1 ? tmp25847 : tmp24514;
  assign tmp25843 = s2 ? tmp25844 : tmp25846;
  assign tmp25850 = s0 ? tmp24514 : tmp25072;
  assign tmp25851 = s0 ? tmp25072 : tmp25177;
  assign tmp25849 = s1 ? tmp25850 : tmp25851;
  assign tmp25853 = s0 ? tmp25177 : tmp25815;
  assign tmp25854 = s0 ? tmp25083 : tmp25337;
  assign tmp25852 = s1 ? tmp25853 : tmp25854;
  assign tmp25848 = s2 ? tmp25849 : tmp25852;
  assign tmp25842 = s3 ? tmp25843 : tmp25848;
  assign tmp25858 = s0 ? tmp25337 : tmp25796;
  assign tmp25857 = s1 ? tmp25858 : tmp25796;
  assign tmp25860 = s0 ? tmp25177 : tmp25796;
  assign tmp25859 = s1 ? tmp25860 : tmp24514;
  assign tmp25856 = s2 ? tmp25857 : tmp25859;
  assign tmp25862 = s1 ? tmp25802 : tmp25860;
  assign tmp25864 = s0 ? tmp25072 : tmp25796;
  assign tmp25863 = s1 ? tmp25854 : tmp25864;
  assign tmp25861 = s2 ? tmp25862 : tmp25863;
  assign tmp25855 = s3 ? tmp25856 : tmp25861;
  assign tmp25841 = s4 ? tmp25842 : tmp25855;
  assign tmp25816 = s5 ? tmp25817 : tmp25841;
  assign tmp25792 = s6 ? tmp25793 : tmp25816;
  assign tmp25869 = s1 ? tmp24514 : tmp25815;
  assign tmp25868 = s2 ? tmp25869 : tmp25796;
  assign tmp25867 = s3 ? tmp25806 : tmp25868;
  assign tmp25866 = s4 ? tmp25794 : tmp25867;
  assign tmp25874 = s1 ? tmp25796 : tmp25823;
  assign tmp25873 = s2 ? tmp25820 : tmp25874;
  assign tmp25876 = s1 ? tmp25803 : tmp25796;
  assign tmp25875 = s2 ? tmp25876 : tmp25828;
  assign tmp25872 = s3 ? tmp25873 : tmp25875;
  assign tmp25878 = s2 ? tmp25832 : tmp25337;
  assign tmp25880 = s1 ? tmp25837 : tmp25796;
  assign tmp25881 = s1 ? tmp24870 : tmp25815;
  assign tmp25879 = s2 ? tmp25880 : tmp25881;
  assign tmp25877 = s3 ? tmp25878 : tmp25879;
  assign tmp25871 = s4 ? tmp25872 : tmp25877;
  assign tmp25885 = s1 ? tmp25829 : tmp25601;
  assign tmp25884 = s2 ? tmp25885 : tmp24514;
  assign tmp25887 = s1 ? tmp25072 : tmp25177;
  assign tmp25888 = s1 ? tmp25083 : tmp25337;
  assign tmp25886 = s2 ? tmp25887 : tmp25888;
  assign tmp25883 = s3 ? tmp25884 : tmp25886;
  assign tmp25882 = s4 ? tmp25883 : tmp25796;
  assign tmp25870 = s5 ? tmp25871 : tmp25882;
  assign tmp25865 = s6 ? tmp25866 : tmp25870;
  assign tmp25791 = s7 ? tmp25792 : tmp25865;
  assign tmp25894 = s1 ? tmp25847 : tmp25796;
  assign tmp25893 = s2 ? tmp25799 : tmp25894;
  assign tmp25892 = s3 ? tmp25795 : tmp25893;
  assign tmp25891 = s4 ? tmp25892 : tmp25805;
  assign tmp25899 = s1 ? tmp25797 : tmp25821;
  assign tmp25898 = s2 ? tmp25820 : tmp25899;
  assign tmp25902 = s0 ? tmp24514 : tmp25803;
  assign tmp25901 = s1 ? tmp25902 : tmp25797;
  assign tmp25900 = s2 ? tmp25901 : tmp25828;
  assign tmp25897 = s3 ? tmp25898 : tmp25900;
  assign tmp25896 = s4 ? tmp25897 : tmp25830;
  assign tmp25895 = s5 ? tmp25896 : tmp25841;
  assign tmp25890 = s6 ? tmp25891 : tmp25895;
  assign tmp25904 = s4 ? tmp25892 : tmp25867;
  assign tmp25909 = s1 ? tmp25796 : tmp25821;
  assign tmp25908 = s2 ? tmp25820 : tmp25909;
  assign tmp25907 = s3 ? tmp25908 : tmp25875;
  assign tmp25906 = s4 ? tmp25907 : tmp25877;
  assign tmp25905 = s5 ? tmp25906 : tmp25882;
  assign tmp25903 = s6 ? tmp25904 : tmp25905;
  assign tmp25889 = s7 ? tmp25890 : tmp25903;
  assign tmp25790 = s8 ? tmp25791 : tmp25889;
  assign tmp25917 = s1 ? tmp25837 : tmp25858;
  assign tmp25916 = s2 ? tmp25917 : tmp25839;
  assign tmp25915 = s3 ? tmp25831 : tmp25916;
  assign tmp25914 = s4 ? tmp25897 : tmp25915;
  assign tmp25922 = s0 ? tmp25601 : tmp25801;
  assign tmp25921 = s1 ? tmp25922 : tmp25801;
  assign tmp25920 = s2 ? tmp25844 : tmp25921;
  assign tmp25919 = s3 ? tmp25920 : tmp25848;
  assign tmp25924 = s2 ? tmp25880 : tmp25859;
  assign tmp25927 = s0 ? tmp25083 : tmp25838;
  assign tmp25926 = s1 ? tmp25927 : tmp25864;
  assign tmp25925 = s2 ? tmp25862 : tmp25926;
  assign tmp25923 = s3 ? tmp25924 : tmp25925;
  assign tmp25918 = s4 ? tmp25919 : tmp25923;
  assign tmp25913 = s5 ? tmp25914 : tmp25918;
  assign tmp25912 = s6 ? tmp25891 : tmp25913;
  assign tmp25911 = s7 ? tmp25912 : tmp25903;
  assign tmp25910 = s8 ? tmp25889 : tmp25911;
  assign tmp25789 = s9 ? tmp25790 : tmp25910;
  assign tmp25936 = s0 ? tmp25811 : tmp25072;
  assign tmp25935 = s1 ? tmp25936 : tmp24514;
  assign tmp25934 = s2 ? tmp25807 : tmp25935;
  assign tmp25933 = s3 ? tmp25934 : tmp25812;
  assign tmp25932 = s4 ? tmp25892 : tmp25933;
  assign tmp25942 = s0 ? tmp25838 : tmp25811;
  assign tmp25941 = s1 ? tmp25942 : tmp25858;
  assign tmp25940 = s2 ? tmp25941 : tmp25839;
  assign tmp25939 = s3 ? tmp25831 : tmp25940;
  assign tmp25938 = s4 ? tmp25897 : tmp25939;
  assign tmp25937 = s5 ? tmp25938 : tmp25841;
  assign tmp25931 = s6 ? tmp25932 : tmp25937;
  assign tmp25945 = s3 ? tmp25934 : tmp25868;
  assign tmp25944 = s4 ? tmp25892 : tmp25945;
  assign tmp25943 = s6 ? tmp25944 : tmp25905;
  assign tmp25930 = s7 ? tmp25931 : tmp25943;
  assign tmp25929 = s8 ? tmp25930 : tmp25931;
  assign tmp25947 = s7 ? tmp25865 : tmp25903;
  assign tmp25948 = s7 ? tmp25903 : tmp25943;
  assign tmp25946 = s8 ? tmp25947 : tmp25948;
  assign tmp25928 = s9 ? tmp25929 : tmp25946;
  assign tmp25788 = s10 ? tmp25789 : tmp25928;
  assign tmp25712 = s12 ? tmp25713 : tmp25788;
  assign tmp25267 = s13 ? tmp25268 : tmp25712;
  assign tmp24858 = s14 ? tmp24859 : tmp25267;
  assign tmp23953 = s15 ? tmp23954 : tmp24858;
  assign tmp25964 = l1 ? tmp23984 : 1;
  assign tmp25963 = s0 ? tmp23987 : tmp25964;
  assign tmp25962 = s1 ? tmp25963 : tmp23982;
  assign tmp25961 = s2 ? tmp25962 : tmp24013;
  assign tmp25960 = s3 ? tmp25961 : tmp23982;
  assign tmp25968 = s0 ? tmp25964 : tmp23987;
  assign tmp25967 = s1 ? tmp25968 : tmp23987;
  assign tmp25966 = s2 ? tmp23982 : tmp25967;
  assign tmp25965 = s3 ? tmp25966 : tmp23982;
  assign tmp25959 = s4 ? tmp25960 : tmp25965;
  assign tmp25958 = s5 ? tmp23990 : tmp25959;
  assign tmp25957 = s6 ? tmp23961 : tmp25958;
  assign tmp25973 = s2 ? tmp25962 : tmp24007;
  assign tmp25972 = s3 ? tmp25973 : tmp23982;
  assign tmp25971 = s4 ? tmp25972 : tmp24035;
  assign tmp25970 = s5 ? tmp24025 : tmp25971;
  assign tmp25969 = s6 ? tmp24018 : tmp25970;
  assign tmp25956 = s7 ? tmp25957 : tmp25969;
  assign tmp25983 = l2 ? tmp23984 : 1;
  assign tmp25982 = l1 ? tmp25983 : tmp23966;
  assign tmp25981 = s0 ? tmp23987 : tmp25982;
  assign tmp25980 = s1 ? tmp23994 : tmp25981;
  assign tmp25979 = s2 ? tmp23993 : tmp25980;
  assign tmp25985 = s0 ? tmp25982 : tmp23987;
  assign tmp25984 = s2 ? tmp25985 : tmp24000;
  assign tmp25978 = s3 ? tmp25979 : tmp25984;
  assign tmp25977 = s4 ? tmp25978 : tmp24047;
  assign tmp25976 = s5 ? tmp25977 : tmp25959;
  assign tmp25975 = s6 ? tmp23961 : tmp25976;
  assign tmp25991 = s1 ? tmp23963 : tmp25981;
  assign tmp25990 = s2 ? tmp23970 : tmp25991;
  assign tmp25989 = s3 ? tmp25990 : tmp24029;
  assign tmp25996 = l2 ? tmp23984 : tmp23965;
  assign tmp25995 = l1 ? tmp25996 : tmp23966;
  assign tmp25997 = s0 ? tmp23963 : tmp25995;
  assign tmp25994 = s1 ? tmp25995 : tmp25997;
  assign tmp25993 = s2 ? tmp24004 : tmp25994;
  assign tmp25992 = s3 ? tmp25993 : tmp24048;
  assign tmp25988 = s4 ? tmp25989 : tmp25992;
  assign tmp25987 = s5 ? tmp25988 : tmp25971;
  assign tmp25986 = s6 ? tmp24018 : tmp25987;
  assign tmp25974 = s7 ? tmp25975 : tmp25986;
  assign tmp25955 = s8 ? tmp25956 : tmp25974;
  assign tmp26006 = l2 ? tmp23984 : tmp23974;
  assign tmp26005 = l1 ? tmp26006 : 1;
  assign tmp26004 = s0 ? tmp25995 : tmp26005;
  assign tmp26003 = s2 ? tmp25995 : tmp26004;
  assign tmp26009 = s0 ? tmp26005 : tmp23982;
  assign tmp26008 = s1 ? tmp25995 : tmp26009;
  assign tmp26012 = l1 ? tmp23984 : tmp23966;
  assign tmp26011 = s0 ? tmp25995 : tmp26012;
  assign tmp26013 = s0 ? tmp23982 : tmp25995;
  assign tmp26010 = s1 ? tmp26011 : tmp26013;
  assign tmp26007 = s2 ? tmp26008 : tmp26010;
  assign tmp26002 = s3 ? tmp26003 : tmp26007;
  assign tmp26001 = s4 ? tmp25995 : tmp26002;
  assign tmp26019 = s0 ? tmp25995 : tmp23963;
  assign tmp26018 = s1 ? tmp26019 : tmp25997;
  assign tmp26020 = s1 ? tmp25997 : tmp26012;
  assign tmp26017 = s2 ? tmp26018 : tmp26020;
  assign tmp26022 = s1 ? tmp26012 : tmp25985;
  assign tmp26024 = s0 ? tmp25995 : tmp25964;
  assign tmp26023 = s1 ? tmp23982 : tmp26024;
  assign tmp26021 = s2 ? tmp26022 : tmp26023;
  assign tmp26016 = s3 ? tmp26017 : tmp26021;
  assign tmp26027 = s1 ? tmp26013 : tmp26024;
  assign tmp26028 = s1 ? tmp26024 : tmp25995;
  assign tmp26026 = s2 ? tmp26027 : tmp26028;
  assign tmp26031 = s0 ? tmp25964 : tmp23982;
  assign tmp26030 = s1 ? tmp25963 : tmp26031;
  assign tmp26029 = s2 ? tmp26030 : tmp23982;
  assign tmp26025 = s3 ? tmp26026 : tmp26029;
  assign tmp26015 = s4 ? tmp26016 : tmp26025;
  assign tmp26014 = s5 ? tmp26015 : tmp24008;
  assign tmp26000 = s6 ? tmp26001 : tmp26014;
  assign tmp26036 = s1 ? tmp26004 : tmp25995;
  assign tmp26035 = s2 ? tmp25995 : tmp26036;
  assign tmp26038 = s1 ? tmp25995 : tmp23982;
  assign tmp26037 = s2 ? tmp26038 : tmp26010;
  assign tmp26034 = s3 ? tmp26035 : tmp26037;
  assign tmp26033 = s4 ? tmp25995 : tmp26034;
  assign tmp26043 = s1 ? tmp26019 : tmp25995;
  assign tmp26044 = s1 ? tmp25995 : tmp26012;
  assign tmp26042 = s2 ? tmp26043 : tmp26044;
  assign tmp26046 = s1 ? tmp26012 : tmp23987;
  assign tmp26045 = s2 ? tmp26046 : tmp26023;
  assign tmp26041 = s3 ? tmp26042 : tmp26045;
  assign tmp26048 = s2 ? tmp26027 : tmp25995;
  assign tmp26049 = s2 ? tmp25962 : tmp23982;
  assign tmp26047 = s3 ? tmp26048 : tmp26049;
  assign tmp26040 = s4 ? tmp26041 : tmp26047;
  assign tmp26039 = s5 ? tmp26040 : tmp24032;
  assign tmp26032 = s6 ? tmp26033 : tmp26039;
  assign tmp25999 = s7 ? tmp26000 : tmp26032;
  assign tmp25998 = s8 ? tmp25974 : tmp25999;
  assign tmp25954 = s9 ? tmp25955 : tmp25998;
  assign tmp26059 = l1 ? tmp26006 : tmp23966;
  assign tmp26058 = s0 ? tmp25995 : tmp26059;
  assign tmp26057 = s1 ? tmp26058 : tmp25995;
  assign tmp26056 = s2 ? tmp25995 : tmp26057;
  assign tmp26055 = s3 ? tmp25995 : tmp26056;
  assign tmp26054 = s4 ? tmp26055 : tmp26002;
  assign tmp26065 = s0 ? tmp25995 : tmp23972;
  assign tmp26066 = s0 ? tmp23972 : tmp25995;
  assign tmp26064 = s1 ? tmp26065 : tmp26066;
  assign tmp26068 = s0 ? tmp26012 : tmp25982;
  assign tmp26067 = s1 ? tmp26066 : tmp26068;
  assign tmp26063 = s2 ? tmp26064 : tmp26067;
  assign tmp26071 = s0 ? tmp25982 : tmp26012;
  assign tmp26070 = s1 ? tmp26071 : tmp25985;
  assign tmp26069 = s2 ? tmp26070 : tmp26023;
  assign tmp26062 = s3 ? tmp26063 : tmp26069;
  assign tmp26061 = s4 ? tmp26062 : tmp26025;
  assign tmp26060 = s5 ? tmp26061 : tmp25959;
  assign tmp26053 = s6 ? tmp26054 : tmp26060;
  assign tmp26073 = s4 ? tmp26055 : tmp26034;
  assign tmp26078 = s1 ? tmp26065 : tmp25995;
  assign tmp26079 = s1 ? tmp25995 : tmp26068;
  assign tmp26077 = s2 ? tmp26078 : tmp26079;
  assign tmp26076 = s3 ? tmp26077 : tmp26045;
  assign tmp26075 = s4 ? tmp26076 : tmp26047;
  assign tmp26074 = s5 ? tmp26075 : tmp25971;
  assign tmp26072 = s6 ? tmp26073 : tmp26074;
  assign tmp26052 = s7 ? tmp26053 : tmp26072;
  assign tmp26051 = s8 ? tmp26052 : tmp26053;
  assign tmp26081 = s7 ? tmp25969 : tmp26032;
  assign tmp26088 = s1 ? tmp25995 : tmp23963;
  assign tmp26087 = s2 ? tmp24004 : tmp26088;
  assign tmp26086 = s3 ? tmp26087 : tmp24048;
  assign tmp26085 = s4 ? tmp25989 : tmp26086;
  assign tmp26084 = s5 ? tmp26085 : tmp25971;
  assign tmp26083 = s6 ? tmp24018 : tmp26084;
  assign tmp26082 = s7 ? tmp26083 : tmp26072;
  assign tmp26080 = s8 ? tmp26081 : tmp26082;
  assign tmp26050 = s9 ? tmp26051 : tmp26080;
  assign tmp25953 = s10 ? tmp25954 : tmp26050;
  assign tmp26092 = s7 ? tmp25986 : tmp26072;
  assign tmp26091 = s8 ? tmp26081 : tmp26092;
  assign tmp26090 = s9 ? tmp26051 : tmp26091;
  assign tmp26089 = s10 ? tmp25954 : tmp26090;
  assign tmp25952 = s11 ? tmp25953 : tmp26089;
  assign tmp26105 = l1 ? tmp25983 : 1;
  assign tmp26104 = s0 ? tmp23973 : tmp26105;
  assign tmp26103 = s1 ? tmp23973 : tmp26104;
  assign tmp26107 = s0 ? tmp26105 : tmp23973;
  assign tmp26106 = s1 ? tmp24209 : tmp26107;
  assign tmp26102 = s2 ? tmp26103 : tmp26106;
  assign tmp26101 = s3 ? tmp23973 : tmp26102;
  assign tmp26100 = s4 ? tmp23973 : tmp26101;
  assign tmp26113 = s0 ? tmp24210 : tmp26105;
  assign tmp26112 = s1 ? tmp24210 : tmp26113;
  assign tmp26115 = s0 ? tmp23978 : tmp26105;
  assign tmp26114 = s1 ? tmp26105 : tmp26115;
  assign tmp26111 = s2 ? tmp26112 : tmp26114;
  assign tmp26110 = s3 ? tmp24215 : tmp26111;
  assign tmp26119 = s0 ? tmp26105 : tmp23978;
  assign tmp26118 = s1 ? tmp26119 : tmp26115;
  assign tmp26120 = s1 ? tmp26115 : tmp23978;
  assign tmp26117 = s2 ? tmp26118 : tmp26120;
  assign tmp26116 = s3 ? tmp26117 : tmp26105;
  assign tmp26109 = s4 ? tmp26110 : tmp26116;
  assign tmp26108 = s5 ? tmp26109 : tmp26105;
  assign tmp26099 = s6 ? tmp26100 : tmp26108;
  assign tmp26126 = s1 ? tmp24210 : tmp26105;
  assign tmp26125 = s2 ? tmp26126 : tmp26114;
  assign tmp26124 = s3 ? tmp24254 : tmp26125;
  assign tmp26128 = s2 ? tmp26118 : tmp23978;
  assign tmp26127 = s3 ? tmp26128 : tmp26105;
  assign tmp26123 = s4 ? tmp26124 : tmp26127;
  assign tmp26122 = s5 ? tmp26123 : tmp26105;
  assign tmp26121 = s6 ? tmp26100 : tmp26122;
  assign tmp26098 = s7 ? tmp26099 : tmp26121;
  assign tmp26134 = s1 ? tmp23973 : tmp26107;
  assign tmp26133 = s2 ? tmp26103 : tmp26134;
  assign tmp26132 = s3 ? tmp23973 : tmp26133;
  assign tmp26131 = s4 ? tmp23973 : tmp26132;
  assign tmp26139 = s1 ? tmp26105 : tmp23978;
  assign tmp26138 = s2 ? tmp26103 : tmp26139;
  assign tmp26137 = s3 ? tmp24280 : tmp26138;
  assign tmp26142 = s1 ? tmp26119 : tmp23978;
  assign tmp26141 = s2 ? tmp26142 : tmp23978;
  assign tmp26140 = s3 ? tmp26141 : tmp26105;
  assign tmp26136 = s4 ? tmp26137 : tmp26140;
  assign tmp26135 = s5 ? tmp26136 : tmp26105;
  assign tmp26130 = s6 ? tmp26131 : tmp26135;
  assign tmp26149 = l1 ? tmp26006 : tmp23973;
  assign tmp26148 = s0 ? tmp23973 : tmp26149;
  assign tmp26147 = s1 ? tmp23973 : tmp26148;
  assign tmp26146 = s2 ? tmp23973 : tmp26147;
  assign tmp26152 = s0 ? tmp26149 : tmp26105;
  assign tmp26151 = s1 ? tmp23973 : tmp26152;
  assign tmp26150 = s2 ? tmp26151 : tmp26134;
  assign tmp26145 = s3 ? tmp26146 : tmp26150;
  assign tmp26144 = s4 ? tmp23973 : tmp26145;
  assign tmp26157 = s1 ? tmp23973 : tmp26105;
  assign tmp26156 = s2 ? tmp26157 : tmp26139;
  assign tmp26155 = s3 ? tmp24304 : tmp26156;
  assign tmp26154 = s4 ? tmp26155 : tmp26140;
  assign tmp26153 = s5 ? tmp26154 : tmp26105;
  assign tmp26143 = s6 ? tmp26144 : tmp26153;
  assign tmp26129 = s7 ? tmp26130 : tmp26143;
  assign tmp26097 = s8 ? tmp26098 : tmp26129;
  assign tmp26164 = s1 ? tmp26149 : tmp26152;
  assign tmp26166 = s0 ? tmp26105 : tmp26149;
  assign tmp26165 = s1 ? tmp26149 : tmp26166;
  assign tmp26163 = s2 ? tmp26164 : tmp26165;
  assign tmp26162 = s3 ? tmp26149 : tmp26163;
  assign tmp26161 = s4 ? tmp26149 : tmp26162;
  assign tmp26172 = s0 ? tmp26149 : tmp23973;
  assign tmp26171 = s1 ? tmp26172 : tmp26148;
  assign tmp26174 = s0 ? tmp23973 : tmp26005;
  assign tmp26175 = l1 ? tmp25983 : tmp23973;
  assign tmp26173 = s1 ? tmp26174 : tmp26175;
  assign tmp26170 = s2 ? tmp26171 : tmp26173;
  assign tmp26178 = s0 ? tmp26175 : tmp26105;
  assign tmp26177 = s1 ? tmp26175 : tmp26178;
  assign tmp26179 = s1 ? tmp26105 : tmp26005;
  assign tmp26176 = s2 ? tmp26177 : tmp26179;
  assign tmp26169 = s3 ? tmp26170 : tmp26176;
  assign tmp26183 = s0 ? tmp26105 : tmp26005;
  assign tmp26182 = s1 ? tmp26183 : tmp26005;
  assign tmp26181 = s2 ? tmp26182 : tmp26005;
  assign tmp26180 = s3 ? tmp26181 : tmp26105;
  assign tmp26168 = s4 ? tmp26169 : tmp26180;
  assign tmp26167 = s5 ? tmp26168 : tmp26105;
  assign tmp26160 = s6 ? tmp26161 : tmp26167;
  assign tmp26189 = s1 ? tmp26172 : tmp26149;
  assign tmp26190 = s1 ? tmp26005 : tmp26175;
  assign tmp26188 = s2 ? tmp26189 : tmp26190;
  assign tmp26192 = s1 ? tmp26175 : tmp26105;
  assign tmp26191 = s2 ? tmp26192 : tmp26179;
  assign tmp26187 = s3 ? tmp26188 : tmp26191;
  assign tmp26186 = s4 ? tmp26187 : tmp26180;
  assign tmp26185 = s5 ? tmp26186 : tmp26105;
  assign tmp26184 = s6 ? tmp26161 : tmp26185;
  assign tmp26159 = s7 ? tmp26160 : tmp26184;
  assign tmp26158 = s8 ? tmp26129 : tmp26159;
  assign tmp26096 = s9 ? tmp26097 : tmp26158;
  assign tmp26194 = s8 ? tmp26159 : tmp26160;
  assign tmp26200 = s2 ? tmp26157 : tmp26106;
  assign tmp26199 = s3 ? tmp23973 : tmp26200;
  assign tmp26198 = s4 ? tmp23973 : tmp26199;
  assign tmp26197 = s6 ? tmp26198 : tmp26122;
  assign tmp26205 = s1 ? tmp26149 : tmp26105;
  assign tmp26204 = s2 ? tmp26205 : tmp26165;
  assign tmp26203 = s3 ? tmp26149 : tmp26204;
  assign tmp26202 = s4 ? tmp26149 : tmp26203;
  assign tmp26201 = s6 ? tmp26202 : tmp26185;
  assign tmp26196 = s7 ? tmp26197 : tmp26201;
  assign tmp26210 = s2 ? tmp26157 : tmp26134;
  assign tmp26209 = s3 ? tmp26146 : tmp26210;
  assign tmp26208 = s4 ? tmp23973 : tmp26209;
  assign tmp26207 = s6 ? tmp26208 : tmp26153;
  assign tmp26206 = s7 ? tmp26207 : tmp26201;
  assign tmp26195 = s8 ? tmp26196 : tmp26206;
  assign tmp26193 = s9 ? tmp26194 : tmp26195;
  assign tmp26095 = s10 ? tmp26096 : tmp26193;
  assign tmp26214 = s7 ? tmp26121 : tmp26184;
  assign tmp26215 = s7 ? tmp26143 : tmp26184;
  assign tmp26213 = s8 ? tmp26214 : tmp26215;
  assign tmp26212 = s9 ? tmp26194 : tmp26213;
  assign tmp26211 = s10 ? tmp26096 : tmp26212;
  assign tmp26094 = s11 ? tmp26095 : tmp26211;
  assign tmp26093 = s12 ? tmp24077 : tmp26094;
  assign tmp25951 = s13 ? tmp25952 : tmp26093;
  assign tmp26225 = l1 ? tmp25983 : tmp23974;
  assign tmp26228 = s0 ? tmp26225 : tmp26175;
  assign tmp26227 = s2 ? tmp26225 : tmp26228;
  assign tmp26231 = s0 ? tmp26175 : tmp23997;
  assign tmp26230 = s1 ? tmp26225 : tmp26231;
  assign tmp26233 = s0 ? tmp23997 : tmp26225;
  assign tmp26232 = s1 ? tmp26225 : tmp26233;
  assign tmp26229 = s2 ? tmp26230 : tmp26232;
  assign tmp26226 = s3 ? tmp26227 : tmp26229;
  assign tmp26224 = s4 ? tmp26225 : tmp26226;
  assign tmp26239 = s0 ? tmp26225 : tmp24093;
  assign tmp26240 = s0 ? tmp24093 : tmp26225;
  assign tmp26238 = s1 ? tmp26239 : tmp26240;
  assign tmp26242 = s0 ? tmp24093 : tmp25982;
  assign tmp26241 = s1 ? tmp26242 : tmp26225;
  assign tmp26237 = s2 ? tmp26238 : tmp26241;
  assign tmp26245 = s0 ? tmp26225 : tmp23997;
  assign tmp26244 = s1 ? tmp26225 : tmp26245;
  assign tmp26248 = l1 ? 1 : tmp25983;
  assign tmp26247 = s0 ? tmp23997 : tmp26248;
  assign tmp26249 = s0 ? tmp25982 : tmp25983;
  assign tmp26246 = s1 ? tmp26247 : tmp26249;
  assign tmp26243 = s2 ? tmp26244 : tmp26246;
  assign tmp26236 = s3 ? tmp26237 : tmp26243;
  assign tmp26253 = s0 ? tmp23997 : tmp25982;
  assign tmp26252 = s1 ? tmp26253 : tmp26249;
  assign tmp26254 = s1 ? tmp26249 : tmp25982;
  assign tmp26251 = s2 ? tmp26252 : tmp26254;
  assign tmp26257 = s0 ? tmp23997 : tmp25983;
  assign tmp26258 = s0 ? tmp25983 : tmp26248;
  assign tmp26256 = s1 ? tmp26257 : tmp26258;
  assign tmp26259 = s1 ? tmp26247 : tmp26248;
  assign tmp26255 = s2 ? tmp26256 : tmp26259;
  assign tmp26250 = s3 ? tmp26251 : tmp26255;
  assign tmp26235 = s4 ? tmp26236 : tmp26250;
  assign tmp26234 = s5 ? tmp26235 : tmp23997;
  assign tmp26223 = s6 ? tmp26224 : tmp26234;
  assign tmp26264 = s1 ? tmp26228 : tmp25982;
  assign tmp26263 = s2 ? tmp26225 : tmp26264;
  assign tmp26266 = s1 ? tmp26225 : tmp23997;
  assign tmp26265 = s2 ? tmp26266 : tmp26232;
  assign tmp26262 = s3 ? tmp26263 : tmp26265;
  assign tmp26261 = s4 ? tmp26225 : tmp26262;
  assign tmp26271 = s1 ? tmp26239 : tmp26225;
  assign tmp26272 = s1 ? tmp25982 : tmp26225;
  assign tmp26270 = s2 ? tmp26271 : tmp26272;
  assign tmp26276 = ~(l2 ? tmp23968 : tmp23967);
  assign tmp26275 = l1 ? tmp25983 : tmp26276;
  assign tmp26277 = s0 ? tmp26275 : tmp23997;
  assign tmp26274 = s1 ? tmp26275 : tmp26277;
  assign tmp26273 = s2 ? tmp26274 : tmp26246;
  assign tmp26269 = s3 ? tmp26270 : tmp26273;
  assign tmp26279 = s2 ? tmp26252 : tmp25982;
  assign tmp26281 = s1 ? tmp26257 : tmp26248;
  assign tmp26280 = s2 ? tmp26281 : tmp23997;
  assign tmp26278 = s3 ? tmp26279 : tmp26280;
  assign tmp26268 = s4 ? tmp26269 : tmp26278;
  assign tmp26267 = s5 ? tmp26268 : tmp23997;
  assign tmp26260 = s6 ? tmp26261 : tmp26267;
  assign tmp26222 = s7 ? tmp26223 : tmp26260;
  assign tmp26221 = s8 ? tmp24347 : tmp26222;
  assign tmp26220 = s9 ? tmp26221 : tmp26222;
  assign tmp26283 = s8 ? tmp26222 : tmp26223;
  assign tmp26291 = s1 ? tmp26275 : tmp23997;
  assign tmp26290 = s2 ? tmp26291 : tmp26246;
  assign tmp26289 = s3 ? tmp26270 : tmp26290;
  assign tmp26288 = s4 ? tmp26289 : tmp26278;
  assign tmp26287 = s5 ? tmp26288 : tmp23997;
  assign tmp26286 = s6 ? tmp26261 : tmp26287;
  assign tmp26285 = s7 ? tmp24385 : tmp26286;
  assign tmp26284 = s8 ? tmp26285 : tmp26286;
  assign tmp26282 = s9 ? tmp26283 : tmp26284;
  assign tmp26219 = s10 ? tmp26220 : tmp26282;
  assign tmp26295 = s7 ? tmp24362 : tmp26260;
  assign tmp26294 = s8 ? tmp26295 : tmp26260;
  assign tmp26293 = s9 ? tmp26283 : tmp26294;
  assign tmp26292 = s10 ? tmp26220 : tmp26293;
  assign tmp26218 = s11 ? tmp26219 : tmp26292;
  assign tmp26306 = s0 ? tmp24399 : tmp26105;
  assign tmp26305 = s1 ? tmp26306 : tmp24399;
  assign tmp26304 = s2 ? tmp24399 : tmp26305;
  assign tmp26303 = s3 ? tmp24399 : tmp26304;
  assign tmp26308 = s2 ? tmp24403 : tmp26306;
  assign tmp26311 = s0 ? tmp26105 : tmp24410;
  assign tmp26310 = s1 ? tmp24399 : tmp26311;
  assign tmp26309 = s2 ? tmp26310 : tmp24411;
  assign tmp26307 = s3 ? tmp26308 : tmp26309;
  assign tmp26302 = s4 ? tmp26303 : tmp26307;
  assign tmp26317 = s0 ? tmp26105 : tmp23982;
  assign tmp26316 = s1 ? tmp26306 : tmp26317;
  assign tmp26319 = s0 ? tmp26105 : tmp24399;
  assign tmp26318 = s1 ? tmp26319 : tmp26306;
  assign tmp26315 = s2 ? tmp26316 : tmp26318;
  assign tmp26320 = s2 ? tmp26319 : tmp24421;
  assign tmp26314 = s3 ? tmp26315 : tmp26320;
  assign tmp26313 = s4 ? tmp26314 : tmp24422;
  assign tmp26312 = s5 ? tmp26313 : tmp24427;
  assign tmp26301 = s6 ? tmp26302 : tmp26312;
  assign tmp26324 = s2 ? tmp24403 : tmp26305;
  assign tmp26323 = s3 ? tmp26324 : tmp24445;
  assign tmp26322 = s4 ? tmp26303 : tmp26323;
  assign tmp26329 = s1 ? tmp26306 : tmp23982;
  assign tmp26330 = s1 ? tmp24399 : tmp26306;
  assign tmp26328 = s2 ? tmp26329 : tmp26330;
  assign tmp26327 = s3 ? tmp26328 : tmp24420;
  assign tmp26326 = s4 ? tmp26327 : tmp24451;
  assign tmp26325 = s5 ? tmp26326 : tmp24453;
  assign tmp26321 = s6 ? tmp26322 : tmp26325;
  assign tmp26300 = s7 ? tmp26301 : tmp26321;
  assign tmp26336 = l2 ? tmp25280 : 1;
  assign tmp26335 = l1 ? tmp23984 : tmp26336;
  assign tmp26339 = s0 ? tmp26335 : tmp25983;
  assign tmp26338 = s1 ? tmp26339 : tmp26335;
  assign tmp26337 = s2 ? tmp26335 : tmp26338;
  assign tmp26334 = s3 ? tmp26335 : tmp26337;
  assign tmp26343 = s0 ? tmp26335 : tmp25964;
  assign tmp26342 = s1 ? tmp26343 : tmp26335;
  assign tmp26344 = s0 ? tmp26335 : tmp26105;
  assign tmp26341 = s2 ? tmp26342 : tmp26344;
  assign tmp26346 = s1 ? tmp26335 : tmp26311;
  assign tmp26349 = l1 ? 1 : tmp26336;
  assign tmp26348 = s0 ? tmp26349 : tmp26335;
  assign tmp26347 = s1 ? tmp26335 : tmp26348;
  assign tmp26345 = s2 ? tmp26346 : tmp26347;
  assign tmp26340 = s3 ? tmp26341 : tmp26345;
  assign tmp26333 = s4 ? tmp26334 : tmp26340;
  assign tmp26356 = l1 ? tmp23984 : tmp25983;
  assign tmp26355 = s0 ? tmp26105 : tmp26356;
  assign tmp26354 = s1 ? tmp26344 : tmp26355;
  assign tmp26358 = s0 ? tmp26105 : tmp26335;
  assign tmp26357 = s1 ? tmp26358 : tmp26339;
  assign tmp26353 = s2 ? tmp26354 : tmp26357;
  assign tmp26361 = s0 ? tmp25983 : tmp26335;
  assign tmp26363 = l1 ? tmp23983 : tmp26336;
  assign tmp26362 = s0 ? tmp25983 : tmp26363;
  assign tmp26360 = s1 ? tmp26361 : tmp26362;
  assign tmp26365 = s0 ? tmp26349 : tmp24410;
  assign tmp26364 = s1 ? tmp26365 : tmp26335;
  assign tmp26359 = s2 ? tmp26360 : tmp26364;
  assign tmp26352 = s3 ? tmp26353 : tmp26359;
  assign tmp26369 = s0 ? tmp24410 : tmp26335;
  assign tmp26370 = s0 ? tmp26356 : tmp26335;
  assign tmp26368 = s1 ? tmp26369 : tmp26370;
  assign tmp26371 = s1 ? tmp26370 : tmp26343;
  assign tmp26367 = s2 ? tmp26368 : tmp26371;
  assign tmp26374 = s0 ? tmp26363 : tmp26335;
  assign tmp26375 = s0 ? tmp26335 : tmp24399;
  assign tmp26373 = s1 ? tmp26374 : tmp26375;
  assign tmp26372 = s2 ? tmp26373 : tmp24410;
  assign tmp26366 = s3 ? tmp26367 : tmp26372;
  assign tmp26351 = s4 ? tmp26352 : tmp26366;
  assign tmp26380 = s0 ? tmp26363 : tmp24410;
  assign tmp26381 = s0 ? tmp24410 : tmp26349;
  assign tmp26379 = s1 ? tmp26380 : tmp26381;
  assign tmp26384 = l1 ? tmp23983 : tmp25983;
  assign tmp26383 = s0 ? tmp26349 : tmp26384;
  assign tmp26382 = s1 ? tmp26383 : tmp26384;
  assign tmp26378 = s2 ? tmp26379 : tmp26382;
  assign tmp26377 = s3 ? tmp26378 : tmp24434;
  assign tmp26387 = s1 ? tmp24431 : tmp26381;
  assign tmp26389 = s0 ? tmp24410 : tmp26363;
  assign tmp26388 = s1 ? tmp26389 : tmp26384;
  assign tmp26386 = s2 ? tmp26387 : tmp26388;
  assign tmp26391 = s1 ? tmp26365 : tmp24412;
  assign tmp26390 = s2 ? tmp26391 : tmp24441;
  assign tmp26385 = s3 ? tmp26386 : tmp26390;
  assign tmp26376 = s4 ? tmp26377 : tmp26385;
  assign tmp26350 = s5 ? tmp26351 : tmp26376;
  assign tmp26332 = s6 ? tmp26333 : tmp26350;
  assign tmp26396 = s1 ? tmp26344 : tmp26335;
  assign tmp26395 = s2 ? tmp26342 : tmp26396;
  assign tmp26398 = s1 ? tmp26335 : tmp24410;
  assign tmp26397 = s2 ? tmp26398 : tmp26347;
  assign tmp26394 = s3 ? tmp26395 : tmp26397;
  assign tmp26393 = s4 ? tmp26334 : tmp26394;
  assign tmp26403 = s1 ? tmp26344 : tmp26356;
  assign tmp26404 = s1 ? tmp26335 : tmp26339;
  assign tmp26402 = s2 ? tmp26403 : tmp26404;
  assign tmp26406 = s1 ? tmp26335 : tmp26363;
  assign tmp26405 = s2 ? tmp26406 : tmp26364;
  assign tmp26401 = s3 ? tmp26402 : tmp26405;
  assign tmp26408 = s2 ? tmp26368 : tmp26335;
  assign tmp26407 = s3 ? tmp26408 : tmp26372;
  assign tmp26400 = s4 ? tmp26401 : tmp26407;
  assign tmp26412 = s1 ? tmp26380 : tmp26349;
  assign tmp26413 = s1 ? tmp26384 : tmp23982;
  assign tmp26411 = s2 ? tmp26412 : tmp26413;
  assign tmp26410 = s3 ? tmp26411 : tmp24456;
  assign tmp26416 = s1 ? tmp24410 : tmp26349;
  assign tmp26415 = s2 ? tmp26416 : tmp26363;
  assign tmp26414 = s3 ? tmp26415 : tmp24421;
  assign tmp26409 = s4 ? tmp26410 : tmp26414;
  assign tmp26399 = s5 ? tmp26400 : tmp26409;
  assign tmp26392 = s6 ? tmp26393 : tmp26399;
  assign tmp26331 = s7 ? tmp26332 : tmp26392;
  assign tmp26299 = s8 ? tmp26300 : tmp26331;
  assign tmp26424 = s0 ? tmp26335 : tmp26356;
  assign tmp26423 = s1 ? tmp26424 : tmp26335;
  assign tmp26422 = s2 ? tmp26423 : tmp26344;
  assign tmp26421 = s3 ? tmp26422 : tmp26345;
  assign tmp26420 = s4 ? tmp26335 : tmp26421;
  assign tmp26429 = s1 ? tmp26358 : tmp26335;
  assign tmp26428 = s2 ? tmp26354 : tmp26429;
  assign tmp26433 = l1 ? tmp25983 : tmp26336;
  assign tmp26432 = s0 ? tmp26433 : tmp26363;
  assign tmp26431 = s1 ? tmp26335 : tmp26432;
  assign tmp26430 = s2 ? tmp26431 : tmp26364;
  assign tmp26427 = s3 ? tmp26428 : tmp26430;
  assign tmp26436 = s1 ? tmp26370 : tmp26424;
  assign tmp26435 = s2 ? tmp26368 : tmp26436;
  assign tmp26434 = s3 ? tmp26435 : tmp26372;
  assign tmp26426 = s4 ? tmp26427 : tmp26434;
  assign tmp26425 = s5 ? tmp26426 : tmp26376;
  assign tmp26419 = s6 ? tmp26420 : tmp26425;
  assign tmp26440 = s2 ? tmp26423 : tmp26396;
  assign tmp26439 = s3 ? tmp26440 : tmp26397;
  assign tmp26438 = s4 ? tmp26335 : tmp26439;
  assign tmp26444 = s2 ? tmp26403 : tmp26335;
  assign tmp26443 = s3 ? tmp26444 : tmp26405;
  assign tmp26442 = s4 ? tmp26443 : tmp26407;
  assign tmp26441 = s5 ? tmp26442 : tmp26409;
  assign tmp26437 = s6 ? tmp26438 : tmp26441;
  assign tmp26418 = s7 ? tmp26419 : tmp26437;
  assign tmp26417 = s8 ? tmp26331 : tmp26418;
  assign tmp26298 = s9 ? tmp26299 : tmp26417;
  assign tmp26446 = s8 ? tmp26331 : tmp26332;
  assign tmp26454 = s1 ? tmp26374 : tmp24399;
  assign tmp26453 = s2 ? tmp26454 : tmp24410;
  assign tmp26452 = s3 ? tmp26408 : tmp26453;
  assign tmp26451 = s4 ? tmp26443 : tmp26452;
  assign tmp26450 = s5 ? tmp26451 : tmp26409;
  assign tmp26449 = s6 ? tmp26438 : tmp26450;
  assign tmp26448 = s7 ? tmp26321 : tmp26449;
  assign tmp26457 = s4 ? tmp26401 : tmp26452;
  assign tmp26456 = s5 ? tmp26457 : tmp26409;
  assign tmp26455 = s6 ? tmp26393 : tmp26456;
  assign tmp26447 = s8 ? tmp26448 : tmp26455;
  assign tmp26445 = s9 ? tmp26446 : tmp26447;
  assign tmp26297 = s10 ? tmp26298 : tmp26445;
  assign tmp26461 = s7 ? tmp26321 : tmp26437;
  assign tmp26460 = s8 ? tmp26461 : tmp26392;
  assign tmp26459 = s9 ? tmp26446 : tmp26460;
  assign tmp26458 = s10 ? tmp26298 : tmp26459;
  assign tmp26296 = s11 ? tmp26297 : tmp26458;
  assign tmp26217 = s12 ? tmp26218 : tmp26296;
  assign tmp26473 = ~(l2 ? tmp23968 : 0);
  assign tmp26472 = l1 ? tmp24499 : tmp26473;
  assign tmp26475 = l1 ? tmp23983 : tmp26473;
  assign tmp26474 = s0 ? tmp26475 : tmp26472;
  assign tmp26471 = s1 ? tmp26472 : tmp26474;
  assign tmp26479 = l1 ? 1 : tmp26473;
  assign tmp26478 = s0 ? tmp26472 : tmp26479;
  assign tmp26477 = s1 ? tmp26478 : tmp26472;
  assign tmp26476 = s2 ? tmp26472 : tmp26477;
  assign tmp26470 = s3 ? tmp26471 : tmp26476;
  assign tmp26483 = s0 ? tmp26472 : tmp26475;
  assign tmp26482 = s1 ? tmp26483 : tmp26472;
  assign tmp26485 = s0 ? tmp26472 : tmp23997;
  assign tmp26486 = s0 ? tmp26475 : tmp23997;
  assign tmp26484 = s1 ? tmp26485 : tmp26486;
  assign tmp26481 = s2 ? tmp26482 : tmp26484;
  assign tmp26488 = s1 ? tmp26475 : tmp24513;
  assign tmp26490 = s0 ? tmp24514 : tmp26472;
  assign tmp26489 = s1 ? tmp26472 : tmp26490;
  assign tmp26487 = s2 ? tmp26488 : tmp26489;
  assign tmp26480 = s3 ? tmp26481 : tmp26487;
  assign tmp26469 = s4 ? tmp26470 : tmp26480;
  assign tmp26496 = s0 ? tmp26479 : tmp26472;
  assign tmp26495 = s1 ? tmp26478 : tmp26496;
  assign tmp26497 = s1 ? tmp26496 : tmp26478;
  assign tmp26494 = s2 ? tmp26495 : tmp26497;
  assign tmp26501 = l1 ? tmp24499 : tmp25983;
  assign tmp26500 = s0 ? tmp26472 : tmp26501;
  assign tmp26499 = s1 ? tmp24514 : tmp26500;
  assign tmp26498 = s2 ? tmp26496 : tmp26499;
  assign tmp26493 = s3 ? tmp26494 : tmp26498;
  assign tmp26505 = s0 ? tmp23987 : tmp26384;
  assign tmp26504 = s1 ? tmp26490 : tmp26505;
  assign tmp26506 = s1 ? tmp26505 : tmp26483;
  assign tmp26503 = s2 ? tmp26504 : tmp26506;
  assign tmp26508 = s1 ? tmp26500 : tmp24535;
  assign tmp26507 = s2 ? tmp26508 : tmp24514;
  assign tmp26502 = s3 ? tmp26503 : tmp26507;
  assign tmp26492 = s4 ? tmp26493 : tmp26502;
  assign tmp26514 = l1 ? tmp24400 : tmp25983;
  assign tmp26513 = s0 ? tmp26472 : tmp26514;
  assign tmp26512 = s1 ? tmp26513 : tmp24514;
  assign tmp26516 = s0 ? tmp26501 : tmp26472;
  assign tmp26515 = s1 ? tmp26490 : tmp26516;
  assign tmp26511 = s2 ? tmp26512 : tmp26515;
  assign tmp26510 = s3 ? tmp26511 : tmp24545;
  assign tmp26520 = s0 ? tmp26514 : tmp26472;
  assign tmp26519 = s1 ? tmp26520 : tmp26500;
  assign tmp26518 = s2 ? tmp24536 : tmp26519;
  assign tmp26517 = s3 ? tmp26518 : tmp24553;
  assign tmp26509 = s4 ? tmp26510 : tmp26517;
  assign tmp26491 = s5 ? tmp26492 : tmp26509;
  assign tmp26468 = s6 ? tmp26469 : tmp26491;
  assign tmp26525 = s1 ? tmp26485 : tmp26475;
  assign tmp26524 = s2 ? tmp26482 : tmp26525;
  assign tmp26527 = s1 ? tmp26475 : tmp24514;
  assign tmp26526 = s2 ? tmp26527 : tmp26489;
  assign tmp26523 = s3 ? tmp26524 : tmp26526;
  assign tmp26522 = s4 ? tmp26470 : tmp26523;
  assign tmp26532 = s1 ? tmp26472 : tmp26478;
  assign tmp26531 = s2 ? tmp26477 : tmp26532;
  assign tmp26533 = s2 ? tmp26472 : tmp26499;
  assign tmp26530 = s3 ? tmp26531 : tmp26533;
  assign tmp26535 = s2 ? tmp26504 : tmp26472;
  assign tmp26537 = s1 ? tmp26500 : tmp24536;
  assign tmp26536 = s2 ? tmp26537 : tmp24514;
  assign tmp26534 = s3 ? tmp26535 : tmp26536;
  assign tmp26529 = s4 ? tmp26530 : tmp26534;
  assign tmp26541 = s1 ? tmp26472 : tmp24536;
  assign tmp26540 = s2 ? tmp26512 : tmp26541;
  assign tmp26542 = s2 ? tmp24514 : tmp24579;
  assign tmp26539 = s3 ? tmp26540 : tmp26542;
  assign tmp26544 = s2 ? tmp24514 : tmp26472;
  assign tmp26543 = s3 ? tmp26544 : tmp24536;
  assign tmp26538 = s4 ? tmp26539 : tmp26543;
  assign tmp26528 = s5 ? tmp26529 : tmp26538;
  assign tmp26521 = s6 ? tmp26522 : tmp26528;
  assign tmp26467 = s7 ? tmp26468 : tmp26521;
  assign tmp26550 = s2 ? tmp24628 : tmp26519;
  assign tmp26549 = s3 ? tmp26550 : tmp24553;
  assign tmp26548 = s4 ? tmp26510 : tmp26549;
  assign tmp26547 = s5 ? tmp26492 : tmp26548;
  assign tmp26546 = s6 ? tmp26469 : tmp26547;
  assign tmp26545 = s7 ? tmp26546 : tmp26521;
  assign tmp26466 = s8 ? tmp26467 : tmp26545;
  assign tmp26557 = s1 ? tmp26472 : tmp26516;
  assign tmp26556 = s2 ? tmp26488 : tmp26557;
  assign tmp26555 = s3 ? tmp26481 : tmp26556;
  assign tmp26554 = s4 ? tmp26470 : tmp26555;
  assign tmp26563 = s0 ? tmp26514 : tmp24514;
  assign tmp26562 = s1 ? tmp26563 : tmp26500;
  assign tmp26561 = s2 ? tmp26496 : tmp26562;
  assign tmp26560 = s3 ? tmp26494 : tmp26561;
  assign tmp26567 = s0 ? tmp26384 : tmp24536;
  assign tmp26566 = s1 ? tmp26500 : tmp26567;
  assign tmp26565 = s2 ? tmp26566 : tmp24514;
  assign tmp26564 = s3 ? tmp26503 : tmp26565;
  assign tmp26559 = s4 ? tmp26560 : tmp26564;
  assign tmp26571 = s1 ? tmp26513 : tmp26514;
  assign tmp26570 = s2 ? tmp26571 : tmp26516;
  assign tmp26569 = s3 ? tmp26570 : tmp24545;
  assign tmp26574 = s1 ? tmp24536 : tmp26514;
  assign tmp26573 = s2 ? tmp26574 : tmp26519;
  assign tmp26576 = s1 ? tmp26514 : tmp24549;
  assign tmp26575 = s2 ? tmp26576 : tmp24554;
  assign tmp26572 = s3 ? tmp26573 : tmp26575;
  assign tmp26568 = s4 ? tmp26569 : tmp26572;
  assign tmp26558 = s5 ? tmp26559 : tmp26568;
  assign tmp26553 = s6 ? tmp26554 : tmp26558;
  assign tmp26580 = s2 ? tmp26527 : tmp26557;
  assign tmp26579 = s3 ? tmp26524 : tmp26580;
  assign tmp26578 = s4 ? tmp26470 : tmp26579;
  assign tmp26584 = s2 ? tmp26472 : tmp26562;
  assign tmp26583 = s3 ? tmp26531 : tmp26584;
  assign tmp26582 = s4 ? tmp26583 : tmp26534;
  assign tmp26587 = s2 ? tmp26571 : tmp26557;
  assign tmp26586 = s3 ? tmp26587 : tmp24696;
  assign tmp26590 = s1 ? tmp26472 : tmp26500;
  assign tmp26589 = s2 ? tmp26514 : tmp26590;
  assign tmp26588 = s3 ? tmp26589 : tmp24536;
  assign tmp26585 = s4 ? tmp26586 : tmp26588;
  assign tmp26581 = s5 ? tmp26582 : tmp26585;
  assign tmp26577 = s6 ? tmp26578 : tmp26581;
  assign tmp26552 = s7 ? tmp26553 : tmp26577;
  assign tmp26551 = s8 ? tmp26545 : tmp26552;
  assign tmp26465 = s9 ? tmp26466 : tmp26551;
  assign tmp26598 = s1 ? tmp26472 : tmp26520;
  assign tmp26597 = s2 ? tmp26488 : tmp26598;
  assign tmp26596 = s3 ? tmp26481 : tmp26597;
  assign tmp26595 = s4 ? tmp26470 : tmp26596;
  assign tmp26603 = s1 ? tmp26520 : tmp26516;
  assign tmp26602 = s2 ? tmp26571 : tmp26603;
  assign tmp26601 = s3 ? tmp26602 : tmp24545;
  assign tmp26600 = s4 ? tmp26601 : tmp26572;
  assign tmp26599 = s5 ? tmp26559 : tmp26600;
  assign tmp26594 = s6 ? tmp26595 : tmp26599;
  assign tmp26607 = s2 ? tmp26527 : tmp26598;
  assign tmp26606 = s3 ? tmp26524 : tmp26607;
  assign tmp26605 = s4 ? tmp26470 : tmp26606;
  assign tmp26611 = s2 ? tmp26571 : tmp26541;
  assign tmp26610 = s3 ? tmp26611 : tmp26542;
  assign tmp26613 = s2 ? tmp26514 : tmp26472;
  assign tmp26612 = s3 ? tmp26613 : tmp24536;
  assign tmp26609 = s4 ? tmp26610 : tmp26612;
  assign tmp26608 = s5 ? tmp26582 : tmp26609;
  assign tmp26604 = s6 ? tmp26605 : tmp26608;
  assign tmp26593 = s7 ? tmp26594 : tmp26604;
  assign tmp26592 = s8 ? tmp26593 : tmp26594;
  assign tmp26622 = s0 ? tmp24588 : tmp26501;
  assign tmp26621 = s1 ? tmp24514 : tmp26622;
  assign tmp26620 = s2 ? tmp24588 : tmp26621;
  assign tmp26619 = s3 ? tmp24687 : tmp26620;
  assign tmp26625 = s1 ? tmp24602 : tmp26505;
  assign tmp26624 = s2 ? tmp26625 : tmp24588;
  assign tmp26627 = s1 ? tmp26622 : tmp24536;
  assign tmp26626 = s2 ? tmp26627 : tmp24514;
  assign tmp26623 = s3 ? tmp26624 : tmp26626;
  assign tmp26618 = s4 ? tmp26619 : tmp26623;
  assign tmp26632 = s0 ? tmp24588 : tmp26514;
  assign tmp26631 = s1 ? tmp26632 : tmp24514;
  assign tmp26630 = s2 ? tmp26631 : tmp24647;
  assign tmp26629 = s3 ? tmp26630 : tmp26542;
  assign tmp26628 = s4 ? tmp26629 : tmp24722;
  assign tmp26617 = s5 ? tmp26618 : tmp26628;
  assign tmp26616 = s6 ? tmp24683 : tmp26617;
  assign tmp26635 = s4 ? tmp26586 : tmp26612;
  assign tmp26634 = s5 ? tmp26582 : tmp26635;
  assign tmp26633 = s6 ? tmp26578 : tmp26634;
  assign tmp26615 = s7 ? tmp26616 : tmp26633;
  assign tmp26614 = s8 ? tmp26615 : tmp26604;
  assign tmp26591 = s9 ? tmp26592 : tmp26614;
  assign tmp26464 = s10 ? tmp26465 : tmp26591;
  assign tmp26639 = s7 ? tmp26616 : tmp26577;
  assign tmp26638 = s8 ? tmp26639 : tmp26604;
  assign tmp26637 = s9 ? tmp26592 : tmp26638;
  assign tmp26636 = s10 ? tmp26465 : tmp26637;
  assign tmp26463 = s11 ? tmp26464 : tmp26636;
  assign tmp26648 = s3 ? tmp24768 : tmp26542;
  assign tmp26647 = s4 ? tmp26648 : tmp24841;
  assign tmp26646 = s5 ? tmp24778 : tmp26647;
  assign tmp26645 = s6 ? tmp24773 : tmp26646;
  assign tmp26644 = s7 ? tmp24741 : tmp26645;
  assign tmp26651 = s5 ? tmp24808 : tmp26647;
  assign tmp26650 = s6 ? tmp24806 : tmp26651;
  assign tmp26649 = s7 ? tmp24791 : tmp26650;
  assign tmp26643 = s8 ? tmp26644 : tmp26649;
  assign tmp26652 = s8 ? tmp26649 : tmp24817;
  assign tmp26642 = s9 ? tmp26643 : tmp26652;
  assign tmp26657 = s5 ? tmp24826 : tmp26647;
  assign tmp26656 = s6 ? tmp24773 : tmp26657;
  assign tmp26655 = s7 ? tmp24818 : tmp26656;
  assign tmp26654 = s8 ? tmp26655 : tmp24818;
  assign tmp26661 = s5 ? tmp24826 : tmp24845;
  assign tmp26660 = s6 ? tmp24773 : tmp26661;
  assign tmp26659 = s7 ? tmp26645 : tmp26660;
  assign tmp26662 = s7 ? tmp26650 : tmp26656;
  assign tmp26658 = s8 ? tmp26659 : tmp26662;
  assign tmp26653 = s9 ? tmp26654 : tmp26658;
  assign tmp26641 = s10 ? tmp26642 : tmp26653;
  assign tmp26666 = s7 ? tmp26645 : tmp24824;
  assign tmp26665 = s8 ? tmp26666 : tmp26662;
  assign tmp26664 = s9 ? tmp26654 : tmp26665;
  assign tmp26663 = s10 ? tmp26642 : tmp26664;
  assign tmp26640 = s11 ? tmp26641 : tmp26663;
  assign tmp26462 = s12 ? tmp26463 : tmp26640;
  assign tmp26216 = s13 ? tmp26217 : tmp26462;
  assign tmp25950 = s14 ? tmp25951 : tmp26216;
  assign tmp26680 = s0 ? tmp25385 : tmp23982;
  assign tmp26679 = s1 ? tmp26680 : tmp25299;
  assign tmp26678 = s2 ? tmp25299 : tmp26679;
  assign tmp26677 = s3 ? tmp25429 : tmp26678;
  assign tmp26676 = s4 ? tmp26677 : tmp25434;
  assign tmp26686 = s0 ? tmp25299 : tmp24399;
  assign tmp26685 = s1 ? tmp25444 : tmp26686;
  assign tmp26684 = s2 ? tmp25442 : tmp26685;
  assign tmp26687 = s2 ? tmp25430 : tmp25448;
  assign tmp26683 = s3 ? tmp26684 : tmp26687;
  assign tmp26682 = s4 ? tmp26683 : tmp25449;
  assign tmp26681 = s5 ? tmp26682 : tmp25455;
  assign tmp26675 = s6 ? tmp26676 : tmp26681;
  assign tmp26689 = s4 ? tmp26677 : tmp25473;
  assign tmp26694 = s1 ? tmp25299 : tmp26686;
  assign tmp26693 = s2 ? tmp25481 : tmp26694;
  assign tmp26692 = s3 ? tmp26693 : tmp25483;
  assign tmp26697 = s1 ? tmp24399 : tmp25299;
  assign tmp26696 = s2 ? tmp25451 : tmp26697;
  assign tmp26695 = s3 ? tmp26696 : tmp25454;
  assign tmp26691 = s4 ? tmp26692 : tmp26695;
  assign tmp26700 = s2 ? tmp25071 : tmp25492;
  assign tmp26699 = s3 ? tmp25489 : tmp26700;
  assign tmp26701 = s3 ? tmp25496 : tmp25497;
  assign tmp26698 = s4 ? tmp26699 : tmp26701;
  assign tmp26690 = s5 ? tmp26691 : tmp26698;
  assign tmp26688 = s6 ? tmp26689 : tmp26690;
  assign tmp26674 = s7 ? tmp26675 : tmp26688;
  assign tmp26708 = s0 ? tmp25385 : tmp25299;
  assign tmp26707 = s1 ? tmp26708 : tmp25299;
  assign tmp26709 = s1 ? tmp25384 : tmp25299;
  assign tmp26706 = s2 ? tmp26707 : tmp26709;
  assign tmp26705 = s3 ? tmp25429 : tmp26706;
  assign tmp26704 = s4 ? tmp26705 : tmp25434;
  assign tmp26715 = s0 ? tmp25299 : tmp24514;
  assign tmp26714 = s1 ? tmp25444 : tmp26715;
  assign tmp26713 = s2 ? tmp25442 : tmp26714;
  assign tmp26717 = s0 ? tmp24514 : tmp25299;
  assign tmp26718 = s1 ? tmp25395 : tmp25299;
  assign tmp26716 = s2 ? tmp26717 : tmp26718;
  assign tmp26712 = s3 ? tmp26713 : tmp26716;
  assign tmp26721 = s1 ? tmp25452 : tmp24419;
  assign tmp26722 = s1 ? tmp24419 : tmp25433;
  assign tmp26720 = s2 ? tmp26721 : tmp26722;
  assign tmp26719 = s3 ? tmp26720 : tmp25454;
  assign tmp26711 = s4 ? tmp26712 : tmp26719;
  assign tmp26726 = s1 ? tmp25465 : tmp25405;
  assign tmp26725 = s2 ? tmp26726 : tmp25466;
  assign tmp26724 = s3 ? tmp26725 : tmp25467;
  assign tmp26723 = s4 ? tmp25456 : tmp26724;
  assign tmp26710 = s5 ? tmp26711 : tmp26723;
  assign tmp26703 = s6 ? tmp26704 : tmp26710;
  assign tmp26730 = s2 ? tmp25410 : tmp25299;
  assign tmp26729 = s3 ? tmp25474 : tmp26730;
  assign tmp26728 = s4 ? tmp26705 : tmp26729;
  assign tmp26735 = s1 ? tmp25299 : tmp26715;
  assign tmp26734 = s2 ? tmp25481 : tmp26735;
  assign tmp26736 = s2 ? tmp25299 : tmp26718;
  assign tmp26733 = s3 ? tmp26734 : tmp26736;
  assign tmp26738 = s2 ? tmp26721 : tmp25299;
  assign tmp26737 = s3 ? tmp26738 : tmp25486;
  assign tmp26732 = s4 ? tmp26733 : tmp26737;
  assign tmp26742 = s1 ? tmp25337 : tmp25396;
  assign tmp26741 = s2 ? tmp26742 : tmp25299;
  assign tmp26740 = s3 ? tmp26741 : tmp25497;
  assign tmp26739 = s4 ? tmp26699 : tmp26740;
  assign tmp26731 = s5 ? tmp26732 : tmp26739;
  assign tmp26727 = s6 ? tmp26728 : tmp26731;
  assign tmp26702 = s7 ? tmp26703 : tmp26727;
  assign tmp26673 = s8 ? tmp26674 : tmp26702;
  assign tmp26751 = s0 ? tmp25299 : tmp24400;
  assign tmp26750 = s1 ? tmp25444 : tmp26751;
  assign tmp26749 = s2 ? tmp25442 : tmp26750;
  assign tmp26753 = s0 ? tmp24400 : tmp25299;
  assign tmp26752 = s2 ? tmp26753 : tmp25448;
  assign tmp26748 = s3 ? tmp26749 : tmp26752;
  assign tmp26747 = s4 ? tmp26748 : tmp25449;
  assign tmp26746 = s5 ? tmp26747 : tmp25455;
  assign tmp26745 = s6 ? tmp25427 : tmp26746;
  assign tmp26759 = s1 ? tmp25299 : tmp26751;
  assign tmp26758 = s2 ? tmp25481 : tmp26759;
  assign tmp26757 = s3 ? tmp26758 : tmp25483;
  assign tmp26756 = s4 ? tmp26757 : tmp25484;
  assign tmp26755 = s5 ? tmp26756 : tmp25487;
  assign tmp26754 = s6 ? tmp25472 : tmp26755;
  assign tmp26744 = s7 ? tmp26745 : tmp26754;
  assign tmp26743 = s8 ? tmp26702 : tmp26744;
  assign tmp26672 = s9 ? tmp26673 : tmp26743;
  assign tmp26763 = s6 ? tmp26676 : tmp26746;
  assign tmp26765 = s5 ? tmp26756 : tmp26698;
  assign tmp26764 = s6 ? tmp26689 : tmp26765;
  assign tmp26762 = s7 ? tmp26763 : tmp26764;
  assign tmp26761 = s8 ? tmp26762 : tmp26763;
  assign tmp26771 = s3 ? tmp26696 : tmp25486;
  assign tmp26770 = s4 ? tmp26692 : tmp26771;
  assign tmp26769 = s5 ? tmp26770 : tmp26698;
  assign tmp26768 = s6 ? tmp26689 : tmp26769;
  assign tmp26773 = s5 ? tmp26756 : tmp25529;
  assign tmp26772 = s6 ? tmp25472 : tmp26773;
  assign tmp26767 = s7 ? tmp26768 : tmp26772;
  assign tmp26774 = s7 ? tmp26727 : tmp26764;
  assign tmp26766 = s8 ? tmp26767 : tmp26774;
  assign tmp26760 = s9 ? tmp26761 : tmp26766;
  assign tmp26671 = s10 ? tmp26672 : tmp26760;
  assign tmp26778 = s7 ? tmp26688 : tmp26754;
  assign tmp26777 = s8 ? tmp26778 : tmp26774;
  assign tmp26776 = s9 ? tmp26761 : tmp26777;
  assign tmp26775 = s10 ? tmp26672 : tmp26776;
  assign tmp26670 = s11 ? tmp26671 : tmp26775;
  assign tmp26789 = s0 ? tmp24400 : tmp26248;
  assign tmp26788 = s1 ? tmp26789 : tmp25553;
  assign tmp26787 = s2 ? tmp26788 : tmp25565;
  assign tmp26786 = s3 ? tmp26787 : tmp25566;
  assign tmp26785 = s4 ? tmp25551 : tmp26786;
  assign tmp26795 = s0 ? tmp25553 : tmp26514;
  assign tmp26794 = s1 ? tmp26795 : tmp24514;
  assign tmp26797 = s0 ? tmp26514 : tmp25553;
  assign tmp26796 = s1 ? tmp26797 : tmp25560;
  assign tmp26793 = s2 ? tmp26794 : tmp26796;
  assign tmp26792 = s3 ? tmp26793 : tmp25575;
  assign tmp26801 = s0 ? tmp26248 : tmp24410;
  assign tmp26800 = s1 ? tmp25581 : tmp26801;
  assign tmp26802 = s1 ? tmp26801 : tmp26789;
  assign tmp26799 = s2 ? tmp26800 : tmp26802;
  assign tmp26798 = s3 ? tmp26799 : tmp25584;
  assign tmp26791 = s4 ? tmp26792 : tmp26798;
  assign tmp26790 = s5 ? tmp26791 : tmp25587;
  assign tmp26784 = s6 ? tmp26785 : tmp26790;
  assign tmp26805 = s3 ? tmp26787 : tmp25610;
  assign tmp26804 = s4 ? tmp25551 : tmp26805;
  assign tmp26809 = s2 ? tmp26794 : tmp25616;
  assign tmp26808 = s3 ? tmp26809 : tmp25617;
  assign tmp26811 = s2 ? tmp26800 : tmp24400;
  assign tmp26810 = s3 ? tmp26811 : tmp25620;
  assign tmp26807 = s4 ? tmp26808 : tmp26810;
  assign tmp26806 = s5 ? tmp26807 : tmp25622;
  assign tmp26803 = s6 ? tmp26804 : tmp26806;
  assign tmp26783 = s7 ? tmp26784 : tmp26803;
  assign tmp26817 = l1 ? tmp25554 : tmp26336;
  assign tmp26818 = s0 ? tmp26349 : tmp26817;
  assign tmp26816 = s1 ? tmp26817 : tmp26818;
  assign tmp26821 = s0 ? tmp24514 : tmp26817;
  assign tmp26820 = s1 ? tmp26821 : tmp26817;
  assign tmp26823 = s0 ? tmp26817 : tmp26349;
  assign tmp26822 = s1 ? tmp26823 : tmp26817;
  assign tmp26819 = s2 ? tmp26820 : tmp26822;
  assign tmp26815 = s3 ? tmp26816 : tmp26819;
  assign tmp26828 = l1 ? tmp24400 : tmp26336;
  assign tmp26827 = s0 ? tmp26828 : tmp26248;
  assign tmp26826 = s1 ? tmp26827 : tmp26817;
  assign tmp26830 = s0 ? tmp26817 : tmp24410;
  assign tmp26829 = s1 ? tmp26830 : tmp26365;
  assign tmp26825 = s2 ? tmp26826 : tmp26829;
  assign tmp26832 = s1 ? tmp26349 : tmp25046;
  assign tmp26831 = s2 ? tmp26832 : tmp26817;
  assign tmp26824 = s3 ? tmp26825 : tmp26831;
  assign tmp26814 = s4 ? tmp26815 : tmp26824;
  assign tmp26838 = s0 ? tmp26817 : tmp26514;
  assign tmp26837 = s1 ? tmp26838 : tmp24514;
  assign tmp26840 = s0 ? tmp26514 : tmp26817;
  assign tmp26839 = s1 ? tmp26840 : tmp26823;
  assign tmp26836 = s2 ? tmp26837 : tmp26839;
  assign tmp26843 = s0 ? tmp26817 : tmp24870;
  assign tmp26842 = s1 ? tmp26843 : tmp26817;
  assign tmp26841 = s2 ? tmp26818 : tmp26842;
  assign tmp26835 = s3 ? tmp26836 : tmp26841;
  assign tmp26847 = s0 ? tmp25026 : tmp26817;
  assign tmp26848 = s0 ? tmp26248 : tmp26349;
  assign tmp26846 = s1 ? tmp26847 : tmp26848;
  assign tmp26849 = s1 ? tmp26848 : tmp26827;
  assign tmp26845 = s2 ? tmp26846 : tmp26849;
  assign tmp26852 = s0 ? tmp26349 : tmp25553;
  assign tmp26851 = s1 ? tmp26817 : tmp26852;
  assign tmp26850 = s2 ? tmp26851 : tmp25585;
  assign tmp26844 = s3 ? tmp26845 : tmp26850;
  assign tmp26834 = s4 ? tmp26835 : tmp26844;
  assign tmp26857 = s0 ? tmp24870 : tmp26817;
  assign tmp26856 = s1 ? tmp26843 : tmp26857;
  assign tmp26859 = s0 ? tmp26817 : tmp24514;
  assign tmp26858 = s1 ? tmp26859 : tmp24514;
  assign tmp26855 = s2 ? tmp26856 : tmp26858;
  assign tmp26854 = s3 ? tmp26855 : tmp25592;
  assign tmp26863 = s0 ? tmp25553 : tmp26817;
  assign tmp26862 = s1 ? tmp25600 : tmp26863;
  assign tmp26864 = s1 ? tmp26857 : tmp24514;
  assign tmp26861 = s2 ? tmp26862 : tmp26864;
  assign tmp26867 = s0 ? tmp26817 : tmp25553;
  assign tmp26866 = s1 ? tmp26867 : tmp25591;
  assign tmp26865 = s2 ? tmp26866 : tmp25605;
  assign tmp26860 = s3 ? tmp26861 : tmp26865;
  assign tmp26853 = s4 ? tmp26854 : tmp26860;
  assign tmp26833 = s5 ? tmp26834 : tmp26853;
  assign tmp26813 = s6 ? tmp26814 : tmp26833;
  assign tmp26872 = s1 ? tmp26830 : tmp26349;
  assign tmp26871 = s2 ? tmp26826 : tmp26872;
  assign tmp26874 = s1 ? tmp26349 : tmp25026;
  assign tmp26873 = s2 ? tmp26874 : tmp26817;
  assign tmp26870 = s3 ? tmp26871 : tmp26873;
  assign tmp26869 = s4 ? tmp26815 : tmp26870;
  assign tmp26879 = s1 ? tmp26817 : tmp26823;
  assign tmp26878 = s2 ? tmp26837 : tmp26879;
  assign tmp26880 = s2 ? tmp26817 : tmp26842;
  assign tmp26877 = s3 ? tmp26878 : tmp26880;
  assign tmp26882 = s2 ? tmp26846 : tmp26828;
  assign tmp26884 = s1 ? tmp26817 : tmp25553;
  assign tmp26883 = s2 ? tmp26884 : tmp25621;
  assign tmp26881 = s3 ? tmp26882 : tmp26883;
  assign tmp26876 = s4 ? tmp26877 : tmp26881;
  assign tmp26887 = s2 ? tmp26842 : tmp26858;
  assign tmp26886 = s3 ? tmp26887 : tmp25625;
  assign tmp26890 = s1 ? tmp25553 : tmp26817;
  assign tmp26889 = s2 ? tmp26890 : tmp26817;
  assign tmp26891 = s1 ? tmp26867 : tmp25553;
  assign tmp26888 = s3 ? tmp26889 : tmp26891;
  assign tmp26885 = s4 ? tmp26886 : tmp26888;
  assign tmp26875 = s5 ? tmp26876 : tmp26885;
  assign tmp26868 = s6 ? tmp26869 : tmp26875;
  assign tmp26812 = s7 ? tmp26813 : tmp26868;
  assign tmp26782 = s8 ? tmp26783 : tmp26812;
  assign tmp26899 = s0 ? tmp26817 : tmp26828;
  assign tmp26898 = s1 ? tmp26899 : tmp26817;
  assign tmp26897 = s2 ? tmp26820 : tmp26898;
  assign tmp26896 = s3 ? tmp26816 : tmp26897;
  assign tmp26903 = s0 ? tmp26828 : tmp26514;
  assign tmp26902 = s1 ? tmp26903 : tmp26817;
  assign tmp26901 = s2 ? tmp26902 : tmp26829;
  assign tmp26900 = s3 ? tmp26901 : tmp26831;
  assign tmp26895 = s4 ? tmp26896 : tmp26900;
  assign tmp26908 = s1 ? tmp26840 : tmp26899;
  assign tmp26907 = s2 ? tmp26837 : tmp26908;
  assign tmp26910 = s0 ? tmp26828 : tmp26817;
  assign tmp26909 = s2 ? tmp26910 : tmp26842;
  assign tmp26906 = s3 ? tmp26907 : tmp26909;
  assign tmp26913 = s1 ? tmp26848 : tmp26903;
  assign tmp26912 = s2 ? tmp26846 : tmp26913;
  assign tmp26911 = s3 ? tmp26912 : tmp26850;
  assign tmp26905 = s4 ? tmp26906 : tmp26911;
  assign tmp26904 = s5 ? tmp26905 : tmp26853;
  assign tmp26894 = s6 ? tmp26895 : tmp26904;
  assign tmp26917 = s2 ? tmp26902 : tmp26872;
  assign tmp26916 = s3 ? tmp26917 : tmp26873;
  assign tmp26915 = s4 ? tmp26896 : tmp26916;
  assign tmp26922 = s1 ? tmp26817 : tmp26899;
  assign tmp26921 = s2 ? tmp26837 : tmp26922;
  assign tmp26920 = s3 ? tmp26921 : tmp26880;
  assign tmp26919 = s4 ? tmp26920 : tmp26881;
  assign tmp26918 = s5 ? tmp26919 : tmp26885;
  assign tmp26914 = s6 ? tmp26915 : tmp26918;
  assign tmp26893 = s7 ? tmp26894 : tmp26914;
  assign tmp26927 = s2 ? tmp26817 : tmp26822;
  assign tmp26926 = s3 ? tmp26816 : tmp26927;
  assign tmp26925 = s4 ? tmp26926 : tmp26900;
  assign tmp26932 = s1 ? tmp26838 : tmp26514;
  assign tmp26931 = s2 ? tmp26932 : tmp26839;
  assign tmp26930 = s3 ? tmp26931 : tmp26841;
  assign tmp26929 = s4 ? tmp26930 : tmp26911;
  assign tmp26938 = l1 ? tmp25554 : tmp25983;
  assign tmp26937 = s0 ? tmp25553 : tmp26938;
  assign tmp26936 = s1 ? tmp26817 : tmp26937;
  assign tmp26935 = s2 ? tmp26856 : tmp26936;
  assign tmp26934 = s3 ? tmp26935 : tmp25592;
  assign tmp26942 = s0 ? tmp26514 : tmp24400;
  assign tmp26941 = s1 ? tmp26857 : tmp26942;
  assign tmp26940 = s2 ? tmp26862 : tmp26941;
  assign tmp26939 = s3 ? tmp26940 : tmp26865;
  assign tmp26933 = s4 ? tmp26934 : tmp26939;
  assign tmp26928 = s5 ? tmp26929 : tmp26933;
  assign tmp26924 = s6 ? tmp26925 : tmp26928;
  assign tmp26944 = s4 ? tmp26926 : tmp26916;
  assign tmp26948 = s2 ? tmp26932 : tmp26879;
  assign tmp26947 = s3 ? tmp26948 : tmp26880;
  assign tmp26946 = s4 ? tmp26947 : tmp26881;
  assign tmp26952 = s1 ? tmp26817 : tmp24514;
  assign tmp26951 = s2 ? tmp26842 : tmp26952;
  assign tmp26950 = s3 ? tmp26951 : tmp25625;
  assign tmp26949 = s4 ? tmp26950 : tmp26888;
  assign tmp26945 = s5 ? tmp26946 : tmp26949;
  assign tmp26943 = s6 ? tmp26944 : tmp26945;
  assign tmp26923 = s7 ? tmp26924 : tmp26943;
  assign tmp26892 = s8 ? tmp26893 : tmp26923;
  assign tmp26781 = s9 ? tmp26782 : tmp26892;
  assign tmp26962 = s0 ? tmp24400 : tmp26514;
  assign tmp26961 = s1 ? tmp26899 : tmp26962;
  assign tmp26960 = s2 ? tmp26856 : tmp26961;
  assign tmp26959 = s3 ? tmp26960 : tmp25592;
  assign tmp26958 = s4 ? tmp26959 : tmp26939;
  assign tmp26957 = s5 ? tmp26929 : tmp26958;
  assign tmp26956 = s6 ? tmp26925 : tmp26957;
  assign tmp26968 = s1 ? tmp26899 : tmp24514;
  assign tmp26967 = s2 ? tmp26842 : tmp26968;
  assign tmp26966 = s3 ? tmp26967 : tmp25625;
  assign tmp26965 = s4 ? tmp26966 : tmp26888;
  assign tmp26964 = s5 ? tmp26946 : tmp26965;
  assign tmp26963 = s6 ? tmp26944 : tmp26964;
  assign tmp26955 = s7 ? tmp26956 : tmp26963;
  assign tmp26954 = s8 ? tmp26955 : tmp26956;
  assign tmp26972 = s5 ? tmp26807 : tmp25706;
  assign tmp26971 = s6 ? tmp26804 : tmp26972;
  assign tmp26976 = s3 ? tmp26889 : tmp25553;
  assign tmp26975 = s4 ? tmp26950 : tmp26976;
  assign tmp26974 = s5 ? tmp26946 : tmp26975;
  assign tmp26973 = s6 ? tmp26944 : tmp26974;
  assign tmp26970 = s7 ? tmp26971 : tmp26973;
  assign tmp26980 = s3 ? tmp26889 : tmp25671;
  assign tmp26979 = s4 ? tmp26966 : tmp26980;
  assign tmp26978 = s5 ? tmp26946 : tmp26979;
  assign tmp26977 = s6 ? tmp26944 : tmp26978;
  assign tmp26969 = s8 ? tmp26970 : tmp26977;
  assign tmp26953 = s9 ? tmp26954 : tmp26969;
  assign tmp26780 = s10 ? tmp26781 : tmp26953;
  assign tmp26984 = s7 ? tmp26803 : tmp26943;
  assign tmp26983 = s8 ? tmp26984 : tmp26963;
  assign tmp26982 = s9 ? tmp26954 : tmp26983;
  assign tmp26981 = s10 ? tmp26781 : tmp26982;
  assign tmp26779 = s11 ? tmp26780 : tmp26981;
  assign tmp26669 = s12 ? tmp26670 : tmp26779;
  assign tmp26668 = s13 ? tmp26669 : tmp25712;
  assign tmp26667 = s14 ? tmp24859 : tmp26668;
  assign tmp25949 = s15 ? tmp25950 : tmp26667;
  assign tmp23952 = s16 ? tmp23953 : tmp25949;
  assign tmp26992 = s8 ? tmp25974 : tmp24057;
  assign tmp26991 = s9 ? tmp25955 : tmp26992;
  assign tmp26994 = s8 ? tmp25956 : tmp25957;
  assign tmp26996 = s7 ? tmp25969 : tmp24066;
  assign tmp26997 = s7 ? tmp26083 : tmp25969;
  assign tmp26995 = s8 ? tmp26996 : tmp26997;
  assign tmp26993 = s9 ? tmp26994 : tmp26995;
  assign tmp26990 = s10 ? tmp26991 : tmp26993;
  assign tmp27001 = s7 ? tmp25986 : tmp25969;
  assign tmp27000 = s8 ? tmp26996 : tmp27001;
  assign tmp26999 = s9 ? tmp26994 : tmp27000;
  assign tmp26998 = s10 ? tmp26991 : tmp26999;
  assign tmp26989 = s11 ? tmp26990 : tmp26998;
  assign tmp27010 = s3 ? tmp24298 : tmp26200;
  assign tmp27009 = s4 ? tmp23973 : tmp27010;
  assign tmp27008 = s6 ? tmp27009 : tmp26122;
  assign tmp27007 = s7 ? tmp26099 : tmp27008;
  assign tmp27006 = s8 ? tmp26129 : tmp27007;
  assign tmp27005 = s9 ? tmp26097 : tmp27006;
  assign tmp27012 = s8 ? tmp27007 : tmp26099;
  assign tmp27014 = s7 ? tmp26197 : tmp27008;
  assign tmp27015 = s7 ? tmp26207 : tmp27008;
  assign tmp27013 = s8 ? tmp27014 : tmp27015;
  assign tmp27011 = s9 ? tmp27012 : tmp27013;
  assign tmp27004 = s10 ? tmp27005 : tmp27011;
  assign tmp27019 = s7 ? tmp26121 : tmp27008;
  assign tmp27020 = s7 ? tmp26143 : tmp27008;
  assign tmp27018 = s8 ? tmp27019 : tmp27020;
  assign tmp27017 = s9 ? tmp27012 : tmp27018;
  assign tmp27016 = s10 ? tmp27005 : tmp27017;
  assign tmp27003 = s11 ? tmp27004 : tmp27016;
  assign tmp27002 = s12 ? tmp24077 : tmp27003;
  assign tmp26988 = s13 ? tmp26989 : tmp27002;
  assign tmp27026 = s8 ? tmp26222 : tmp24373;
  assign tmp27025 = s9 ? tmp26221 : tmp27026;
  assign tmp27029 = s7 ? tmp26286 : tmp24362;
  assign tmp27028 = s8 ? tmp24384 : tmp27029;
  assign tmp27027 = s9 ? tmp24382 : tmp27028;
  assign tmp27024 = s10 ? tmp27025 : tmp27027;
  assign tmp27033 = s7 ? tmp26260 : tmp24362;
  assign tmp27032 = s8 ? tmp24362 : tmp27033;
  assign tmp27031 = s9 ? tmp24382 : tmp27032;
  assign tmp27030 = s10 ? tmp27025 : tmp27031;
  assign tmp27023 = s11 ? tmp27024 : tmp27030;
  assign tmp27042 = s2 ? tmp24399 : tmp26306;
  assign tmp27041 = s3 ? tmp27042 : tmp26309;
  assign tmp27040 = s4 ? tmp26303 : tmp27041;
  assign tmp27044 = s4 ? tmp26314 : tmp24451;
  assign tmp27043 = s5 ? tmp27044 : tmp24427;
  assign tmp27039 = s6 ? tmp27040 : tmp27043;
  assign tmp27047 = s3 ? tmp26304 : tmp24445;
  assign tmp27046 = s4 ? tmp26303 : tmp27047;
  assign tmp27045 = s6 ? tmp27046 : tmp26325;
  assign tmp27038 = s7 ? tmp27039 : tmp27045;
  assign tmp27037 = s8 ? tmp26331 : tmp27038;
  assign tmp27036 = s9 ? tmp26299 : tmp27037;
  assign tmp27049 = s8 ? tmp26300 : tmp26301;
  assign tmp27051 = s7 ? tmp26321 : tmp27045;
  assign tmp27052 = s7 ? tmp26455 : tmp26321;
  assign tmp27050 = s8 ? tmp27051 : tmp27052;
  assign tmp27048 = s9 ? tmp27049 : tmp27050;
  assign tmp27035 = s10 ? tmp27036 : tmp27048;
  assign tmp27056 = s7 ? tmp26392 : tmp26321;
  assign tmp27055 = s8 ? tmp27051 : tmp27056;
  assign tmp27054 = s9 ? tmp27049 : tmp27055;
  assign tmp27053 = s10 ? tmp27036 : tmp27054;
  assign tmp27034 = s11 ? tmp27035 : tmp27053;
  assign tmp27022 = s12 ? tmp27023 : tmp27034;
  assign tmp27068 = ~(l2 ? tmp23968 : tmp24501);
  assign tmp27067 = l1 ? tmp24499 : tmp27068;
  assign tmp27069 = s0 ? tmp26475 : tmp27067;
  assign tmp27066 = s1 ? tmp27067 : tmp27069;
  assign tmp27072 = s0 ? tmp27067 : tmp26479;
  assign tmp27071 = s1 ? tmp27072 : tmp27067;
  assign tmp27070 = s2 ? tmp27067 : tmp27071;
  assign tmp27065 = s3 ? tmp27066 : tmp27070;
  assign tmp27076 = s0 ? tmp27067 : tmp26475;
  assign tmp27075 = s1 ? tmp27076 : tmp27067;
  assign tmp27078 = s0 ? tmp27067 : tmp23997;
  assign tmp27077 = s1 ? tmp27078 : tmp26486;
  assign tmp27074 = s2 ? tmp27075 : tmp27077;
  assign tmp27081 = s0 ? tmp24514 : tmp27067;
  assign tmp27080 = s1 ? tmp27067 : tmp27081;
  assign tmp27079 = s2 ? tmp26488 : tmp27080;
  assign tmp27073 = s3 ? tmp27074 : tmp27079;
  assign tmp27064 = s4 ? tmp27065 : tmp27073;
  assign tmp27087 = s0 ? tmp26479 : tmp27067;
  assign tmp27086 = s1 ? tmp27072 : tmp27087;
  assign tmp27088 = s1 ? tmp27087 : tmp27072;
  assign tmp27085 = s2 ? tmp27086 : tmp27088;
  assign tmp27091 = s0 ? tmp27067 : tmp24527;
  assign tmp27090 = s1 ? tmp24514 : tmp27091;
  assign tmp27089 = s2 ? tmp27087 : tmp27090;
  assign tmp27084 = s3 ? tmp27085 : tmp27089;
  assign tmp27096 = l1 ? tmp24400 : tmp23983;
  assign tmp27095 = s0 ? tmp27096 : tmp27067;
  assign tmp27094 = s1 ? tmp27095 : tmp24531;
  assign tmp27097 = s1 ? tmp24531 : tmp27076;
  assign tmp27093 = s2 ? tmp27094 : tmp27097;
  assign tmp27099 = s1 ? tmp27091 : tmp24535;
  assign tmp27098 = s2 ? tmp27099 : tmp24514;
  assign tmp27092 = s3 ? tmp27093 : tmp27098;
  assign tmp27083 = s4 ? tmp27084 : tmp27092;
  assign tmp27104 = s0 ? tmp27067 : tmp26514;
  assign tmp27103 = s1 ? tmp27104 : tmp24514;
  assign tmp27106 = s0 ? tmp24536 : tmp27067;
  assign tmp27107 = s0 ? tmp24527 : tmp27067;
  assign tmp27105 = s1 ? tmp27106 : tmp27107;
  assign tmp27102 = s2 ? tmp27103 : tmp27105;
  assign tmp27101 = s3 ? tmp27102 : tmp24545;
  assign tmp27111 = s0 ? tmp26514 : tmp27067;
  assign tmp27110 = s1 ? tmp27111 : tmp27091;
  assign tmp27109 = s2 ? tmp24536 : tmp27110;
  assign tmp27108 = s3 ? tmp27109 : tmp24553;
  assign tmp27100 = s4 ? tmp27101 : tmp27108;
  assign tmp27082 = s5 ? tmp27083 : tmp27100;
  assign tmp27063 = s6 ? tmp27064 : tmp27082;
  assign tmp27116 = s1 ? tmp27078 : tmp26475;
  assign tmp27115 = s2 ? tmp27075 : tmp27116;
  assign tmp27117 = s2 ? tmp26527 : tmp27080;
  assign tmp27114 = s3 ? tmp27115 : tmp27117;
  assign tmp27113 = s4 ? tmp27065 : tmp27114;
  assign tmp27122 = s1 ? tmp27067 : tmp27072;
  assign tmp27121 = s2 ? tmp27071 : tmp27122;
  assign tmp27123 = s2 ? tmp27067 : tmp27090;
  assign tmp27120 = s3 ? tmp27121 : tmp27123;
  assign tmp27125 = s2 ? tmp27094 : tmp27067;
  assign tmp27127 = s1 ? tmp27091 : tmp24536;
  assign tmp27126 = s2 ? tmp27127 : tmp24514;
  assign tmp27124 = s3 ? tmp27125 : tmp27126;
  assign tmp27119 = s4 ? tmp27120 : tmp27124;
  assign tmp27131 = s1 ? tmp27067 : tmp27107;
  assign tmp27130 = s2 ? tmp27103 : tmp27131;
  assign tmp27129 = s3 ? tmp27130 : tmp24576;
  assign tmp27134 = s1 ? tmp27067 : tmp27091;
  assign tmp27133 = s2 ? tmp24514 : tmp27134;
  assign tmp27132 = s3 ? tmp27133 : tmp24536;
  assign tmp27128 = s4 ? tmp27129 : tmp27132;
  assign tmp27118 = s5 ? tmp27119 : tmp27128;
  assign tmp27112 = s6 ? tmp27113 : tmp27118;
  assign tmp27062 = s7 ? tmp27063 : tmp27112;
  assign tmp27143 = l1 ? tmp24499 : tmp23984;
  assign tmp27142 = s0 ? tmp27067 : tmp27143;
  assign tmp27141 = s1 ? tmp24514 : tmp27142;
  assign tmp27140 = s2 ? tmp27087 : tmp27141;
  assign tmp27139 = s3 ? tmp27085 : tmp27140;
  assign tmp27146 = s1 ? tmp27095 : tmp26505;
  assign tmp27147 = s1 ? tmp26505 : tmp27076;
  assign tmp27145 = s2 ? tmp27146 : tmp27147;
  assign tmp27149 = s1 ? tmp27142 : tmp24535;
  assign tmp27148 = s2 ? tmp27149 : tmp24514;
  assign tmp27144 = s3 ? tmp27145 : tmp27148;
  assign tmp27138 = s4 ? tmp27139 : tmp27144;
  assign tmp27153 = s1 ? tmp27081 : tmp27107;
  assign tmp27152 = s2 ? tmp27103 : tmp27153;
  assign tmp27151 = s3 ? tmp27152 : tmp24545;
  assign tmp27155 = s2 ? tmp24628 : tmp27110;
  assign tmp27154 = s3 ? tmp27155 : tmp24553;
  assign tmp27150 = s4 ? tmp27151 : tmp27154;
  assign tmp27137 = s5 ? tmp27138 : tmp27150;
  assign tmp27136 = s6 ? tmp27064 : tmp27137;
  assign tmp27160 = s2 ? tmp27067 : tmp27141;
  assign tmp27159 = s3 ? tmp27121 : tmp27160;
  assign tmp27162 = s2 ? tmp27146 : tmp27067;
  assign tmp27164 = s1 ? tmp27142 : tmp24536;
  assign tmp27163 = s2 ? tmp27164 : tmp24514;
  assign tmp27161 = s3 ? tmp27162 : tmp27163;
  assign tmp27158 = s4 ? tmp27159 : tmp27161;
  assign tmp27157 = s5 ? tmp27158 : tmp27128;
  assign tmp27156 = s6 ? tmp27113 : tmp27157;
  assign tmp27135 = s7 ? tmp27136 : tmp27156;
  assign tmp27061 = s8 ? tmp27062 : tmp27135;
  assign tmp27173 = s0 ? tmp24588 : tmp27143;
  assign tmp27172 = s1 ? tmp24514 : tmp27173;
  assign tmp27171 = s2 ? tmp24608 : tmp27172;
  assign tmp27170 = s3 ? tmp24663 : tmp27171;
  assign tmp27177 = s0 ? tmp27096 : tmp24588;
  assign tmp27176 = s1 ? tmp27177 : tmp24531;
  assign tmp27175 = s2 ? tmp27176 : tmp24671;
  assign tmp27179 = s1 ? tmp27173 : tmp24535;
  assign tmp27178 = s2 ? tmp27179 : tmp24514;
  assign tmp27174 = s3 ? tmp27175 : tmp27178;
  assign tmp27169 = s4 ? tmp27170 : tmp27174;
  assign tmp27184 = s0 ? tmp27143 : tmp24588;
  assign tmp27183 = s1 ? tmp24625 : tmp27184;
  assign tmp27182 = s2 ? tmp26631 : tmp27183;
  assign tmp27181 = s3 ? tmp27182 : tmp24545;
  assign tmp27188 = s0 ? tmp26514 : tmp24588;
  assign tmp27187 = s1 ? tmp27188 : tmp27173;
  assign tmp27186 = s2 ? tmp24536 : tmp27187;
  assign tmp27185 = s3 ? tmp27186 : tmp24553;
  assign tmp27180 = s4 ? tmp27181 : tmp27185;
  assign tmp27168 = s5 ? tmp27169 : tmp27180;
  assign tmp27167 = s6 ? tmp24657 : tmp27168;
  assign tmp27193 = s2 ? tmp24588 : tmp27172;
  assign tmp27192 = s3 ? tmp24687 : tmp27193;
  assign tmp27195 = s2 ? tmp27176 : tmp24588;
  assign tmp27197 = s1 ? tmp27173 : tmp24536;
  assign tmp27196 = s2 ? tmp27197 : tmp24514;
  assign tmp27194 = s3 ? tmp27195 : tmp27196;
  assign tmp27191 = s4 ? tmp27192 : tmp27194;
  assign tmp27199 = s3 ? tmp26630 : tmp24696;
  assign tmp27202 = s1 ? tmp24588 : tmp27143;
  assign tmp27201 = s2 ? tmp24514 : tmp27202;
  assign tmp27200 = s3 ? tmp27201 : tmp24536;
  assign tmp27198 = s4 ? tmp27199 : tmp27200;
  assign tmp27190 = s5 ? tmp27191 : tmp27198;
  assign tmp27189 = s6 ? tmp24683 : tmp27190;
  assign tmp27166 = s7 ? tmp27167 : tmp27189;
  assign tmp27165 = s8 ? tmp27135 : tmp27166;
  assign tmp27060 = s9 ? tmp27061 : tmp27165;
  assign tmp27212 = s0 ? tmp27096 : tmp24498;
  assign tmp27211 = s1 ? tmp27212 : tmp24531;
  assign tmp27210 = s2 ? tmp27211 : tmp24532;
  assign tmp27209 = s3 ? tmp27210 : tmp24533;
  assign tmp27208 = s4 ? tmp24519 : tmp27209;
  assign tmp27217 = s0 ? tmp24498 : tmp26514;
  assign tmp27216 = s1 ? tmp27217 : tmp24514;
  assign tmp27215 = s2 ? tmp27216 : tmp24542;
  assign tmp27214 = s3 ? tmp27215 : tmp24545;
  assign tmp27221 = s0 ? tmp26514 : tmp24498;
  assign tmp27220 = s1 ? tmp27221 : tmp24526;
  assign tmp27219 = s2 ? tmp24536 : tmp27220;
  assign tmp27218 = s3 ? tmp27219 : tmp24553;
  assign tmp27213 = s4 ? tmp27214 : tmp27218;
  assign tmp27207 = s5 ? tmp27208 : tmp27213;
  assign tmp27206 = s6 ? tmp24495 : tmp27207;
  assign tmp27226 = s2 ? tmp27211 : tmp24498;
  assign tmp27225 = s3 ? tmp27226 : tmp24570;
  assign tmp27224 = s4 ? tmp24564 : tmp27225;
  assign tmp27229 = s2 ? tmp27216 : tmp24708;
  assign tmp27228 = s3 ? tmp27229 : tmp24576;
  assign tmp27227 = s4 ? tmp27228 : tmp24709;
  assign tmp27223 = s5 ? tmp27224 : tmp27227;
  assign tmp27222 = s6 ? tmp24556 : tmp27223;
  assign tmp27205 = s7 ? tmp27206 : tmp27222;
  assign tmp27204 = s8 ? tmp27205 : tmp27206;
  assign tmp27236 = s2 ? tmp24514 : tmp27067;
  assign tmp27235 = s3 ? tmp27236 : tmp24536;
  assign tmp27234 = s4 ? tmp27129 : tmp27235;
  assign tmp27233 = s5 ? tmp27119 : tmp27234;
  assign tmp27232 = s6 ? tmp27113 : tmp27233;
  assign tmp27243 = s0 ? tmp27143 : tmp24514;
  assign tmp27242 = s1 ? tmp27243 : tmp24514;
  assign tmp27241 = s2 ? tmp27242 : tmp24579;
  assign tmp27240 = s3 ? tmp26630 : tmp27241;
  assign tmp27239 = s4 ? tmp27240 : tmp24722;
  assign tmp27238 = s5 ? tmp27191 : tmp27239;
  assign tmp27237 = s6 ? tmp24683 : tmp27238;
  assign tmp27231 = s7 ? tmp27232 : tmp27237;
  assign tmp27246 = s5 ? tmp27158 : tmp27234;
  assign tmp27245 = s6 ? tmp27113 : tmp27246;
  assign tmp27249 = s4 ? tmp27228 : tmp24717;
  assign tmp27248 = s5 ? tmp27224 : tmp27249;
  assign tmp27247 = s6 ? tmp24556 : tmp27248;
  assign tmp27244 = s7 ? tmp27245 : tmp27247;
  assign tmp27230 = s8 ? tmp27231 : tmp27244;
  assign tmp27203 = s9 ? tmp27204 : tmp27230;
  assign tmp27059 = s10 ? tmp27060 : tmp27203;
  assign tmp27256 = s4 ? tmp27240 : tmp27200;
  assign tmp27255 = s5 ? tmp27191 : tmp27256;
  assign tmp27254 = s6 ? tmp24683 : tmp27255;
  assign tmp27253 = s7 ? tmp27112 : tmp27254;
  assign tmp27257 = s7 ? tmp27156 : tmp27222;
  assign tmp27252 = s8 ? tmp27253 : tmp27257;
  assign tmp27251 = s9 ? tmp27204 : tmp27252;
  assign tmp27250 = s10 ? tmp27060 : tmp27251;
  assign tmp27058 = s11 ? tmp27059 : tmp27250;
  assign tmp27057 = s12 ? tmp27058 : tmp24736;
  assign tmp27021 = s13 ? tmp27022 : tmp27057;
  assign tmp26987 = s14 ? tmp26988 : tmp27021;
  assign tmp27270 = s1 ? tmp26962 : tmp25553;
  assign tmp27269 = s2 ? tmp27270 : tmp25565;
  assign tmp27268 = s3 ? tmp27269 : tmp25566;
  assign tmp27267 = s4 ? tmp25676 : tmp27268;
  assign tmp27275 = s1 ? tmp26797 : tmp25679;
  assign tmp27274 = s2 ? tmp26794 : tmp27275;
  assign tmp27273 = s3 ? tmp27274 : tmp25685;
  assign tmp27278 = s1 ? tmp26801 : tmp26962;
  assign tmp27277 = s2 ? tmp26800 : tmp27278;
  assign tmp27276 = s3 ? tmp27277 : tmp25584;
  assign tmp27272 = s4 ? tmp27273 : tmp27276;
  assign tmp27271 = s5 ? tmp27272 : tmp25587;
  assign tmp27266 = s6 ? tmp27267 : tmp27271;
  assign tmp27281 = s3 ? tmp27269 : tmp25610;
  assign tmp27280 = s4 ? tmp25676 : tmp27281;
  assign tmp27285 = s2 ? tmp26794 : tmp25693;
  assign tmp27284 = s3 ? tmp27285 : tmp25617;
  assign tmp27283 = s4 ? tmp27284 : tmp26810;
  assign tmp27282 = s5 ? tmp27283 : tmp25694;
  assign tmp27279 = s6 ? tmp27280 : tmp27282;
  assign tmp27265 = s7 ? tmp27266 : tmp27279;
  assign tmp27264 = s8 ? tmp26893 : tmp27265;
  assign tmp27263 = s9 ? tmp26782 : tmp27264;
  assign tmp27290 = s5 ? tmp27283 : tmp25700;
  assign tmp27289 = s6 ? tmp27280 : tmp27290;
  assign tmp27288 = s7 ? tmp27266 : tmp27289;
  assign tmp27287 = s8 ? tmp27288 : tmp27266;
  assign tmp27292 = s7 ? tmp26971 : tmp27279;
  assign tmp27296 = s4 ? tmp26886 : tmp26980;
  assign tmp27295 = s5 ? tmp26919 : tmp27296;
  assign tmp27294 = s6 ? tmp26915 : tmp27295;
  assign tmp27293 = s7 ? tmp27294 : tmp27289;
  assign tmp27291 = s8 ? tmp27292 : tmp27293;
  assign tmp27286 = s9 ? tmp27287 : tmp27291;
  assign tmp27262 = s10 ? tmp27263 : tmp27286;
  assign tmp27300 = s7 ? tmp26803 : tmp27279;
  assign tmp27301 = s7 ? tmp26914 : tmp27289;
  assign tmp27299 = s8 ? tmp27300 : tmp27301;
  assign tmp27298 = s9 ? tmp27287 : tmp27299;
  assign tmp27297 = s10 ? tmp27263 : tmp27298;
  assign tmp27261 = s11 ? tmp27262 : tmp27297;
  assign tmp27260 = s12 ? tmp25269 : tmp27261;
  assign tmp27259 = s13 ? tmp27260 : tmp25712;
  assign tmp27258 = s14 ? tmp24859 : tmp27259;
  assign tmp26986 = s15 ? tmp26987 : tmp27258;
  assign tmp27315 = s1 ? tmp27067 : tmp27111;
  assign tmp27314 = s2 ? tmp26488 : tmp27315;
  assign tmp27313 = s3 ? tmp27074 : tmp27314;
  assign tmp27312 = s4 ? tmp27065 : tmp27313;
  assign tmp27320 = s1 ? tmp26563 : tmp27091;
  assign tmp27319 = s2 ? tmp27087 : tmp27320;
  assign tmp27318 = s3 ? tmp27085 : tmp27319;
  assign tmp27324 = s0 ? tmp23983 : tmp24536;
  assign tmp27323 = s1 ? tmp27091 : tmp27324;
  assign tmp27322 = s2 ? tmp27323 : tmp24514;
  assign tmp27321 = s3 ? tmp27093 : tmp27322;
  assign tmp27317 = s4 ? tmp27318 : tmp27321;
  assign tmp27328 = s1 ? tmp27104 : tmp26514;
  assign tmp27327 = s2 ? tmp27328 : tmp27107;
  assign tmp27326 = s3 ? tmp27327 : tmp24545;
  assign tmp27331 = s1 ? tmp24536 : tmp27143;
  assign tmp27330 = s2 ? tmp27331 : tmp27110;
  assign tmp27329 = s3 ? tmp27330 : tmp26575;
  assign tmp27325 = s4 ? tmp27326 : tmp27329;
  assign tmp27316 = s5 ? tmp27317 : tmp27325;
  assign tmp27311 = s6 ? tmp27312 : tmp27316;
  assign tmp27335 = s2 ? tmp26527 : tmp27315;
  assign tmp27334 = s3 ? tmp27115 : tmp27335;
  assign tmp27333 = s4 ? tmp27065 : tmp27334;
  assign tmp27339 = s2 ? tmp27067 : tmp27320;
  assign tmp27338 = s3 ? tmp27121 : tmp27339;
  assign tmp27337 = s4 ? tmp27338 : tmp27124;
  assign tmp27342 = s2 ? tmp27328 : tmp27131;
  assign tmp27341 = s3 ? tmp27342 : tmp24576;
  assign tmp27344 = s2 ? tmp26514 : tmp27134;
  assign tmp27343 = s3 ? tmp27344 : tmp24536;
  assign tmp27340 = s4 ? tmp27341 : tmp27343;
  assign tmp27336 = s5 ? tmp27337 : tmp27340;
  assign tmp27332 = s6 ? tmp27333 : tmp27336;
  assign tmp27310 = s7 ? tmp27311 : tmp27332;
  assign tmp27351 = s1 ? tmp26563 : tmp27142;
  assign tmp27350 = s2 ? tmp27087 : tmp27351;
  assign tmp27349 = s3 ? tmp27085 : tmp27350;
  assign tmp27354 = s1 ? tmp27142 : tmp26567;
  assign tmp27353 = s2 ? tmp27354 : tmp24514;
  assign tmp27352 = s3 ? tmp27145 : tmp27353;
  assign tmp27348 = s4 ? tmp27349 : tmp27352;
  assign tmp27358 = s1 ? tmp27111 : tmp27107;
  assign tmp27357 = s2 ? tmp27328 : tmp27358;
  assign tmp27356 = s3 ? tmp27357 : tmp24545;
  assign tmp27360 = s2 ? tmp26574 : tmp27110;
  assign tmp27359 = s3 ? tmp27360 : tmp26575;
  assign tmp27355 = s4 ? tmp27356 : tmp27359;
  assign tmp27347 = s5 ? tmp27348 : tmp27355;
  assign tmp27346 = s6 ? tmp27312 : tmp27347;
  assign tmp27365 = s2 ? tmp27067 : tmp27351;
  assign tmp27364 = s3 ? tmp27121 : tmp27365;
  assign tmp27363 = s4 ? tmp27364 : tmp27161;
  assign tmp27362 = s5 ? tmp27363 : tmp27340;
  assign tmp27361 = s6 ? tmp27333 : tmp27362;
  assign tmp27345 = s7 ? tmp27346 : tmp27361;
  assign tmp27309 = s8 ? tmp27310 : tmp27345;
  assign tmp27374 = s0 ? tmp27096 : tmp26472;
  assign tmp27373 = s1 ? tmp27374 : tmp26505;
  assign tmp27372 = s2 ? tmp27373 : tmp26506;
  assign tmp27371 = s3 ? tmp27372 : tmp26565;
  assign tmp27370 = s4 ? tmp26560 : tmp27371;
  assign tmp27379 = s0 ? tmp27143 : tmp26472;
  assign tmp27378 = s1 ? tmp26520 : tmp27379;
  assign tmp27377 = s2 ? tmp26571 : tmp27378;
  assign tmp27376 = s3 ? tmp27377 : tmp24545;
  assign tmp27383 = s0 ? tmp26472 : tmp27143;
  assign tmp27382 = s1 ? tmp26520 : tmp27383;
  assign tmp27381 = s2 ? tmp26574 : tmp27382;
  assign tmp27380 = s3 ? tmp27381 : tmp26575;
  assign tmp27375 = s4 ? tmp27376 : tmp27380;
  assign tmp27369 = s5 ? tmp27370 : tmp27375;
  assign tmp27368 = s6 ? tmp26595 : tmp27369;
  assign tmp27388 = s2 ? tmp27373 : tmp26472;
  assign tmp27387 = s3 ? tmp27388 : tmp26536;
  assign tmp27386 = s4 ? tmp26583 : tmp27387;
  assign tmp27392 = s1 ? tmp26472 : tmp27379;
  assign tmp27391 = s2 ? tmp26571 : tmp27392;
  assign tmp27390 = s3 ? tmp27391 : tmp27241;
  assign tmp27395 = s1 ? tmp26472 : tmp27383;
  assign tmp27394 = s2 ? tmp26514 : tmp27395;
  assign tmp27393 = s3 ? tmp27394 : tmp24536;
  assign tmp27389 = s4 ? tmp27390 : tmp27393;
  assign tmp27385 = s5 ? tmp27386 : tmp27389;
  assign tmp27384 = s6 ? tmp26605 : tmp27385;
  assign tmp27367 = s7 ? tmp27368 : tmp27384;
  assign tmp27366 = s8 ? tmp27345 : tmp27367;
  assign tmp27308 = s9 ? tmp27309 : tmp27366;
  assign tmp27397 = s8 ? tmp27345 : tmp27346;
  assign tmp27404 = s2 ? tmp26514 : tmp27067;
  assign tmp27403 = s3 ? tmp27404 : tmp24536;
  assign tmp27402 = s4 ? tmp27341 : tmp27403;
  assign tmp27401 = s5 ? tmp27337 : tmp27402;
  assign tmp27400 = s6 ? tmp27333 : tmp27401;
  assign tmp27407 = s4 ? tmp27390 : tmp26612;
  assign tmp27406 = s5 ? tmp27386 : tmp27407;
  assign tmp27405 = s6 ? tmp26605 : tmp27406;
  assign tmp27399 = s7 ? tmp27400 : tmp27405;
  assign tmp27409 = s5 ? tmp27363 : tmp27402;
  assign tmp27408 = s6 ? tmp27333 : tmp27409;
  assign tmp27398 = s8 ? tmp27399 : tmp27408;
  assign tmp27396 = s9 ? tmp27397 : tmp27398;
  assign tmp27307 = s10 ? tmp27308 : tmp27396;
  assign tmp27413 = s7 ? tmp27332 : tmp27384;
  assign tmp27412 = s8 ? tmp27413 : tmp27361;
  assign tmp27411 = s9 ? tmp27397 : tmp27412;
  assign tmp27410 = s10 ? tmp27308 : tmp27411;
  assign tmp27306 = s11 ? tmp27307 : tmp27410;
  assign tmp27305 = s12 ? tmp27306 : tmp24736;
  assign tmp27304 = s13 ? tmp26217 : tmp27305;
  assign tmp27303 = s14 ? tmp25951 : tmp27304;
  assign tmp27416 = s12 ? tmp25269 : tmp26779;
  assign tmp27415 = s13 ? tmp27416 : tmp25712;
  assign tmp27414 = s14 ? tmp24859 : tmp27415;
  assign tmp27302 = s15 ? tmp27303 : tmp27414;
  assign tmp26985 = s16 ? tmp26986 : tmp27302;
  assign tmp23951 = s17 ? tmp23952 : tmp26985;
  assign s11n = tmp23951;

  assign tmp27424 = ~(l4 ? 1 : 0);
  assign tmp27423 = l3 ? 1 : tmp27424;
  assign tmp27422 = l2 ? 1 : tmp27423;
  assign tmp27421 = l1 ? 1 : tmp27422;
  assign tmp27420 = s7 ? tmp27421 : 1;
  assign tmp27427 = l2 ? tmp27423 : 1;
  assign tmp27426 = l1 ? tmp27427 : tmp27423;
  assign tmp27425 = s7 ? tmp27426 : 1;
  assign tmp27419 = s8 ? tmp27420 : tmp27425;
  assign tmp27429 = s7 ? tmp27427 : 1;
  assign tmp27428 = s8 ? tmp27425 : tmp27429;
  assign tmp27418 = s9 ? tmp27419 : tmp27428;
  assign tmp27431 = s8 ? tmp27425 : tmp27426;
  assign tmp27430 = s9 ? tmp27431 : 1;
  assign tmp27417 = ~(s10 ? tmp27418 : tmp27430);
  assign s10n = tmp27417;

  assign tmp27439 = ~(l4 ? 1 : 0);
  assign tmp27438 = l3 ? 1 : tmp27439;
  assign tmp27437 = l2 ? 1 : tmp27438;
  assign tmp27436 = l1 ? 1 : tmp27437;
  assign tmp27440 = ~(l2 ? tmp27438 : 1);
  assign tmp27435 = s7 ? tmp27436 : tmp27440;
  assign tmp27441 = s7 ? tmp27436 : 0;
  assign tmp27434 = s8 ? tmp27435 : tmp27441;
  assign tmp27444 = ~(l1 ? 1 : tmp27437);
  assign tmp27443 = s7 ? 1 : tmp27444;
  assign tmp27442 = s8 ? tmp27441 : tmp27443;
  assign tmp27433 = s9 ? tmp27434 : tmp27442;
  assign tmp27449 = l2 ? tmp27438 : 1;
  assign tmp27448 = l1 ? tmp27449 : tmp27438;
  assign tmp27447 = s7 ? tmp27436 : tmp27448;
  assign tmp27446 = s8 ? tmp27441 : tmp27447;
  assign tmp27451 = s7 ? tmp27449 : tmp27436;
  assign tmp27450 = ~(s8 ? tmp27451 : 1);
  assign tmp27445 = s9 ? tmp27446 : tmp27450;
  assign tmp27432 = s10 ? tmp27433 : tmp27445;
  assign s9n = tmp27432;

  assign tmp27459 = ~(l4 ? 1 : 0);
  assign tmp27458 = l3 ? 1 : tmp27459;
  assign tmp27457 = l2 ? tmp27458 : 1;
  assign tmp27456 = l1 ? tmp27457 : tmp27458;
  assign tmp27461 = l2 ? 1 : tmp27458;
  assign tmp27460 = ~(l1 ? 1 : tmp27461);
  assign tmp27455 = s7 ? tmp27456 : tmp27460;
  assign tmp27463 = l1 ? 1 : tmp27461;
  assign tmp27464 = ~(l1 ? tmp27457 : tmp27458);
  assign tmp27462 = s7 ? tmp27463 : tmp27464;
  assign tmp27454 = s8 ? tmp27455 : tmp27462;
  assign tmp27466 = s7 ? tmp27456 : 0;
  assign tmp27465 = s8 ? tmp27462 : tmp27466;
  assign tmp27453 = s9 ? tmp27454 : tmp27465;
  assign tmp27469 = s7 ? tmp27456 : tmp27463;
  assign tmp27468 = s8 ? tmp27455 : tmp27469;
  assign tmp27471 = s7 ? tmp27463 : 1;
  assign tmp27470 = ~(s8 ? tmp27471 : tmp27469);
  assign tmp27467 = s9 ? tmp27468 : tmp27470;
  assign tmp27452 = s10 ? tmp27453 : tmp27467;
  assign s8n = tmp27452;

  assign tmp27488 = l4 ? 1 : 0;
  assign tmp27487 = ~(l3 ? tmp27488 : 1);
  assign tmp27486 = l2 ? 1 : tmp27487;
  assign tmp27490 = l3 ? 1 : 0;
  assign tmp27492 = ~(l4 ? 1 : 0);
  assign tmp27491 = ~(l3 ? 1 : tmp27492);
  assign tmp27489 = ~(l2 ? tmp27490 : tmp27491);
  assign tmp27485 = l1 ? tmp27486 : tmp27489;
  assign tmp27496 = l3 ? 1 : tmp27492;
  assign tmp27495 = l2 ? tmp27496 : 1;
  assign tmp27497 = l2 ? tmp27490 : 0;
  assign tmp27494 = l1 ? tmp27495 : tmp27497;
  assign tmp27499 = l2 ? 1 : tmp27492;
  assign tmp27498 = ~(l1 ? tmp27499 : tmp27489);
  assign tmp27493 = ~(s0 ? tmp27494 : tmp27498);
  assign tmp27484 = s1 ? tmp27485 : tmp27493;
  assign tmp27504 = l2 ? 1 : 0;
  assign tmp27506 = ~(l3 ? 1 : 0);
  assign tmp27505 = ~(l2 ? tmp27496 : tmp27506);
  assign tmp27503 = l1 ? tmp27504 : tmp27505;
  assign tmp27509 = l3 ? tmp27488 : 0;
  assign tmp27508 = l2 ? tmp27509 : tmp27488;
  assign tmp27510 = l2 ? tmp27509 : tmp27491;
  assign tmp27507 = ~(l1 ? tmp27508 : tmp27510);
  assign tmp27502 = s0 ? tmp27503 : tmp27507;
  assign tmp27513 = ~(l2 ? tmp27490 : tmp27506);
  assign tmp27512 = l1 ? tmp27486 : tmp27513;
  assign tmp27511 = s0 ? tmp27512 : tmp27507;
  assign tmp27501 = s1 ? tmp27502 : tmp27511;
  assign tmp27517 = l2 ? tmp27496 : 0;
  assign tmp27516 = ~(l1 ? tmp27495 : tmp27517);
  assign tmp27515 = s0 ? tmp27512 : tmp27516;
  assign tmp27519 = l1 ? tmp27508 : tmp27510;
  assign tmp27521 = l2 ? tmp27490 : tmp27491;
  assign tmp27520 = l1 ? tmp27508 : tmp27521;
  assign tmp27518 = ~(s0 ? tmp27519 : tmp27520);
  assign tmp27514 = s1 ? tmp27515 : tmp27518;
  assign tmp27500 = s2 ? tmp27501 : tmp27514;
  assign tmp27483 = s3 ? tmp27484 : tmp27500;
  assign tmp27526 = l1 ? tmp27504 : tmp27489;
  assign tmp27525 = s0 ? tmp27526 : tmp27516;
  assign tmp27527 = ~(s0 ? tmp27520 : tmp27519);
  assign tmp27524 = s1 ? tmp27525 : tmp27527;
  assign tmp27530 = ~(l1 ? tmp27495 : 0);
  assign tmp27529 = s0 ? tmp27485 : tmp27530;
  assign tmp27532 = l1 ? tmp27495 : tmp27490;
  assign tmp27533 = l1 ? tmp27495 : 0;
  assign tmp27531 = ~(s0 ? tmp27532 : tmp27533);
  assign tmp27528 = s1 ? tmp27529 : tmp27531;
  assign tmp27523 = s2 ? tmp27524 : tmp27528;
  assign tmp27536 = s0 ? tmp27532 : tmp27494;
  assign tmp27537 = s0 ? tmp27533 : 0;
  assign tmp27535 = s1 ? tmp27536 : tmp27537;
  assign tmp27539 = ~(s0 ? 1 : tmp27507);
  assign tmp27538 = s1 ? tmp27519 : tmp27539;
  assign tmp27534 = ~(s2 ? tmp27535 : tmp27538);
  assign tmp27522 = s3 ? tmp27523 : tmp27534;
  assign tmp27482 = s4 ? tmp27483 : tmp27522;
  assign tmp27546 = l1 ? tmp27499 : tmp27489;
  assign tmp27545 = s0 ? tmp27546 : tmp27516;
  assign tmp27548 = l1 ? tmp27495 : tmp27517;
  assign tmp27549 = ~(l1 ? tmp27504 : tmp27505);
  assign tmp27547 = ~(s0 ? tmp27548 : tmp27549);
  assign tmp27544 = s1 ? tmp27545 : tmp27547;
  assign tmp27554 = l3 ? 1 : tmp27488;
  assign tmp27553 = ~(l2 ? tmp27490 : tmp27554);
  assign tmp27552 = ~(l1 ? tmp27499 : tmp27553);
  assign tmp27551 = s0 ? tmp27548 : tmp27552;
  assign tmp27555 = s0 ? tmp27519 : tmp27517;
  assign tmp27550 = ~(s1 ? tmp27551 : tmp27555);
  assign tmp27543 = s2 ? tmp27544 : tmp27550;
  assign tmp27560 = l2 ? 1 : tmp27490;
  assign tmp27559 = ~(l1 ? tmp27560 : tmp27513);
  assign tmp27558 = s0 ? tmp27517 : tmp27559;
  assign tmp27561 = s0 ? tmp27517 : tmp27508;
  assign tmp27557 = s1 ? tmp27558 : tmp27561;
  assign tmp27563 = ~(l2 ? tmp27509 : tmp27488);
  assign tmp27562 = ~(s1 ? 1 : tmp27563);
  assign tmp27556 = ~(s2 ? tmp27557 : tmp27562);
  assign tmp27542 = s3 ? tmp27543 : tmp27556;
  assign tmp27569 = l2 ? tmp27490 : tmp27488;
  assign tmp27568 = ~(l1 ? tmp27508 : tmp27569);
  assign tmp27567 = s0 ? 1 : tmp27568;
  assign tmp27570 = ~(s0 ? tmp27495 : tmp27533);
  assign tmp27566 = s1 ? tmp27567 : tmp27570;
  assign tmp27572 = s0 ? tmp27495 : tmp27533;
  assign tmp27574 = l1 ? tmp27504 : tmp27553;
  assign tmp27575 = ~(l2 ? tmp27496 : 1);
  assign tmp27573 = ~(s0 ? tmp27574 : tmp27575);
  assign tmp27571 = ~(s1 ? tmp27572 : tmp27573);
  assign tmp27565 = s2 ? tmp27566 : tmp27571;
  assign tmp27579 = l1 ? tmp27560 : tmp27499;
  assign tmp27578 = s0 ? tmp27574 : tmp27579;
  assign tmp27580 = ~(s0 ? tmp27533 : tmp27508);
  assign tmp27577 = s1 ? tmp27578 : tmp27580;
  assign tmp27576 = s2 ? tmp27577 : 1;
  assign tmp27564 = s3 ? tmp27565 : tmp27576;
  assign tmp27541 = s4 ? tmp27542 : tmp27564;
  assign tmp27585 = s0 ? tmp27508 : 0;
  assign tmp27584 = s1 ? tmp27585 : 0;
  assign tmp27588 = l1 ? tmp27504 : tmp27575;
  assign tmp27587 = s0 ? 1 : tmp27588;
  assign tmp27586 = ~(s1 ? tmp27587 : tmp27588);
  assign tmp27583 = s2 ? tmp27584 : tmp27586;
  assign tmp27591 = s0 ? tmp27588 : 1;
  assign tmp27590 = s1 ? tmp27591 : 1;
  assign tmp27594 = l1 ? tmp27504 : tmp27563;
  assign tmp27593 = s0 ? 1 : tmp27594;
  assign tmp27592 = s1 ? 1 : tmp27593;
  assign tmp27589 = ~(s2 ? tmp27590 : tmp27592);
  assign tmp27582 = s3 ? tmp27583 : tmp27589;
  assign tmp27598 = s0 ? tmp27594 : 1;
  assign tmp27597 = s1 ? tmp27598 : 1;
  assign tmp27601 = l1 ? tmp27499 : tmp27553;
  assign tmp27600 = s0 ? 1 : tmp27601;
  assign tmp27599 = s1 ? tmp27600 : tmp27588;
  assign tmp27596 = s2 ? tmp27597 : tmp27599;
  assign tmp27606 = ~(l2 ? 1 : tmp27492);
  assign tmp27605 = ~(l1 ? tmp27508 : tmp27606);
  assign tmp27604 = s0 ? 1 : tmp27605;
  assign tmp27603 = s1 ? 1 : tmp27604;
  assign tmp27607 = s1 ? tmp27593 : 1;
  assign tmp27602 = s2 ? tmp27603 : tmp27607;
  assign tmp27595 = ~(s3 ? tmp27596 : tmp27602);
  assign tmp27581 = ~(s4 ? tmp27582 : tmp27595);
  assign tmp27540 = s5 ? tmp27541 : tmp27581;
  assign tmp27481 = s6 ? tmp27482 : tmp27540;
  assign tmp27480 = s7 ? tmp27481 : tmp27575;
  assign tmp27615 = l3 ? tmp27488 : 1;
  assign tmp27614 = l2 ? tmp27488 : tmp27615;
  assign tmp27613 = l1 ? tmp27614 : tmp27521;
  assign tmp27617 = l1 ? 1 : tmp27497;
  assign tmp27618 = l1 ? tmp27488 : tmp27521;
  assign tmp27616 = s0 ? tmp27617 : tmp27618;
  assign tmp27612 = s1 ? tmp27613 : tmp27616;
  assign tmp27623 = l2 ? tmp27488 : 1;
  assign tmp27624 = l2 ? tmp27490 : tmp27506;
  assign tmp27622 = l1 ? tmp27623 : tmp27624;
  assign tmp27625 = l1 ? tmp27488 : tmp27510;
  assign tmp27621 = s0 ? tmp27622 : tmp27625;
  assign tmp27627 = l1 ? tmp27614 : tmp27624;
  assign tmp27626 = s0 ? tmp27627 : tmp27625;
  assign tmp27620 = s1 ? tmp27621 : tmp27626;
  assign tmp27629 = s0 ? tmp27627 : tmp27617;
  assign tmp27630 = s0 ? tmp27625 : tmp27618;
  assign tmp27628 = s1 ? tmp27629 : tmp27630;
  assign tmp27619 = s2 ? tmp27620 : tmp27628;
  assign tmp27611 = s3 ? tmp27612 : tmp27619;
  assign tmp27635 = l1 ? tmp27623 : tmp27521;
  assign tmp27636 = l1 ? 1 : tmp27504;
  assign tmp27634 = s0 ? tmp27635 : tmp27636;
  assign tmp27637 = s0 ? tmp27618 : tmp27625;
  assign tmp27633 = s1 ? tmp27634 : tmp27637;
  assign tmp27640 = l1 ? 1 : 0;
  assign tmp27639 = s0 ? tmp27613 : tmp27640;
  assign tmp27642 = l1 ? 1 : tmp27490;
  assign tmp27641 = s0 ? tmp27642 : tmp27640;
  assign tmp27638 = s1 ? tmp27639 : tmp27641;
  assign tmp27632 = s2 ? tmp27633 : tmp27638;
  assign tmp27645 = s0 ? tmp27642 : tmp27617;
  assign tmp27646 = s0 ? tmp27640 : 0;
  assign tmp27644 = s1 ? tmp27645 : tmp27646;
  assign tmp27649 = ~(l1 ? tmp27488 : tmp27510);
  assign tmp27648 = ~(s0 ? 1 : tmp27649);
  assign tmp27647 = s1 ? tmp27625 : tmp27648;
  assign tmp27643 = s2 ? tmp27644 : tmp27647;
  assign tmp27631 = s3 ? tmp27632 : tmp27643;
  assign tmp27610 = s4 ? tmp27611 : tmp27631;
  assign tmp27655 = s0 ? tmp27618 : tmp27636;
  assign tmp27656 = s0 ? tmp27636 : tmp27622;
  assign tmp27654 = s1 ? tmp27655 : tmp27656;
  assign tmp27659 = l1 ? tmp27488 : tmp27569;
  assign tmp27658 = s0 ? tmp27636 : tmp27659;
  assign tmp27660 = s0 ? tmp27625 : tmp27617;
  assign tmp27657 = s1 ? tmp27658 : tmp27660;
  assign tmp27653 = s2 ? tmp27654 : tmp27657;
  assign tmp27665 = l2 ? tmp27488 : tmp27506;
  assign tmp27664 = l1 ? tmp27665 : tmp27624;
  assign tmp27663 = s0 ? tmp27617 : tmp27664;
  assign tmp27667 = l1 ? tmp27488 : tmp27508;
  assign tmp27666 = s0 ? tmp27617 : tmp27667;
  assign tmp27662 = s1 ? tmp27663 : tmp27666;
  assign tmp27669 = ~(l1 ? tmp27488 : tmp27508);
  assign tmp27668 = ~(s1 ? 1 : tmp27669);
  assign tmp27661 = s2 ? tmp27662 : tmp27668;
  assign tmp27652 = s3 ? tmp27653 : tmp27661;
  assign tmp27674 = ~(l1 ? tmp27488 : tmp27569);
  assign tmp27673 = s0 ? 1 : tmp27674;
  assign tmp27675 = ~(s0 ? 1 : tmp27640);
  assign tmp27672 = s1 ? tmp27673 : tmp27675;
  assign tmp27677 = s0 ? 1 : tmp27640;
  assign tmp27679 = l1 ? tmp27623 : tmp27569;
  assign tmp27678 = s0 ? tmp27679 : 1;
  assign tmp27676 = ~(s1 ? tmp27677 : tmp27678);
  assign tmp27671 = s2 ? tmp27672 : tmp27676;
  assign tmp27684 = ~(l2 ? tmp27490 : tmp27488);
  assign tmp27683 = l1 ? tmp27504 : tmp27684;
  assign tmp27685 = ~(l1 ? tmp27665 : tmp27606);
  assign tmp27682 = s0 ? tmp27683 : tmp27685;
  assign tmp27686 = ~(s0 ? tmp27640 : tmp27488);
  assign tmp27681 = s1 ? tmp27682 : tmp27686;
  assign tmp27680 = s2 ? tmp27681 : 1;
  assign tmp27670 = ~(s3 ? tmp27671 : tmp27680);
  assign tmp27651 = s4 ? tmp27652 : tmp27670;
  assign tmp27691 = s0 ? tmp27667 : 0;
  assign tmp27690 = s1 ? tmp27691 : 0;
  assign tmp27695 = ~(l2 ? tmp27490 : 1);
  assign tmp27694 = l1 ? tmp27504 : tmp27695;
  assign tmp27693 = s0 ? 1 : tmp27694;
  assign tmp27697 = l1 ? tmp27504 : 0;
  assign tmp27696 = s0 ? tmp27697 : tmp27694;
  assign tmp27692 = ~(s1 ? tmp27693 : tmp27696);
  assign tmp27689 = s2 ? tmp27690 : tmp27692;
  assign tmp27700 = s0 ? tmp27697 : 1;
  assign tmp27699 = s1 ? tmp27700 : 1;
  assign tmp27703 = l1 ? tmp27504 : tmp27492;
  assign tmp27702 = s0 ? 1 : tmp27703;
  assign tmp27701 = s1 ? 1 : tmp27702;
  assign tmp27698 = ~(s2 ? tmp27699 : tmp27701);
  assign tmp27688 = s3 ? tmp27689 : tmp27698;
  assign tmp27707 = s0 ? tmp27703 : 1;
  assign tmp27706 = s1 ? tmp27707 : 1;
  assign tmp27710 = l1 ? tmp27499 : tmp27684;
  assign tmp27709 = s0 ? 1 : tmp27710;
  assign tmp27711 = s0 ? tmp27694 : tmp27697;
  assign tmp27708 = s1 ? tmp27709 : tmp27711;
  assign tmp27705 = s2 ? tmp27706 : tmp27708;
  assign tmp27715 = ~(l1 ? tmp27488 : tmp27606);
  assign tmp27714 = s0 ? 1 : tmp27715;
  assign tmp27713 = s1 ? 1 : tmp27714;
  assign tmp27716 = s1 ? tmp27702 : 1;
  assign tmp27712 = s2 ? tmp27713 : tmp27716;
  assign tmp27704 = ~(s3 ? tmp27705 : tmp27712);
  assign tmp27687 = s4 ? tmp27688 : tmp27704;
  assign tmp27650 = s5 ? tmp27651 : tmp27687;
  assign tmp27609 = s6 ? tmp27610 : tmp27650;
  assign tmp27608 = ~(s7 ? tmp27609 : tmp27495);
  assign tmp27479 = s8 ? tmp27480 : tmp27608;
  assign tmp27718 = s7 ? tmp27609 : tmp27495;
  assign tmp27724 = s0 ? tmp27526 : tmp27546;
  assign tmp27723 = s1 ? tmp27485 : tmp27724;
  assign tmp27729 = ~(l2 ? tmp27509 : tmp27491);
  assign tmp27728 = l1 ? tmp27499 : tmp27729;
  assign tmp27727 = s0 ? tmp27526 : tmp27728;
  assign tmp27730 = s0 ? tmp27485 : tmp27728;
  assign tmp27726 = s1 ? tmp27727 : tmp27730;
  assign tmp27732 = s0 ? tmp27485 : tmp27526;
  assign tmp27733 = s0 ? tmp27728 : tmp27546;
  assign tmp27731 = s1 ? tmp27732 : tmp27733;
  assign tmp27725 = s2 ? tmp27726 : tmp27731;
  assign tmp27722 = s3 ? tmp27723 : tmp27725;
  assign tmp27739 = ~(l2 ? 1 : tmp27491);
  assign tmp27738 = l1 ? tmp27504 : tmp27739;
  assign tmp27737 = s0 ? tmp27526 : tmp27738;
  assign tmp27740 = s0 ? tmp27546 : tmp27728;
  assign tmp27736 = s1 ? tmp27737 : tmp27740;
  assign tmp27744 = l2 ? 1 : tmp27496;
  assign tmp27743 = l1 ? tmp27504 : tmp27744;
  assign tmp27742 = s0 ? tmp27485 : tmp27743;
  assign tmp27745 = s0 ? tmp27574 : tmp27743;
  assign tmp27741 = s1 ? tmp27742 : tmp27745;
  assign tmp27735 = s2 ? tmp27736 : tmp27741;
  assign tmp27748 = s0 ? tmp27574 : tmp27526;
  assign tmp27750 = l1 ? 1 : tmp27744;
  assign tmp27749 = s0 ? tmp27743 : tmp27750;
  assign tmp27747 = s1 ? tmp27748 : tmp27749;
  assign tmp27752 = s0 ? tmp27750 : tmp27728;
  assign tmp27751 = s1 ? tmp27728 : tmp27752;
  assign tmp27746 = s2 ? tmp27747 : tmp27751;
  assign tmp27734 = s3 ? tmp27735 : tmp27746;
  assign tmp27721 = s4 ? tmp27722 : tmp27734;
  assign tmp27760 = l2 ? 1 : tmp27491;
  assign tmp27759 = ~(l1 ? 1 : tmp27760);
  assign tmp27758 = s0 ? tmp27546 : tmp27759;
  assign tmp27762 = l1 ? 1 : tmp27760;
  assign tmp27763 = ~(l1 ? tmp27504 : tmp27489);
  assign tmp27761 = ~(s0 ? tmp27762 : tmp27763);
  assign tmp27757 = s1 ? tmp27758 : tmp27761;
  assign tmp27765 = s0 ? tmp27762 : tmp27498;
  assign tmp27767 = l1 ? 1 : tmp27489;
  assign tmp27766 = ~(s0 ? tmp27728 : tmp27767);
  assign tmp27764 = ~(s1 ? tmp27765 : tmp27766);
  assign tmp27756 = s2 ? tmp27757 : tmp27764;
  assign tmp27771 = l1 ? tmp27560 : tmp27489;
  assign tmp27770 = s0 ? tmp27767 : tmp27771;
  assign tmp27772 = s0 ? tmp27767 : tmp27649;
  assign tmp27769 = s1 ? tmp27770 : tmp27772;
  assign tmp27773 = s1 ? tmp27750 : tmp27563;
  assign tmp27768 = s2 ? tmp27769 : tmp27773;
  assign tmp27755 = s3 ? tmp27756 : tmp27768;
  assign tmp27777 = s0 ? tmp27750 : tmp27546;
  assign tmp27778 = s0 ? tmp27697 : tmp27743;
  assign tmp27776 = s1 ? tmp27777 : tmp27778;
  assign tmp27780 = s0 ? tmp27526 : tmp27697;
  assign tmp27779 = s1 ? tmp27778 : tmp27780;
  assign tmp27775 = s2 ? tmp27776 : tmp27779;
  assign tmp27784 = l1 ? tmp27560 : tmp27744;
  assign tmp27783 = s0 ? tmp27526 : tmp27784;
  assign tmp27785 = s0 ? tmp27743 : tmp27492;
  assign tmp27782 = s1 ? tmp27783 : tmp27785;
  assign tmp27781 = s2 ? tmp27782 : tmp27750;
  assign tmp27774 = s3 ? tmp27775 : tmp27781;
  assign tmp27754 = s4 ? tmp27755 : tmp27774;
  assign tmp27791 = ~(l1 ? 1 : tmp27744);
  assign tmp27790 = s0 ? tmp27625 : tmp27791;
  assign tmp27789 = s1 ? tmp27790 : tmp27791;
  assign tmp27793 = s0 ? tmp27750 : tmp27574;
  assign tmp27794 = s0 ? tmp27504 : tmp27574;
  assign tmp27792 = ~(s1 ? tmp27793 : tmp27794);
  assign tmp27788 = s2 ? tmp27789 : tmp27792;
  assign tmp27797 = s0 ? tmp27504 : tmp27750;
  assign tmp27796 = s1 ? tmp27797 : tmp27750;
  assign tmp27799 = s0 ? tmp27750 : tmp27743;
  assign tmp27798 = s1 ? tmp27750 : tmp27799;
  assign tmp27795 = ~(s2 ? tmp27796 : tmp27798);
  assign tmp27787 = s3 ? tmp27788 : tmp27795;
  assign tmp27802 = s1 ? tmp27749 : tmp27750;
  assign tmp27804 = s0 ? tmp27574 : tmp27504;
  assign tmp27803 = s1 ? tmp27777 : tmp27804;
  assign tmp27801 = s2 ? tmp27802 : tmp27803;
  assign tmp27809 = ~(l2 ? 1 : tmp27496);
  assign tmp27808 = ~(l1 ? tmp27488 : tmp27809);
  assign tmp27807 = s0 ? tmp27750 : tmp27808;
  assign tmp27806 = s1 ? tmp27750 : tmp27807;
  assign tmp27810 = s1 ? tmp27799 : tmp27750;
  assign tmp27805 = s2 ? tmp27806 : tmp27810;
  assign tmp27800 = ~(s3 ? tmp27801 : tmp27805);
  assign tmp27786 = ~(s4 ? tmp27787 : tmp27800);
  assign tmp27753 = s5 ? tmp27754 : tmp27786;
  assign tmp27720 = s6 ? tmp27721 : tmp27753;
  assign tmp27719 = ~(s7 ? tmp27720 : tmp27575);
  assign tmp27717 = ~(s8 ? tmp27718 : tmp27719);
  assign tmp27478 = s9 ? tmp27479 : tmp27717;
  assign tmp27820 = ~(l2 ? tmp27490 : 0);
  assign tmp27819 = l1 ? tmp27504 : tmp27820;
  assign tmp27818 = s0 ? tmp27819 : tmp27546;
  assign tmp27817 = s1 ? tmp27485 : tmp27818;
  assign tmp27824 = l1 ? tmp27504 : tmp27513;
  assign tmp27823 = s0 ? tmp27824 : tmp27728;
  assign tmp27825 = s0 ? tmp27512 : tmp27728;
  assign tmp27822 = s1 ? tmp27823 : tmp27825;
  assign tmp27827 = s0 ? tmp27512 : tmp27819;
  assign tmp27826 = s1 ? tmp27827 : tmp27733;
  assign tmp27821 = s2 ? tmp27822 : tmp27826;
  assign tmp27816 = s3 ? tmp27817 : tmp27821;
  assign tmp27833 = ~(l2 ? 1 : 0);
  assign tmp27832 = l1 ? tmp27504 : tmp27833;
  assign tmp27831 = s0 ? tmp27526 : tmp27832;
  assign tmp27830 = s1 ? tmp27831 : tmp27740;
  assign tmp27836 = l1 ? tmp27504 : 1;
  assign tmp27835 = s0 ? tmp27485 : tmp27836;
  assign tmp27838 = l1 ? tmp27504 : tmp27506;
  assign tmp27837 = s0 ? tmp27838 : tmp27836;
  assign tmp27834 = s1 ? tmp27835 : tmp27837;
  assign tmp27829 = s2 ? tmp27830 : tmp27834;
  assign tmp27841 = s0 ? tmp27838 : tmp27819;
  assign tmp27842 = s0 ? tmp27836 : 1;
  assign tmp27840 = s1 ? tmp27841 : tmp27842;
  assign tmp27844 = s0 ? 1 : tmp27728;
  assign tmp27843 = s1 ? tmp27728 : tmp27844;
  assign tmp27839 = s2 ? tmp27840 : tmp27843;
  assign tmp27828 = s3 ? tmp27829 : tmp27839;
  assign tmp27815 = s4 ? tmp27816 : tmp27828;
  assign tmp27851 = ~(l1 ? 1 : tmp27504);
  assign tmp27850 = s0 ? tmp27546 : tmp27851;
  assign tmp27853 = ~(l1 ? tmp27504 : tmp27513);
  assign tmp27852 = ~(s0 ? tmp27636 : tmp27853);
  assign tmp27849 = s1 ? tmp27850 : tmp27852;
  assign tmp27856 = ~(l1 ? tmp27499 : tmp27684);
  assign tmp27855 = s0 ? tmp27636 : tmp27856;
  assign tmp27858 = l1 ? 1 : tmp27820;
  assign tmp27857 = ~(s0 ? tmp27728 : tmp27858);
  assign tmp27854 = ~(s1 ? tmp27855 : tmp27857);
  assign tmp27848 = s2 ? tmp27849 : tmp27854;
  assign tmp27862 = l1 ? tmp27560 : tmp27513;
  assign tmp27861 = s0 ? tmp27858 : tmp27862;
  assign tmp27863 = s0 ? tmp27858 : tmp27669;
  assign tmp27860 = s1 ? tmp27861 : tmp27863;
  assign tmp27864 = s1 ? 1 : tmp27563;
  assign tmp27859 = s2 ? tmp27860 : tmp27864;
  assign tmp27847 = s3 ? tmp27848 : tmp27859;
  assign tmp27868 = s0 ? tmp27697 : tmp27836;
  assign tmp27867 = s1 ? tmp27709 : tmp27868;
  assign tmp27870 = s0 ? tmp27683 : tmp27697;
  assign tmp27869 = s1 ? tmp27868 : tmp27870;
  assign tmp27866 = s2 ? tmp27867 : tmp27869;
  assign tmp27873 = s0 ? tmp27683 : tmp27579;
  assign tmp27874 = s0 ? tmp27836 : tmp27492;
  assign tmp27872 = s1 ? tmp27873 : tmp27874;
  assign tmp27871 = s2 ? tmp27872 : 1;
  assign tmp27865 = s3 ? tmp27866 : tmp27871;
  assign tmp27846 = s4 ? tmp27847 : tmp27865;
  assign tmp27875 = ~(s4 ? tmp27688 : tmp27704);
  assign tmp27845 = s5 ? tmp27846 : tmp27875;
  assign tmp27814 = s6 ? tmp27815 : tmp27845;
  assign tmp27813 = s7 ? tmp27814 : tmp27575;
  assign tmp27812 = s8 ? tmp27813 : tmp27814;
  assign tmp27811 = s9 ? tmp27812 : tmp27575;
  assign tmp27477 = s10 ? tmp27478 : tmp27811;
  assign tmp27887 = ~(l3 ? tmp27488 : 0);
  assign tmp27886 = l2 ? 1 : tmp27887;
  assign tmp27888 = ~(l2 ? tmp27490 : tmp27509);
  assign tmp27885 = l1 ? tmp27886 : tmp27888;
  assign tmp27891 = l2 ? tmp27490 : 1;
  assign tmp27890 = l1 ? tmp27490 : tmp27891;
  assign tmp27892 = ~(l1 ? tmp27886 : tmp27506);
  assign tmp27889 = ~(s0 ? tmp27890 : tmp27892);
  assign tmp27884 = s1 ? tmp27885 : tmp27889;
  assign tmp27897 = l2 ? 1 : tmp27506;
  assign tmp27898 = ~(l2 ? tmp27496 : tmp27490);
  assign tmp27896 = l1 ? tmp27897 : tmp27898;
  assign tmp27895 = s0 ? tmp27896 : tmp27887;
  assign tmp27900 = l1 ? tmp27886 : tmp27506;
  assign tmp27899 = s0 ? tmp27900 : tmp27887;
  assign tmp27894 = s1 ? tmp27895 : tmp27899;
  assign tmp27902 = s0 ? tmp27900 : tmp27575;
  assign tmp27904 = ~(l1 ? tmp27886 : tmp27888);
  assign tmp27903 = ~(s0 ? tmp27509 : tmp27904);
  assign tmp27901 = s1 ? tmp27902 : tmp27903;
  assign tmp27893 = s2 ? tmp27894 : tmp27901;
  assign tmp27883 = s3 ? tmp27884 : tmp27893;
  assign tmp27909 = l1 ? tmp27897 : tmp27506;
  assign tmp27910 = ~(l1 ? tmp27490 : tmp27495);
  assign tmp27908 = s0 ? tmp27909 : tmp27910;
  assign tmp27911 = s0 ? tmp27885 : tmp27887;
  assign tmp27907 = s1 ? tmp27908 : tmp27911;
  assign tmp27913 = s0 ? tmp27885 : tmp27575;
  assign tmp27914 = ~(s0 ? tmp27490 : tmp27495);
  assign tmp27912 = s1 ? tmp27913 : tmp27914;
  assign tmp27906 = s2 ? tmp27907 : tmp27912;
  assign tmp27917 = s0 ? tmp27495 : 0;
  assign tmp27916 = s1 ? tmp27890 : tmp27917;
  assign tmp27919 = ~(s0 ? 1 : tmp27887);
  assign tmp27918 = s1 ? tmp27509 : tmp27919;
  assign tmp27915 = ~(s2 ? tmp27916 : tmp27918);
  assign tmp27905 = s3 ? tmp27906 : tmp27915;
  assign tmp27882 = s4 ? tmp27883 : tmp27905;
  assign tmp27926 = ~(l1 ? tmp27897 : tmp27898);
  assign tmp27925 = ~(s0 ? tmp27495 : tmp27926);
  assign tmp27924 = s1 ? tmp27902 : tmp27925;
  assign tmp27929 = ~(l1 ? tmp27886 : tmp27820);
  assign tmp27928 = s0 ? tmp27495 : tmp27929;
  assign tmp27930 = s0 ? tmp27509 : tmp27495;
  assign tmp27927 = ~(s1 ? tmp27928 : tmp27930);
  assign tmp27923 = s2 ? tmp27924 : tmp27927;
  assign tmp27934 = ~(l1 ? 1 : tmp27506);
  assign tmp27933 = s0 ? tmp27495 : tmp27934;
  assign tmp27936 = l2 ? tmp27509 : 0;
  assign tmp27935 = s0 ? tmp27495 : tmp27936;
  assign tmp27932 = s1 ? tmp27933 : tmp27935;
  assign tmp27937 = ~(s1 ? 1 : tmp27887);
  assign tmp27931 = ~(s2 ? tmp27932 : tmp27937);
  assign tmp27922 = s3 ? tmp27923 : tmp27931;
  assign tmp27942 = l1 ? tmp27886 : tmp27820;
  assign tmp27941 = s0 ? 1 : tmp27942;
  assign tmp27944 = l1 ? tmp27490 : tmp27495;
  assign tmp27943 = ~(s0 ? tmp27944 : 0);
  assign tmp27940 = s1 ? tmp27941 : tmp27943;
  assign tmp27946 = s0 ? tmp27944 : 0;
  assign tmp27948 = l1 ? tmp27897 : tmp27820;
  assign tmp27947 = ~(s0 ? tmp27948 : tmp27910);
  assign tmp27945 = ~(s1 ? tmp27946 : tmp27947);
  assign tmp27939 = s2 ? tmp27940 : tmp27945;
  assign tmp27951 = s0 ? tmp27858 : 1;
  assign tmp27950 = s1 ? tmp27951 : 1;
  assign tmp27949 = s2 ? tmp27950 : 1;
  assign tmp27938 = s3 ? tmp27939 : tmp27949;
  assign tmp27921 = s4 ? tmp27922 : tmp27938;
  assign tmp27956 = s0 ? tmp27936 : 0;
  assign tmp27955 = s1 ? tmp27956 : 0;
  assign tmp27960 = ~(l2 ? tmp27496 : 0);
  assign tmp27959 = l1 ? 1 : tmp27960;
  assign tmp27958 = s0 ? 1 : tmp27959;
  assign tmp27957 = ~(s1 ? tmp27958 : tmp27959);
  assign tmp27954 = s2 ? tmp27955 : tmp27957;
  assign tmp27953 = s3 ? tmp27954 : 0;
  assign tmp27964 = s0 ? 1 : tmp27858;
  assign tmp27963 = s1 ? tmp27964 : tmp27959;
  assign tmp27962 = s2 ? 1 : tmp27963;
  assign tmp27961 = ~(s3 ? tmp27962 : 1);
  assign tmp27952 = ~(s4 ? tmp27953 : tmp27961);
  assign tmp27920 = s5 ? tmp27921 : tmp27952;
  assign tmp27881 = s6 ? tmp27882 : tmp27920;
  assign tmp27880 = s7 ? tmp27881 : tmp27575;
  assign tmp27971 = l2 ? tmp27488 : tmp27509;
  assign tmp27972 = l2 ? tmp27490 : tmp27509;
  assign tmp27970 = l1 ? tmp27971 : tmp27972;
  assign tmp27974 = l1 ? tmp27560 : tmp27891;
  assign tmp27975 = l1 ? tmp27971 : tmp27490;
  assign tmp27973 = s0 ? tmp27974 : tmp27975;
  assign tmp27969 = s1 ? tmp27970 : tmp27973;
  assign tmp27980 = l2 ? tmp27488 : tmp27490;
  assign tmp27979 = l1 ? tmp27980 : tmp27490;
  assign tmp27981 = l1 ? tmp27971 : tmp27509;
  assign tmp27978 = s0 ? tmp27979 : tmp27981;
  assign tmp27982 = s0 ? tmp27975 : tmp27981;
  assign tmp27977 = s1 ? tmp27978 : tmp27982;
  assign tmp27985 = l1 ? 1 : tmp27891;
  assign tmp27984 = s0 ? tmp27975 : tmp27985;
  assign tmp27986 = s0 ? tmp27981 : tmp27970;
  assign tmp27983 = s1 ? tmp27984 : tmp27986;
  assign tmp27976 = s2 ? tmp27977 : tmp27983;
  assign tmp27968 = s3 ? tmp27969 : tmp27976;
  assign tmp27991 = l1 ? tmp27560 : 1;
  assign tmp27990 = s0 ? tmp27979 : tmp27991;
  assign tmp27992 = s0 ? tmp27970 : tmp27981;
  assign tmp27989 = s1 ? tmp27990 : tmp27992;
  assign tmp27994 = s0 ? tmp27970 : 1;
  assign tmp27996 = l1 ? tmp27560 : tmp27490;
  assign tmp27995 = s0 ? tmp27996 : 1;
  assign tmp27993 = s1 ? tmp27994 : tmp27995;
  assign tmp27988 = s2 ? tmp27989 : tmp27993;
  assign tmp27999 = s0 ? 1 : 0;
  assign tmp27998 = s1 ? tmp27974 : tmp27999;
  assign tmp28002 = ~(l1 ? tmp27971 : tmp27509);
  assign tmp28001 = ~(s0 ? 1 : tmp28002);
  assign tmp28000 = s1 ? tmp27981 : tmp28001;
  assign tmp27997 = s2 ? tmp27998 : tmp28000;
  assign tmp27987 = s3 ? tmp27988 : tmp27997;
  assign tmp27967 = s4 ? tmp27968 : tmp27987;
  assign tmp28008 = s0 ? tmp27975 : 1;
  assign tmp28009 = s0 ? 1 : tmp27979;
  assign tmp28007 = s1 ? tmp28008 : tmp28009;
  assign tmp28011 = s0 ? 1 : tmp27975;
  assign tmp28014 = l2 ? tmp27488 : 0;
  assign tmp28013 = l1 ? tmp28014 : tmp27509;
  assign tmp28012 = s0 ? tmp28013 : tmp27985;
  assign tmp28010 = s1 ? tmp28011 : tmp28012;
  assign tmp28006 = s2 ? tmp28007 : tmp28010;
  assign tmp28018 = l1 ? tmp28014 : tmp27490;
  assign tmp28017 = s0 ? tmp27985 : tmp28018;
  assign tmp28020 = ~(l1 ? 1 : tmp27887);
  assign tmp28019 = s0 ? tmp27985 : tmp28020;
  assign tmp28016 = s1 ? tmp28017 : tmp28019;
  assign tmp28021 = ~(s1 ? 1 : tmp28002);
  assign tmp28015 = s2 ? tmp28016 : tmp28021;
  assign tmp28005 = s3 ? tmp28006 : tmp28015;
  assign tmp28026 = ~(l1 ? tmp27971 : tmp27497);
  assign tmp28025 = s0 ? 1 : tmp28026;
  assign tmp28027 = ~(s0 ? tmp27991 : tmp27697);
  assign tmp28024 = s1 ? tmp28025 : tmp28027;
  assign tmp28029 = s0 ? tmp27991 : tmp27697;
  assign tmp28028 = ~(s1 ? tmp28029 : tmp27990);
  assign tmp28023 = s2 ? tmp28024 : tmp28028;
  assign tmp28033 = l1 ? 1 : tmp27506;
  assign tmp28034 = ~(l1 ? tmp28014 : 0);
  assign tmp28032 = s0 ? tmp28033 : tmp28034;
  assign tmp28035 = ~(s0 ? tmp27697 : 0);
  assign tmp28031 = s1 ? tmp28032 : tmp28035;
  assign tmp28030 = s2 ? tmp28031 : 1;
  assign tmp28022 = ~(s3 ? tmp28023 : tmp28030);
  assign tmp28004 = s4 ? tmp28005 : tmp28022;
  assign tmp28041 = l1 ? 1 : tmp27887;
  assign tmp28040 = s0 ? tmp28041 : 1;
  assign tmp28039 = s1 ? tmp28040 : 1;
  assign tmp28042 = s0 ? 1 : tmp28033;
  assign tmp28038 = s2 ? tmp28039 : tmp28042;
  assign tmp28037 = s3 ? tmp28038 : 1;
  assign tmp28046 = s0 ? tmp28033 : 1;
  assign tmp28045 = s1 ? tmp28042 : tmp28046;
  assign tmp28044 = s2 ? 1 : tmp28045;
  assign tmp28043 = s3 ? tmp28044 : 1;
  assign tmp28036 = ~(s4 ? tmp28037 : tmp28043);
  assign tmp28003 = s5 ? tmp28004 : tmp28036;
  assign tmp27966 = s6 ? tmp27967 : tmp28003;
  assign tmp27965 = ~(s7 ? tmp27966 : tmp27495);
  assign tmp27879 = s8 ? tmp27880 : tmp27965;
  assign tmp28048 = s7 ? tmp27966 : tmp27495;
  assign tmp28054 = l1 ? tmp27886 : tmp27684;
  assign tmp28056 = ~(l1 ? tmp27886 : tmp27553);
  assign tmp28055 = ~(s0 ? tmp27890 : tmp28056);
  assign tmp28053 = s1 ? tmp28054 : tmp28055;
  assign tmp28060 = l1 ? tmp27897 : tmp27695;
  assign tmp28061 = ~(l1 ? tmp27509 : tmp27508);
  assign tmp28059 = s0 ? tmp28060 : tmp28061;
  assign tmp28063 = l1 ? tmp27886 : tmp27695;
  assign tmp28062 = s0 ? tmp28063 : tmp28061;
  assign tmp28058 = s1 ? tmp28059 : tmp28062;
  assign tmp28065 = s0 ? tmp28063 : tmp27695;
  assign tmp28067 = l1 ? tmp27509 : tmp27508;
  assign tmp28068 = l1 ? tmp27509 : tmp27569;
  assign tmp28066 = ~(s0 ? tmp28067 : tmp28068);
  assign tmp28064 = s1 ? tmp28065 : tmp28066;
  assign tmp28057 = s2 ? tmp28058 : tmp28064;
  assign tmp28052 = s3 ? tmp28053 : tmp28057;
  assign tmp28073 = l1 ? tmp27897 : tmp27553;
  assign tmp28074 = ~(l1 ? tmp27490 : 1);
  assign tmp28072 = s0 ? tmp28073 : tmp28074;
  assign tmp28075 = ~(s0 ? tmp28068 : tmp28067);
  assign tmp28071 = s1 ? tmp28072 : tmp28075;
  assign tmp28077 = s0 ? tmp28054 : tmp27697;
  assign tmp28080 = l2 ? tmp27490 : tmp27554;
  assign tmp28079 = l1 ? tmp27490 : tmp28080;
  assign tmp28081 = ~(l1 ? tmp27504 : 0);
  assign tmp28078 = ~(s0 ? tmp28079 : tmp28081);
  assign tmp28076 = s1 ? tmp28077 : tmp28078;
  assign tmp28070 = s2 ? tmp28071 : tmp28076;
  assign tmp28084 = ~(s0 ? tmp27697 : tmp27750);
  assign tmp28083 = s1 ? tmp27890 : tmp28084;
  assign tmp28086 = ~(s0 ? tmp27750 : tmp28061);
  assign tmp28085 = s1 ? tmp28067 : tmp28086;
  assign tmp28082 = ~(s2 ? tmp28083 : tmp28085);
  assign tmp28069 = s3 ? tmp28070 : tmp28082;
  assign tmp28051 = s4 ? tmp28052 : tmp28069;
  assign tmp28093 = l1 ? tmp27886 : tmp27553;
  assign tmp28092 = s0 ? tmp28093 : 0;
  assign tmp28095 = ~(l1 ? tmp27897 : tmp27695);
  assign tmp28094 = ~(s0 ? 1 : tmp28095);
  assign tmp28091 = s1 ? tmp28092 : tmp28094;
  assign tmp28098 = ~(l1 ? tmp27886 : tmp27489);
  assign tmp28097 = s0 ? 1 : tmp28098;
  assign tmp28100 = l1 ? 1 : tmp27563;
  assign tmp28099 = ~(s0 ? tmp28100 : tmp27695);
  assign tmp28096 = ~(s1 ? tmp28097 : tmp28099);
  assign tmp28090 = s2 ? tmp28091 : tmp28096;
  assign tmp28104 = ~(l1 ? 1 : tmp27695);
  assign tmp28103 = s0 ? tmp27891 : tmp28104;
  assign tmp28106 = ~(l1 ? 1 : tmp27729);
  assign tmp28105 = s0 ? tmp27891 : tmp28106;
  assign tmp28102 = s1 ? tmp28103 : tmp28105;
  assign tmp28108 = ~(l1 ? tmp27509 : tmp27510);
  assign tmp28107 = ~(s1 ? tmp27750 : tmp28108);
  assign tmp28101 = ~(s2 ? tmp28102 : tmp28107);
  assign tmp28089 = s3 ? tmp28090 : tmp28101;
  assign tmp28113 = ~(l1 ? tmp27509 : tmp27521);
  assign tmp28112 = s0 ? tmp27750 : tmp28113;
  assign tmp28115 = l1 ? tmp27490 : 1;
  assign tmp28114 = ~(s0 ? tmp28115 : tmp27791);
  assign tmp28111 = s1 ? tmp28112 : tmp28114;
  assign tmp28117 = s0 ? tmp28115 : tmp27791;
  assign tmp28119 = l1 ? tmp27897 : tmp27489;
  assign tmp28118 = ~(s0 ? tmp28119 : tmp28074);
  assign tmp28116 = ~(s1 ? tmp28117 : tmp28118);
  assign tmp28110 = s2 ? tmp28111 : tmp28116;
  assign tmp28122 = s0 ? tmp27767 : tmp27750;
  assign tmp28121 = s1 ? tmp28122 : tmp27750;
  assign tmp28120 = s2 ? tmp28121 : tmp27750;
  assign tmp28109 = s3 ? tmp28110 : tmp28120;
  assign tmp28088 = s4 ? tmp28089 : tmp28109;
  assign tmp28128 = l1 ? 1 : tmp27729;
  assign tmp28127 = s0 ? tmp28128 : tmp27750;
  assign tmp28126 = s1 ? tmp28127 : tmp27750;
  assign tmp28130 = l1 ? 1 : tmp27553;
  assign tmp28129 = s0 ? tmp27750 : tmp28130;
  assign tmp28125 = s2 ? tmp28126 : tmp28129;
  assign tmp28124 = s3 ? tmp28125 : tmp27750;
  assign tmp28134 = s0 ? tmp27750 : tmp27767;
  assign tmp28135 = s0 ? tmp28130 : tmp27750;
  assign tmp28133 = s1 ? tmp28134 : tmp28135;
  assign tmp28132 = s2 ? tmp27750 : tmp28133;
  assign tmp28131 = s3 ? tmp28132 : tmp27750;
  assign tmp28123 = s4 ? tmp28124 : tmp28131;
  assign tmp28087 = s5 ? tmp28088 : tmp28123;
  assign tmp28050 = s6 ? tmp28051 : tmp28087;
  assign tmp28049 = ~(s7 ? tmp28050 : tmp27575);
  assign tmp28047 = ~(s8 ? tmp28048 : tmp28049);
  assign tmp27878 = s9 ? tmp27879 : tmp28047;
  assign tmp28144 = s0 ? tmp27909 : tmp27887;
  assign tmp28143 = s1 ? tmp28144 : tmp27899;
  assign tmp28146 = s0 ? tmp27900 : tmp27695;
  assign tmp28148 = l1 ? tmp27509 : tmp27972;
  assign tmp28147 = ~(s0 ? tmp27509 : tmp28148);
  assign tmp28145 = s1 ? tmp28146 : tmp28147;
  assign tmp28142 = s2 ? tmp28143 : tmp28145;
  assign tmp28141 = s3 ? tmp27884 : tmp28142;
  assign tmp28152 = s0 ? tmp27909 : tmp28074;
  assign tmp28153 = ~(s0 ? tmp28148 : tmp27509);
  assign tmp28151 = s1 ? tmp28152 : tmp28153;
  assign tmp28155 = s0 ? tmp27885 : tmp27697;
  assign tmp28156 = ~(s0 ? tmp27490 : tmp28081);
  assign tmp28154 = s1 ? tmp28155 : tmp28156;
  assign tmp28150 = s2 ? tmp28151 : tmp28154;
  assign tmp28159 = ~(s0 ? tmp27697 : 1);
  assign tmp28158 = s1 ? tmp27890 : tmp28159;
  assign tmp28157 = ~(s2 ? tmp28158 : tmp27918);
  assign tmp28149 = s3 ? tmp28150 : tmp28157;
  assign tmp28140 = s4 ? tmp28141 : tmp28149;
  assign tmp28165 = s0 ? tmp27900 : 0;
  assign tmp28167 = ~(l1 ? tmp27897 : tmp27506);
  assign tmp28166 = ~(s0 ? 1 : tmp28167);
  assign tmp28164 = s1 ? tmp28165 : tmp28166;
  assign tmp28169 = s0 ? 1 : tmp27892;
  assign tmp28170 = s0 ? tmp27509 : tmp27891;
  assign tmp28168 = ~(s1 ? tmp28169 : tmp28170);
  assign tmp28163 = s2 ? tmp28164 : tmp28168;
  assign tmp28173 = s0 ? tmp27891 : tmp27934;
  assign tmp28174 = s0 ? tmp27891 : tmp28020;
  assign tmp28172 = s1 ? tmp28173 : tmp28174;
  assign tmp28171 = ~(s2 ? tmp28172 : tmp27937);
  assign tmp28162 = s3 ? tmp28163 : tmp28171;
  assign tmp28179 = ~(l1 ? tmp27509 : tmp27497);
  assign tmp28178 = s0 ? 1 : tmp28179;
  assign tmp28180 = ~(s0 ? tmp28115 : 0);
  assign tmp28177 = s1 ? tmp28178 : tmp28180;
  assign tmp28182 = s0 ? tmp28115 : 0;
  assign tmp28183 = ~(s0 ? tmp27909 : tmp28074);
  assign tmp28181 = ~(s1 ? tmp28182 : tmp28183);
  assign tmp28176 = s2 ? tmp28177 : tmp28181;
  assign tmp28185 = s1 ? tmp28046 : 1;
  assign tmp28184 = s2 ? tmp28185 : 1;
  assign tmp28175 = s3 ? tmp28176 : tmp28184;
  assign tmp28161 = s4 ? tmp28162 : tmp28175;
  assign tmp28186 = s4 ? tmp28037 : tmp28043;
  assign tmp28160 = s5 ? tmp28161 : tmp28186;
  assign tmp28139 = s6 ? tmp28140 : tmp28160;
  assign tmp28138 = s7 ? tmp28139 : tmp27575;
  assign tmp28137 = s8 ? tmp28138 : tmp28139;
  assign tmp28136 = s9 ? tmp28137 : tmp27575;
  assign tmp27877 = s10 ? tmp27878 : tmp28136;
  assign tmp28196 = l1 ? tmp27490 : tmp27833;
  assign tmp28197 = ~(l1 ? tmp27886 : tmp27897);
  assign tmp28195 = ~(s0 ? tmp28196 : tmp28197);
  assign tmp28194 = s1 ? tmp27886 : tmp28195;
  assign tmp28200 = s0 ? tmp27897 : tmp27886;
  assign tmp28202 = l1 ? tmp27886 : tmp27897;
  assign tmp28201 = s0 ? tmp28202 : tmp27886;
  assign tmp28199 = s1 ? tmp28200 : tmp28201;
  assign tmp28205 = ~(l1 ? tmp27495 : tmp27833);
  assign tmp28204 = s0 ? tmp28202 : tmp28205;
  assign tmp28203 = s1 ? tmp28204 : tmp27886;
  assign tmp28198 = s2 ? tmp28199 : tmp28203;
  assign tmp28193 = s3 ? tmp28194 : tmp28198;
  assign tmp28210 = ~(l1 ? tmp27490 : tmp27833);
  assign tmp28209 = s0 ? tmp27897 : tmp28210;
  assign tmp28208 = s1 ? tmp28209 : tmp27886;
  assign tmp28212 = s0 ? tmp27886 : tmp27575;
  assign tmp28214 = l1 ? tmp27490 : 0;
  assign tmp28213 = ~(s0 ? tmp28214 : tmp27495);
  assign tmp28211 = s1 ? tmp28212 : tmp28213;
  assign tmp28207 = s2 ? tmp28208 : tmp28211;
  assign tmp28216 = s1 ? tmp28196 : tmp27917;
  assign tmp28218 = s0 ? 1 : tmp27886;
  assign tmp28217 = ~(s1 ? tmp27886 : tmp28218);
  assign tmp28215 = ~(s2 ? tmp28216 : tmp28217);
  assign tmp28206 = s3 ? tmp28207 : tmp28215;
  assign tmp28192 = s4 ? tmp28193 : tmp28206;
  assign tmp28225 = l1 ? tmp27495 : tmp27833;
  assign tmp28226 = ~(l2 ? 1 : tmp27506);
  assign tmp28224 = ~(s0 ? tmp28225 : tmp28226);
  assign tmp28223 = s1 ? tmp28204 : tmp28224;
  assign tmp28229 = ~(l1 ? tmp27886 : 1);
  assign tmp28228 = s0 ? tmp28225 : tmp28229;
  assign tmp28231 = l1 ? 1 : tmp27886;
  assign tmp28230 = ~(s0 ? tmp28231 : tmp27504);
  assign tmp28227 = ~(s1 ? tmp28228 : tmp28230);
  assign tmp28222 = s2 ? tmp28223 : tmp28227;
  assign tmp28235 = l1 ? 1 : tmp27897;
  assign tmp28234 = s0 ? tmp27504 : tmp28235;
  assign tmp28236 = s0 ? tmp27504 : 1;
  assign tmp28233 = s1 ? tmp28234 : tmp28236;
  assign tmp28239 = l1 ? tmp27886 : 1;
  assign tmp28238 = s0 ? tmp28239 : 1;
  assign tmp28237 = s1 ? 1 : tmp28238;
  assign tmp28232 = s2 ? tmp28233 : tmp28237;
  assign tmp28221 = s3 ? tmp28222 : tmp28232;
  assign tmp28243 = s0 ? 1 : tmp28239;
  assign tmp28244 = ~(s0 ? tmp28214 : 0);
  assign tmp28242 = s1 ? tmp28243 : tmp28244;
  assign tmp28246 = s0 ? tmp28214 : 0;
  assign tmp28248 = l1 ? tmp27897 : 1;
  assign tmp28249 = ~(l1 ? tmp27490 : 0);
  assign tmp28247 = ~(s0 ? tmp28248 : tmp28249);
  assign tmp28245 = ~(s1 ? tmp28246 : tmp28247);
  assign tmp28241 = s2 ? tmp28242 : tmp28245;
  assign tmp28240 = s3 ? tmp28241 : 1;
  assign tmp28220 = s4 ? tmp28221 : tmp28240;
  assign tmp28219 = s5 ? tmp28220 : 1;
  assign tmp28191 = s6 ? tmp28192 : tmp28219;
  assign tmp28190 = s7 ? tmp28191 : tmp27575;
  assign tmp28256 = ~(l2 ? 1 : tmp27887);
  assign tmp28255 = l1 ? tmp27971 : tmp28256;
  assign tmp28258 = l1 ? tmp27560 : tmp27833;
  assign tmp28259 = l1 ? tmp27971 : tmp28226;
  assign tmp28257 = s0 ? tmp28258 : tmp28259;
  assign tmp28254 = s1 ? tmp28255 : tmp28257;
  assign tmp28263 = l1 ? tmp27980 : tmp28226;
  assign tmp28262 = s0 ? tmp28263 : tmp28255;
  assign tmp28264 = s0 ? tmp28259 : tmp28255;
  assign tmp28261 = s1 ? tmp28262 : tmp28264;
  assign tmp28267 = l1 ? 1 : tmp27833;
  assign tmp28266 = s0 ? tmp28259 : tmp28267;
  assign tmp28265 = s1 ? tmp28266 : tmp28255;
  assign tmp28260 = s2 ? tmp28261 : tmp28265;
  assign tmp28253 = s3 ? tmp28254 : tmp28260;
  assign tmp28271 = s0 ? tmp28263 : tmp28258;
  assign tmp28270 = s1 ? tmp28271 : tmp28255;
  assign tmp28273 = s0 ? tmp28255 : 1;
  assign tmp28275 = l1 ? tmp27560 : 0;
  assign tmp28274 = s0 ? tmp28275 : 1;
  assign tmp28272 = s1 ? tmp28273 : tmp28274;
  assign tmp28269 = s2 ? tmp28270 : tmp28272;
  assign tmp28277 = s1 ? tmp28258 : tmp27999;
  assign tmp28280 = ~(l1 ? tmp27971 : tmp28256);
  assign tmp28279 = ~(s0 ? 1 : tmp28280);
  assign tmp28278 = s1 ? tmp28255 : tmp28279;
  assign tmp28276 = s2 ? tmp28277 : tmp28278;
  assign tmp28268 = s3 ? tmp28269 : tmp28276;
  assign tmp28252 = s4 ? tmp28253 : tmp28268;
  assign tmp28286 = s0 ? tmp28267 : tmp28263;
  assign tmp28285 = s1 ? tmp28266 : tmp28286;
  assign tmp28289 = l1 ? tmp27971 : 0;
  assign tmp28288 = s0 ? tmp28267 : tmp28289;
  assign tmp28291 = l1 ? tmp28014 : tmp28256;
  assign tmp28290 = s0 ? tmp28291 : tmp28267;
  assign tmp28287 = s1 ? tmp28288 : tmp28290;
  assign tmp28284 = s2 ? tmp28285 : tmp28287;
  assign tmp28295 = l1 ? tmp28014 : tmp28226;
  assign tmp28294 = s0 ? tmp28267 : tmp28295;
  assign tmp28296 = s0 ? tmp28267 : 0;
  assign tmp28293 = s1 ? tmp28294 : tmp28296;
  assign tmp28299 = l1 ? tmp28014 : 0;
  assign tmp28298 = ~(s0 ? tmp28289 : tmp28299);
  assign tmp28297 = ~(s1 ? 1 : tmp28298);
  assign tmp28292 = s2 ? tmp28293 : tmp28297;
  assign tmp28283 = s3 ? tmp28284 : tmp28292;
  assign tmp28304 = ~(l1 ? tmp27971 : 0);
  assign tmp28303 = s0 ? 1 : tmp28304;
  assign tmp28305 = ~(s0 ? tmp28275 : tmp27697);
  assign tmp28302 = s1 ? tmp28303 : tmp28305;
  assign tmp28307 = s0 ? tmp28275 : tmp27697;
  assign tmp28309 = l1 ? tmp27980 : 0;
  assign tmp28308 = s0 ? tmp28309 : tmp28275;
  assign tmp28306 = ~(s1 ? tmp28307 : tmp28308);
  assign tmp28301 = s2 ? tmp28302 : tmp28306;
  assign tmp28312 = s0 ? 1 : tmp28034;
  assign tmp28311 = s1 ? tmp28312 : tmp28035;
  assign tmp28310 = s2 ? tmp28311 : 1;
  assign tmp28300 = ~(s3 ? tmp28301 : tmp28310);
  assign tmp28282 = s4 ? tmp28283 : tmp28300;
  assign tmp28281 = s5 ? tmp28282 : 0;
  assign tmp28251 = s6 ? tmp28252 : tmp28281;
  assign tmp28250 = ~(s7 ? tmp28251 : tmp27495);
  assign tmp28189 = s8 ? tmp28190 : tmp28250;
  assign tmp28314 = s7 ? tmp28251 : tmp27495;
  assign tmp28320 = l1 ? tmp27886 : tmp27499;
  assign tmp28324 = ~(l3 ? 1 : tmp27488);
  assign tmp28323 = l2 ? 1 : tmp28324;
  assign tmp28322 = ~(l1 ? tmp27886 : tmp28323);
  assign tmp28321 = ~(s0 ? tmp28196 : tmp28322);
  assign tmp28319 = s1 ? tmp28320 : tmp28321;
  assign tmp28328 = l1 ? tmp27897 : tmp27504;
  assign tmp28329 = ~(l1 ? tmp27509 : tmp27606);
  assign tmp28327 = s0 ? tmp28328 : tmp28329;
  assign tmp28331 = l1 ? tmp27886 : tmp27504;
  assign tmp28330 = s0 ? tmp28331 : tmp28329;
  assign tmp28326 = s1 ? tmp28327 : tmp28330;
  assign tmp28333 = s0 ? tmp28331 : tmp27504;
  assign tmp28332 = s1 ? tmp28333 : tmp28329;
  assign tmp28325 = s2 ? tmp28326 : tmp28332;
  assign tmp28318 = s3 ? tmp28319 : tmp28325;
  assign tmp28338 = l1 ? tmp27897 : tmp28323;
  assign tmp28337 = s0 ? tmp28338 : tmp28210;
  assign tmp28336 = s1 ? tmp28337 : tmp28329;
  assign tmp28340 = s0 ? tmp28320 : tmp27697;
  assign tmp28342 = l1 ? tmp27490 : tmp27809;
  assign tmp28341 = ~(s0 ? tmp28342 : tmp28081);
  assign tmp28339 = s1 ? tmp28340 : tmp28341;
  assign tmp28335 = s2 ? tmp28336 : tmp28339;
  assign tmp28344 = s1 ? tmp28196 : tmp28084;
  assign tmp28346 = l1 ? tmp27509 : tmp27606;
  assign tmp28347 = ~(s0 ? tmp27750 : tmp28329);
  assign tmp28345 = s1 ? tmp28346 : tmp28347;
  assign tmp28343 = ~(s2 ? tmp28344 : tmp28345);
  assign tmp28334 = s3 ? tmp28335 : tmp28343;
  assign tmp28317 = s4 ? tmp28318 : tmp28334;
  assign tmp28354 = l1 ? tmp27886 : tmp28323;
  assign tmp28355 = ~(l1 ? 1 : tmp27833);
  assign tmp28353 = s0 ? tmp28354 : tmp28355;
  assign tmp28357 = ~(l1 ? tmp27897 : tmp27504);
  assign tmp28356 = ~(s0 ? tmp28267 : tmp28357);
  assign tmp28352 = s1 ? tmp28353 : tmp28356;
  assign tmp28360 = ~(l1 ? tmp27886 : tmp27744);
  assign tmp28359 = s0 ? tmp28267 : tmp28360;
  assign tmp28362 = l1 ? 1 : tmp27499;
  assign tmp28361 = ~(s0 ? tmp28362 : tmp27636);
  assign tmp28358 = ~(s1 ? tmp28359 : tmp28361);
  assign tmp28351 = s2 ? tmp28352 : tmp28358;
  assign tmp28365 = s0 ? tmp27636 : tmp27750;
  assign tmp28364 = s1 ? tmp27636 : tmp28365;
  assign tmp28368 = l1 ? tmp27509 : tmp27809;
  assign tmp28367 = ~(s0 ? tmp28368 : tmp27791);
  assign tmp28366 = s1 ? tmp27750 : tmp28367;
  assign tmp28363 = s2 ? tmp28364 : tmp28366;
  assign tmp28350 = s3 ? tmp28351 : tmp28363;
  assign tmp28373 = ~(l1 ? tmp27509 : tmp27809);
  assign tmp28372 = s0 ? tmp27750 : tmp28373;
  assign tmp28374 = ~(s0 ? tmp28342 : tmp27791);
  assign tmp28371 = s1 ? tmp28372 : tmp28374;
  assign tmp28376 = s0 ? tmp28342 : tmp27791;
  assign tmp28378 = l1 ? tmp27897 : tmp27744;
  assign tmp28379 = ~(l1 ? tmp27490 : tmp27809);
  assign tmp28377 = ~(s0 ? tmp28378 : tmp28379);
  assign tmp28375 = ~(s1 ? tmp28376 : tmp28377);
  assign tmp28370 = s2 ? tmp28371 : tmp28375;
  assign tmp28369 = s3 ? tmp28370 : tmp27750;
  assign tmp28349 = s4 ? tmp28350 : tmp28369;
  assign tmp28348 = s5 ? tmp28349 : tmp27750;
  assign tmp28316 = s6 ? tmp28317 : tmp28348;
  assign tmp28315 = ~(s7 ? tmp28316 : tmp27575);
  assign tmp28313 = ~(s8 ? tmp28314 : tmp28315);
  assign tmp28188 = s9 ? tmp28189 : tmp28313;
  assign tmp28389 = ~(l1 ? tmp27509 : tmp28256);
  assign tmp28388 = s0 ? tmp27897 : tmp28389;
  assign tmp28390 = s0 ? tmp28202 : tmp28389;
  assign tmp28387 = s1 ? tmp28388 : tmp28390;
  assign tmp28392 = s0 ? tmp28202 : tmp27504;
  assign tmp28391 = s1 ? tmp28392 : tmp28389;
  assign tmp28386 = s2 ? tmp28387 : tmp28391;
  assign tmp28385 = s3 ? tmp28194 : tmp28386;
  assign tmp28395 = s1 ? tmp28209 : tmp28389;
  assign tmp28397 = s0 ? tmp27886 : tmp27697;
  assign tmp28398 = ~(s0 ? tmp28214 : tmp28081);
  assign tmp28396 = s1 ? tmp28397 : tmp28398;
  assign tmp28394 = s2 ? tmp28395 : tmp28396;
  assign tmp28400 = s1 ? tmp28196 : tmp28159;
  assign tmp28402 = l1 ? tmp27509 : tmp28256;
  assign tmp28403 = ~(s0 ? 1 : tmp28389);
  assign tmp28401 = s1 ? tmp28402 : tmp28403;
  assign tmp28399 = ~(s2 ? tmp28400 : tmp28401);
  assign tmp28393 = s3 ? tmp28394 : tmp28399;
  assign tmp28384 = s4 ? tmp28385 : tmp28393;
  assign tmp28409 = s0 ? tmp28202 : tmp28355;
  assign tmp28410 = ~(s0 ? tmp28267 : tmp28226);
  assign tmp28408 = s1 ? tmp28409 : tmp28410;
  assign tmp28412 = s0 ? tmp28267 : tmp28229;
  assign tmp28413 = ~(s0 ? tmp28231 : tmp27636);
  assign tmp28411 = ~(s1 ? tmp28412 : tmp28413);
  assign tmp28407 = s2 ? tmp28408 : tmp28411;
  assign tmp28416 = s0 ? tmp27636 : tmp28235;
  assign tmp28417 = s0 ? tmp27636 : 1;
  assign tmp28415 = s1 ? tmp28416 : tmp28417;
  assign tmp28420 = l1 ? tmp27509 : 0;
  assign tmp28419 = ~(s0 ? tmp28420 : 0);
  assign tmp28418 = s1 ? 1 : tmp28419;
  assign tmp28414 = s2 ? tmp28415 : tmp28418;
  assign tmp28406 = s3 ? tmp28407 : tmp28414;
  assign tmp28425 = ~(l1 ? tmp27509 : 0);
  assign tmp28424 = s0 ? 1 : tmp28425;
  assign tmp28423 = s1 ? tmp28424 : tmp28244;
  assign tmp28422 = s2 ? tmp28423 : tmp28245;
  assign tmp28421 = s3 ? tmp28422 : 1;
  assign tmp28405 = s4 ? tmp28406 : tmp28421;
  assign tmp28404 = s5 ? tmp28405 : 1;
  assign tmp28383 = s6 ? tmp28384 : tmp28404;
  assign tmp28382 = s7 ? tmp28383 : tmp27575;
  assign tmp28381 = s8 ? tmp28382 : tmp28383;
  assign tmp28380 = s9 ? tmp28381 : tmp27575;
  assign tmp28187 = s10 ? tmp28188 : tmp28380;
  assign tmp27876 = s12 ? tmp27877 : tmp28187;
  assign tmp27476 = s13 ? tmp27477 : tmp27876;
  assign tmp28436 = l1 ? 1 : tmp27888;
  assign tmp28438 = l1 ? 1 : tmp27695;
  assign tmp28437 = s0 ? tmp28438 : tmp28033;
  assign tmp28435 = s1 ? tmp28436 : tmp28437;
  assign tmp28442 = l1 ? 1 : tmp27898;
  assign tmp28441 = s0 ? tmp28442 : tmp28041;
  assign tmp28443 = s0 ? tmp28033 : tmp28041;
  assign tmp28440 = s1 ? tmp28441 : tmp28443;
  assign tmp28446 = l1 ? 1 : tmp27575;
  assign tmp28445 = s0 ? tmp28033 : tmp28446;
  assign tmp28447 = s0 ? tmp28041 : tmp28436;
  assign tmp28444 = s1 ? tmp28445 : tmp28447;
  assign tmp28439 = s2 ? tmp28440 : tmp28444;
  assign tmp28434 = s3 ? tmp28435 : tmp28439;
  assign tmp28451 = s0 ? tmp28436 : tmp28041;
  assign tmp28450 = s1 ? tmp28445 : tmp28451;
  assign tmp28453 = s0 ? tmp28436 : tmp28446;
  assign tmp28452 = s1 ? tmp28453 : tmp28445;
  assign tmp28449 = s2 ? tmp28450 : tmp28452;
  assign tmp28456 = s0 ? tmp28446 : 1;
  assign tmp28455 = s1 ? tmp28438 : tmp28456;
  assign tmp28458 = s0 ? tmp28041 : tmp27887;
  assign tmp28459 = s0 ? 1 : tmp28041;
  assign tmp28457 = s1 ? tmp28458 : tmp28459;
  assign tmp28454 = s2 ? tmp28455 : tmp28457;
  assign tmp28448 = s3 ? tmp28449 : tmp28454;
  assign tmp28433 = s4 ? tmp28434 : tmp28448;
  assign tmp28465 = s0 ? tmp28446 : tmp28442;
  assign tmp28464 = s1 ? tmp28445 : tmp28465;
  assign tmp28467 = s0 ? tmp28446 : tmp27858;
  assign tmp28468 = ~(s0 ? tmp27509 : tmp27495);
  assign tmp28466 = s1 ? tmp28467 : tmp28468;
  assign tmp28463 = s2 ? tmp28464 : tmp28466;
  assign tmp28473 = ~(l2 ? tmp27509 : 0);
  assign tmp28472 = l1 ? 1 : tmp28473;
  assign tmp28471 = s0 ? tmp28472 : 1;
  assign tmp28470 = ~(s1 ? 1 : tmp28471);
  assign tmp28469 = ~(s2 ? tmp27932 : tmp28470);
  assign tmp28462 = s3 ? tmp28463 : tmp28469;
  assign tmp28476 = s1 ? tmp27964 : tmp28456;
  assign tmp28478 = s0 ? tmp27858 : tmp28446;
  assign tmp28477 = s1 ? tmp28456 : tmp28478;
  assign tmp28475 = s2 ? tmp28476 : tmp28477;
  assign tmp28474 = s3 ? tmp28475 : tmp27949;
  assign tmp28461 = s4 ? tmp28462 : tmp28474;
  assign tmp28460 = s5 ? tmp28461 : tmp27952;
  assign tmp28432 = s6 ? tmp28433 : tmp28460;
  assign tmp28431 = s7 ? tmp28432 : tmp27575;
  assign tmp28485 = ~(l2 ? tmp27554 : tmp27509);
  assign tmp28484 = l1 ? 1 : tmp28485;
  assign tmp28488 = ~(l2 ? tmp27554 : 1);
  assign tmp28487 = l1 ? 1 : tmp28488;
  assign tmp28490 = ~(l2 ? tmp27554 : tmp27490);
  assign tmp28489 = l1 ? 1 : tmp28490;
  assign tmp28486 = s0 ? tmp28487 : tmp28489;
  assign tmp28483 = s1 ? tmp28484 : tmp28486;
  assign tmp28495 = ~(l2 ? 1 : tmp27490);
  assign tmp28494 = l1 ? 1 : tmp28495;
  assign tmp28497 = ~(l2 ? tmp27488 : tmp27509);
  assign tmp28496 = l1 ? 1 : tmp28497;
  assign tmp28493 = s0 ? tmp28494 : tmp28496;
  assign tmp28498 = s0 ? tmp28489 : tmp28496;
  assign tmp28492 = s1 ? tmp28493 : tmp28498;
  assign tmp28500 = s0 ? tmp28489 : tmp27640;
  assign tmp28501 = s0 ? tmp28496 : tmp28484;
  assign tmp28499 = s1 ? tmp28500 : tmp28501;
  assign tmp28491 = s2 ? tmp28492 : tmp28499;
  assign tmp28482 = s3 ? tmp28483 : tmp28491;
  assign tmp28505 = s0 ? tmp28484 : tmp28496;
  assign tmp28504 = s1 ? tmp28500 : tmp28505;
  assign tmp28507 = s0 ? tmp28484 : tmp27640;
  assign tmp28509 = l1 ? 1 : tmp28324;
  assign tmp28508 = s0 ? tmp28509 : tmp27640;
  assign tmp28506 = s1 ? tmp28507 : tmp28508;
  assign tmp28503 = s2 ? tmp28504 : tmp28506;
  assign tmp28512 = s0 ? tmp27640 : 1;
  assign tmp28511 = s1 ? tmp28487 : tmp28512;
  assign tmp28515 = ~(l1 ? 1 : tmp28497);
  assign tmp28514 = ~(s0 ? tmp27488 : tmp28515);
  assign tmp28513 = s1 ? tmp28496 : tmp28514;
  assign tmp28510 = s2 ? tmp28511 : tmp28513;
  assign tmp28502 = s3 ? tmp28503 : tmp28510;
  assign tmp28481 = s4 ? tmp28482 : tmp28502;
  assign tmp28521 = s0 ? tmp27640 : tmp28494;
  assign tmp28520 = s1 ? tmp28500 : tmp28521;
  assign tmp28525 = ~(l2 ? tmp27554 : 0);
  assign tmp28524 = l1 ? 1 : tmp28525;
  assign tmp28523 = s0 ? tmp27640 : tmp28524;
  assign tmp28526 = s0 ? tmp28496 : tmp27640;
  assign tmp28522 = s1 ? tmp28523 : tmp28526;
  assign tmp28519 = s2 ? tmp28520 : tmp28522;
  assign tmp28529 = s0 ? tmp27640 : tmp28489;
  assign tmp28531 = ~(l2 ? tmp27488 : 0);
  assign tmp28530 = s0 ? tmp27640 : tmp28531;
  assign tmp28528 = s1 ? tmp28529 : tmp28530;
  assign tmp28533 = s0 ? tmp27488 : 0;
  assign tmp28534 = ~(l1 ? 1 : tmp28531);
  assign tmp28532 = ~(s1 ? tmp28533 : tmp28534);
  assign tmp28527 = s2 ? tmp28528 : tmp28532;
  assign tmp28518 = s3 ? tmp28519 : tmp28527;
  assign tmp28538 = s0 ? 1 : tmp28524;
  assign tmp28540 = l1 ? 1 : tmp27492;
  assign tmp28539 = s0 ? tmp27640 : tmp28540;
  assign tmp28537 = s1 ? tmp28538 : tmp28539;
  assign tmp28542 = s0 ? tmp28524 : tmp27640;
  assign tmp28541 = s1 ? tmp28539 : tmp28542;
  assign tmp28536 = s2 ? tmp28537 : tmp28541;
  assign tmp28546 = l1 ? 1 : tmp28531;
  assign tmp28545 = s0 ? tmp28524 : tmp28546;
  assign tmp28547 = s0 ? tmp28540 : 1;
  assign tmp28544 = s1 ? tmp28545 : tmp28547;
  assign tmp28543 = s2 ? tmp28544 : 1;
  assign tmp28535 = s3 ? tmp28536 : tmp28543;
  assign tmp28517 = s4 ? tmp28518 : tmp28535;
  assign tmp28552 = s0 ? tmp28014 : 0;
  assign tmp28553 = ~(s0 ? 1 : tmp28540);
  assign tmp28551 = s1 ? tmp28552 : tmp28553;
  assign tmp28555 = s0 ? tmp28540 : tmp28267;
  assign tmp28554 = ~(s1 ? tmp28555 : tmp28267);
  assign tmp28550 = s2 ? tmp28551 : tmp28554;
  assign tmp28549 = s3 ? tmp28550 : 0;
  assign tmp28559 = s0 ? 1 : tmp27492;
  assign tmp28558 = s1 ? 1 : tmp28559;
  assign tmp28560 = s1 ? tmp28538 : tmp28267;
  assign tmp28557 = s2 ? tmp28558 : tmp28560;
  assign tmp28562 = s1 ? tmp28547 : 1;
  assign tmp28561 = s2 ? tmp28562 : 1;
  assign tmp28556 = ~(s3 ? tmp28557 : tmp28561);
  assign tmp28548 = ~(s4 ? tmp28549 : tmp28556);
  assign tmp28516 = s5 ? tmp28517 : tmp28548;
  assign tmp28480 = s6 ? tmp28481 : tmp28516;
  assign tmp28479 = s7 ? tmp28480 : tmp27575;
  assign tmp28430 = s8 ? tmp28431 : tmp28479;
  assign tmp28570 = ~(l2 ? tmp27554 : tmp27488);
  assign tmp28569 = l1 ? 1 : tmp28570;
  assign tmp28571 = s0 ? tmp28487 : tmp28509;
  assign tmp28568 = s1 ? tmp28569 : tmp28571;
  assign tmp28574 = s0 ? tmp28487 : tmp28540;
  assign tmp28573 = s1 ? tmp28539 : tmp28574;
  assign tmp28576 = s0 ? tmp28487 : tmp27640;
  assign tmp28577 = s0 ? tmp28540 : tmp28569;
  assign tmp28575 = s1 ? tmp28576 : tmp28577;
  assign tmp28572 = s2 ? tmp28573 : tmp28575;
  assign tmp28567 = s3 ? tmp28568 : tmp28572;
  assign tmp28581 = s0 ? tmp28569 : tmp28540;
  assign tmp28580 = s1 ? tmp28508 : tmp28581;
  assign tmp28583 = s0 ? tmp28569 : tmp27640;
  assign tmp28582 = s1 ? tmp28583 : tmp28508;
  assign tmp28579 = s2 ? tmp28580 : tmp28582;
  assign tmp28586 = s0 ? tmp27640 : tmp27750;
  assign tmp28585 = s1 ? tmp28487 : tmp28586;
  assign tmp28589 = ~(l1 ? 1 : tmp27492);
  assign tmp28588 = ~(s0 ? tmp27488 : tmp28589);
  assign tmp28587 = s1 ? tmp28540 : tmp28588;
  assign tmp28584 = s2 ? tmp28585 : tmp28587;
  assign tmp28578 = s3 ? tmp28579 : tmp28584;
  assign tmp28566 = s4 ? tmp28567 : tmp28578;
  assign tmp28594 = s1 ? tmp28508 : tmp27640;
  assign tmp28596 = s0 ? tmp27640 : tmp28509;
  assign tmp28597 = s0 ? tmp28540 : tmp27640;
  assign tmp28595 = s1 ? tmp28596 : tmp28597;
  assign tmp28593 = s2 ? tmp28594 : tmp28595;
  assign tmp28600 = s0 ? tmp27640 : tmp28487;
  assign tmp28599 = s1 ? tmp28600 : tmp28539;
  assign tmp28602 = s0 ? tmp27488 : tmp27791;
  assign tmp28601 = ~(s1 ? tmp28602 : tmp28589);
  assign tmp28598 = s2 ? tmp28599 : tmp28601;
  assign tmp28592 = s3 ? tmp28593 : tmp28598;
  assign tmp28608 = ~(l2 ? tmp27554 : tmp27491);
  assign tmp28607 = l1 ? 1 : tmp28608;
  assign tmp28606 = s0 ? tmp27750 : tmp28607;
  assign tmp28605 = s1 ? tmp28606 : tmp28539;
  assign tmp28609 = s1 ? tmp28539 : tmp28508;
  assign tmp28604 = s2 ? tmp28605 : tmp28609;
  assign tmp28614 = ~(l2 ? tmp27488 : tmp27491);
  assign tmp28613 = l1 ? 1 : tmp28614;
  assign tmp28612 = s0 ? tmp28509 : tmp28613;
  assign tmp28615 = s0 ? tmp28540 : tmp27750;
  assign tmp28611 = s1 ? tmp28612 : tmp28615;
  assign tmp28610 = s2 ? tmp28611 : tmp27750;
  assign tmp28603 = s3 ? tmp28604 : tmp28610;
  assign tmp28591 = s4 ? tmp28592 : tmp28603;
  assign tmp28620 = s0 ? tmp27750 : tmp28540;
  assign tmp28619 = s1 ? tmp28615 : tmp28620;
  assign tmp28621 = s1 ? tmp28597 : tmp27640;
  assign tmp28618 = s2 ? tmp28619 : tmp28621;
  assign tmp28617 = s3 ? tmp28618 : tmp27750;
  assign tmp28625 = s0 ? tmp27750 : tmp27492;
  assign tmp28624 = s1 ? tmp27750 : tmp28625;
  assign tmp28627 = s0 ? tmp27750 : tmp28509;
  assign tmp28626 = s1 ? tmp28627 : tmp27640;
  assign tmp28623 = s2 ? tmp28624 : tmp28626;
  assign tmp28629 = s1 ? tmp28615 : tmp27750;
  assign tmp28628 = s2 ? tmp28629 : tmp27750;
  assign tmp28622 = s3 ? tmp28623 : tmp28628;
  assign tmp28616 = s4 ? tmp28617 : tmp28622;
  assign tmp28590 = s5 ? tmp28591 : tmp28616;
  assign tmp28565 = s6 ? tmp28566 : tmp28590;
  assign tmp28564 = s7 ? tmp28565 : tmp27575;
  assign tmp28563 = s8 ? tmp28479 : tmp28564;
  assign tmp28429 = s9 ? tmp28430 : tmp28563;
  assign tmp28631 = s8 ? tmp28479 : tmp28480;
  assign tmp28630 = s9 ? tmp28631 : tmp27575;
  assign tmp28428 = s10 ? tmp28429 : tmp28630;
  assign tmp28641 = l2 ? tmp27554 : tmp27496;
  assign tmp28640 = l1 ? tmp27560 : tmp28641;
  assign tmp28643 = l2 ? tmp27554 : tmp27490;
  assign tmp28644 = l1 ? tmp27744 : tmp28641;
  assign tmp28642 = s0 ? tmp28643 : tmp28644;
  assign tmp28639 = s1 ? tmp28640 : tmp28642;
  assign tmp28647 = l1 ? tmp27560 : tmp28643;
  assign tmp28646 = s0 ? tmp28647 : tmp28644;
  assign tmp28649 = s0 ? tmp28647 : 1;
  assign tmp28648 = s1 ? tmp28649 : tmp28644;
  assign tmp28645 = s2 ? tmp28646 : tmp28648;
  assign tmp28638 = s3 ? tmp28639 : tmp28645;
  assign tmp28654 = l1 ? tmp28643 : 1;
  assign tmp28653 = s0 ? tmp28640 : tmp28654;
  assign tmp28652 = s1 ? tmp28653 : tmp28644;
  assign tmp28656 = s0 ? tmp28640 : 1;
  assign tmp28657 = s0 ? tmp28643 : 1;
  assign tmp28655 = s1 ? tmp28656 : tmp28657;
  assign tmp28651 = s2 ? tmp28652 : tmp28655;
  assign tmp28661 = l2 ? tmp27554 : 1;
  assign tmp28660 = s0 ? 1 : tmp28661;
  assign tmp28659 = s1 ? tmp28643 : tmp28660;
  assign tmp28665 = ~(l2 ? tmp27554 : tmp27496);
  assign tmp28664 = ~(l1 ? tmp27508 : tmp28665);
  assign tmp28663 = s0 ? tmp28644 : tmp28664;
  assign tmp28667 = l1 ? 1 : tmp28661;
  assign tmp28666 = s0 ? tmp28667 : tmp28644;
  assign tmp28662 = s1 ? tmp28663 : tmp28666;
  assign tmp28658 = s2 ? tmp28659 : tmp28662;
  assign tmp28650 = s3 ? tmp28651 : tmp28658;
  assign tmp28637 = s4 ? tmp28638 : tmp28650;
  assign tmp28673 = s0 ? tmp28644 : 1;
  assign tmp28674 = s0 ? 1 : tmp28647;
  assign tmp28672 = s1 ? tmp28673 : tmp28674;
  assign tmp28678 = l2 ? tmp27554 : tmp27492;
  assign tmp28677 = l1 ? tmp27744 : tmp28678;
  assign tmp28676 = s0 ? 1 : tmp28677;
  assign tmp28680 = l1 ? tmp27508 : tmp28665;
  assign tmp28679 = ~(s0 ? tmp28680 : 0);
  assign tmp28675 = s1 ? tmp28676 : tmp28679;
  assign tmp28671 = s2 ? tmp28672 : tmp28675;
  assign tmp28685 = ~(l2 ? tmp27554 : tmp27492);
  assign tmp28684 = ~(l1 ? tmp27508 : tmp28685);
  assign tmp28683 = s0 ? 1 : tmp28684;
  assign tmp28682 = s1 ? tmp28674 : tmp28683;
  assign tmp28687 = s0 ? tmp28667 : 1;
  assign tmp28688 = s0 ? tmp28677 : tmp28684;
  assign tmp28686 = s1 ? tmp28687 : tmp28688;
  assign tmp28681 = s2 ? tmp28682 : tmp28686;
  assign tmp28670 = s3 ? tmp28671 : tmp28681;
  assign tmp28692 = s0 ? tmp28667 : tmp28677;
  assign tmp28693 = s0 ? tmp28654 : tmp27575;
  assign tmp28691 = s1 ? tmp28692 : tmp28693;
  assign tmp28696 = l1 ? tmp27560 : tmp28678;
  assign tmp28695 = s0 ? tmp28696 : tmp28654;
  assign tmp28694 = s1 ? tmp28693 : tmp28695;
  assign tmp28690 = s2 ? tmp28691 : tmp28694;
  assign tmp28700 = l1 ? tmp27504 : tmp28678;
  assign tmp28702 = ~(l2 ? tmp27496 : tmp27488);
  assign tmp28701 = l1 ? tmp27560 : tmp28702;
  assign tmp28699 = s0 ? tmp28700 : tmp28701;
  assign tmp28704 = l1 ? tmp27508 : tmp28685;
  assign tmp28703 = ~(s0 ? tmp27495 : tmp28704);
  assign tmp28698 = s1 ? tmp28699 : tmp28703;
  assign tmp28706 = s0 ? tmp28661 : 1;
  assign tmp28705 = s1 ? 1 : tmp28706;
  assign tmp28697 = s2 ? tmp28698 : tmp28705;
  assign tmp28689 = s3 ? tmp28690 : tmp28697;
  assign tmp28669 = s4 ? tmp28670 : tmp28689;
  assign tmp28711 = s0 ? tmp28704 : 0;
  assign tmp28712 = ~(s0 ? 1 : tmp28446);
  assign tmp28710 = s1 ? tmp28711 : tmp28712;
  assign tmp28714 = s0 ? tmp28446 : tmp27504;
  assign tmp28715 = s0 ? tmp27588 : tmp27504;
  assign tmp28713 = ~(s1 ? tmp28714 : tmp28715);
  assign tmp28709 = s2 ? tmp28710 : tmp28713;
  assign tmp28719 = l1 ? tmp27504 : tmp28702;
  assign tmp28718 = s0 ? tmp27959 : tmp28719;
  assign tmp28717 = s1 ? tmp27958 : tmp28718;
  assign tmp28716 = ~(s2 ? tmp27590 : tmp28717);
  assign tmp28708 = s3 ? tmp28709 : tmp28716;
  assign tmp28723 = s0 ? tmp28719 : 1;
  assign tmp28724 = s0 ? 1 : tmp28667;
  assign tmp28722 = s1 ? tmp28723 : tmp28724;
  assign tmp28727 = l1 ? tmp27499 : tmp28678;
  assign tmp28726 = s0 ? 1 : tmp28727;
  assign tmp28728 = s0 ? tmp27504 : tmp27588;
  assign tmp28725 = s1 ? tmp28726 : tmp28728;
  assign tmp28721 = s2 ? tmp28722 : tmp28725;
  assign tmp28733 = l2 ? tmp27496 : tmp27488;
  assign tmp28732 = ~(l1 ? tmp27508 : tmp28733);
  assign tmp28731 = s0 ? 1 : tmp28732;
  assign tmp28730 = s1 ? tmp28456 : tmp28731;
  assign tmp28734 = s1 ? tmp28718 : 1;
  assign tmp28729 = s2 ? tmp28730 : tmp28734;
  assign tmp28720 = ~(s3 ? tmp28721 : tmp28729);
  assign tmp28707 = ~(s4 ? tmp28708 : tmp28720);
  assign tmp28668 = s5 ? tmp28669 : tmp28707;
  assign tmp28636 = s6 ? tmp28637 : tmp28668;
  assign tmp28635 = s7 ? tmp28636 : tmp27575;
  assign tmp28741 = l2 ? tmp27488 : tmp27496;
  assign tmp28740 = l1 ? tmp27560 : tmp28741;
  assign tmp28743 = l1 ? tmp27560 : tmp27623;
  assign tmp28744 = l1 ? tmp27744 : tmp28741;
  assign tmp28742 = s0 ? tmp28743 : tmp28744;
  assign tmp28739 = s1 ? tmp28740 : tmp28742;
  assign tmp28747 = s0 ? tmp27560 : tmp28644;
  assign tmp28749 = l1 ? tmp27560 : tmp27980;
  assign tmp28748 = s0 ? tmp28749 : tmp28644;
  assign tmp28746 = s1 ? tmp28747 : tmp28748;
  assign tmp28751 = s0 ? tmp28749 : 1;
  assign tmp28752 = s0 ? tmp28644 : tmp28744;
  assign tmp28750 = s1 ? tmp28751 : tmp28752;
  assign tmp28745 = s2 ? tmp28746 : tmp28750;
  assign tmp28738 = s3 ? tmp28739 : tmp28745;
  assign tmp28756 = s0 ? tmp28740 : tmp27991;
  assign tmp28757 = s0 ? tmp28744 : tmp28644;
  assign tmp28755 = s1 ? tmp28756 : tmp28757;
  assign tmp28759 = s0 ? tmp28740 : 1;
  assign tmp28761 = l1 ? tmp27560 : tmp27488;
  assign tmp28760 = s0 ? tmp28761 : 1;
  assign tmp28758 = s1 ? tmp28759 : tmp28760;
  assign tmp28754 = s2 ? tmp28755 : tmp28758;
  assign tmp28764 = s0 ? tmp28761 : tmp28743;
  assign tmp28765 = s0 ? 1 : tmp27891;
  assign tmp28763 = s1 ? tmp28764 : tmp28765;
  assign tmp28768 = l1 ? tmp27499 : tmp28641;
  assign tmp28767 = s0 ? tmp28644 : tmp28768;
  assign tmp28766 = s1 ? tmp28767 : tmp28666;
  assign tmp28762 = s2 ? tmp28763 : tmp28766;
  assign tmp28753 = s3 ? tmp28754 : tmp28762;
  assign tmp28737 = s4 ? tmp28738 : tmp28753;
  assign tmp28774 = s0 ? tmp28744 : 1;
  assign tmp28775 = s0 ? 1 : tmp27560;
  assign tmp28773 = s1 ? tmp28774 : tmp28775;
  assign tmp28779 = l2 ? tmp27488 : tmp27492;
  assign tmp28778 = l1 ? tmp27744 : tmp28779;
  assign tmp28777 = s0 ? 1 : tmp28778;
  assign tmp28780 = s0 ? tmp28768 : 1;
  assign tmp28776 = s1 ? tmp28777 : tmp28780;
  assign tmp28772 = s2 ? tmp28773 : tmp28776;
  assign tmp28783 = s0 ? 1 : tmp28749;
  assign tmp28785 = ~(l1 ? tmp27488 : tmp28685);
  assign tmp28784 = s0 ? 1 : tmp28785;
  assign tmp28782 = s1 ? tmp28783 : tmp28784;
  assign tmp28787 = s0 ? tmp28677 : tmp28727;
  assign tmp28786 = s1 ? tmp28687 : tmp28787;
  assign tmp28781 = s2 ? tmp28782 : tmp28786;
  assign tmp28771 = s3 ? tmp28772 : tmp28781;
  assign tmp28791 = s0 ? tmp27985 : tmp28778;
  assign tmp28792 = s0 ? tmp27991 : tmp28014;
  assign tmp28790 = s1 ? tmp28791 : tmp28792;
  assign tmp28795 = l1 ? tmp27560 : tmp28779;
  assign tmp28794 = s0 ? tmp28795 : tmp27991;
  assign tmp28793 = s1 ? tmp28792 : tmp28794;
  assign tmp28789 = s2 ? tmp28790 : tmp28793;
  assign tmp28799 = l1 ? tmp27504 : tmp28779;
  assign tmp28798 = s0 ? tmp28799 : tmp28795;
  assign tmp28802 = ~(l2 ? tmp27490 : tmp27492);
  assign tmp28801 = ~(l1 ? tmp27488 : tmp28802);
  assign tmp28800 = s0 ? tmp28014 : tmp28801;
  assign tmp28797 = s1 ? tmp28798 : tmp28800;
  assign tmp28804 = s0 ? tmp27891 : 1;
  assign tmp28803 = s1 ? 1 : tmp28804;
  assign tmp28796 = s2 ? tmp28797 : tmp28803;
  assign tmp28788 = s3 ? tmp28789 : tmp28796;
  assign tmp28770 = s4 ? tmp28771 : tmp28788;
  assign tmp28810 = l1 ? tmp27488 : tmp28685;
  assign tmp28809 = s0 ? tmp28810 : 0;
  assign tmp28812 = l1 ? 1 : tmp27488;
  assign tmp28811 = ~(s0 ? 1 : tmp28812);
  assign tmp28808 = s1 ? tmp28809 : tmp28811;
  assign tmp28814 = s0 ? tmp28812 : tmp27504;
  assign tmp28815 = s0 ? tmp27697 : tmp27504;
  assign tmp28813 = ~(s1 ? tmp28814 : tmp28815);
  assign tmp28807 = s2 ? tmp28808 : tmp28813;
  assign tmp28818 = s0 ? 1 : tmp28267;
  assign tmp28821 = ~(l2 ? 1 : tmp27488);
  assign tmp28820 = l1 ? tmp27504 : tmp28821;
  assign tmp28819 = s0 ? tmp28267 : tmp28820;
  assign tmp28817 = s1 ? tmp28818 : tmp28819;
  assign tmp28816 = ~(s2 ? tmp27699 : tmp28817);
  assign tmp28806 = s3 ? tmp28807 : tmp28816;
  assign tmp28825 = s0 ? tmp28820 : 1;
  assign tmp28824 = s1 ? tmp28825 : tmp28724;
  assign tmp28828 = l1 ? tmp27499 : tmp28779;
  assign tmp28827 = s0 ? 1 : tmp28828;
  assign tmp28829 = s0 ? tmp27504 : tmp27697;
  assign tmp28826 = s1 ? tmp28827 : tmp28829;
  assign tmp28823 = s2 ? tmp28824 : tmp28826;
  assign tmp28832 = s0 ? tmp28812 : 1;
  assign tmp28835 = l2 ? 1 : tmp27488;
  assign tmp28834 = ~(l1 ? tmp27488 : tmp28835);
  assign tmp28833 = s0 ? 1 : tmp28834;
  assign tmp28831 = s1 ? tmp28832 : tmp28833;
  assign tmp28836 = s1 ? tmp28819 : 1;
  assign tmp28830 = s2 ? tmp28831 : tmp28836;
  assign tmp28822 = ~(s3 ? tmp28823 : tmp28830);
  assign tmp28805 = ~(s4 ? tmp28806 : tmp28822);
  assign tmp28769 = s5 ? tmp28770 : tmp28805;
  assign tmp28736 = s6 ? tmp28737 : tmp28769;
  assign tmp28735 = s7 ? tmp28736 : tmp27575;
  assign tmp28634 = s8 ? tmp28635 : tmp28735;
  assign tmp28843 = s0 ? tmp28740 : tmp28744;
  assign tmp28842 = s1 ? tmp28740 : tmp28843;
  assign tmp28846 = s0 ? tmp28749 : tmp27750;
  assign tmp28845 = s1 ? tmp28846 : tmp28752;
  assign tmp28844 = s2 ? tmp28746 : tmp28845;
  assign tmp28841 = s3 ? tmp28842 : tmp28844;
  assign tmp28850 = s0 ? tmp28740 : tmp27784;
  assign tmp28849 = s1 ? tmp28850 : tmp28757;
  assign tmp28852 = s0 ? tmp28740 : tmp27750;
  assign tmp28854 = l1 ? tmp27560 : tmp27971;
  assign tmp28853 = s0 ? tmp28854 : tmp27750;
  assign tmp28851 = s1 ? tmp28852 : tmp28853;
  assign tmp28848 = s2 ? tmp28849 : tmp28851;
  assign tmp28857 = s0 ? tmp28854 : tmp28740;
  assign tmp28860 = l2 ? tmp27490 : tmp27496;
  assign tmp28859 = l1 ? tmp27891 : tmp28860;
  assign tmp28858 = s0 ? tmp27750 : tmp28859;
  assign tmp28856 = s1 ? tmp28857 : tmp28858;
  assign tmp28863 = l1 ? 1 : tmp28641;
  assign tmp28862 = s0 ? tmp28863 : tmp28644;
  assign tmp28861 = s1 ? tmp28767 : tmp28862;
  assign tmp28855 = s2 ? tmp28856 : tmp28861;
  assign tmp28847 = s3 ? tmp28848 : tmp28855;
  assign tmp28840 = s4 ? tmp28841 : tmp28847;
  assign tmp28869 = s0 ? tmp28744 : tmp27750;
  assign tmp28870 = s0 ? tmp27750 : tmp27560;
  assign tmp28868 = s1 ? tmp28869 : tmp28870;
  assign tmp28872 = s0 ? tmp27750 : tmp28778;
  assign tmp28873 = s0 ? tmp28768 : tmp27750;
  assign tmp28871 = s1 ? tmp28872 : tmp28873;
  assign tmp28867 = s2 ? tmp28868 : tmp28871;
  assign tmp28876 = s0 ? tmp27750 : tmp28749;
  assign tmp28877 = s0 ? tmp27750 : tmp28785;
  assign tmp28875 = s1 ? tmp28876 : tmp28877;
  assign tmp28879 = s0 ? tmp28863 : tmp27750;
  assign tmp28878 = s1 ? tmp28879 : tmp28787;
  assign tmp28874 = s2 ? tmp28875 : tmp28878;
  assign tmp28866 = s3 ? tmp28867 : tmp28874;
  assign tmp28884 = l1 ? 1 : tmp28860;
  assign tmp28883 = s0 ? tmp28884 : tmp28778;
  assign tmp28885 = s0 ? tmp27784 : tmp28014;
  assign tmp28882 = s1 ? tmp28883 : tmp28885;
  assign tmp28887 = s0 ? tmp28795 : tmp27784;
  assign tmp28886 = s1 ? tmp28885 : tmp28887;
  assign tmp28881 = s2 ? tmp28882 : tmp28886;
  assign tmp28890 = s0 ? tmp28859 : tmp27750;
  assign tmp28889 = s1 ? tmp27750 : tmp28890;
  assign tmp28888 = s2 ? tmp28797 : tmp28889;
  assign tmp28880 = s3 ? tmp28881 : tmp28888;
  assign tmp28865 = s4 ? tmp28866 : tmp28880;
  assign tmp28895 = s0 ? tmp28810 : tmp27791;
  assign tmp28897 = l1 ? 1 : tmp27971;
  assign tmp28896 = ~(s0 ? tmp27750 : tmp28897);
  assign tmp28894 = s1 ? tmp28895 : tmp28896;
  assign tmp28899 = s0 ? tmp28897 : tmp27504;
  assign tmp28898 = ~(s1 ? tmp28899 : tmp28815);
  assign tmp28893 = s2 ? tmp28894 : tmp28898;
  assign tmp28902 = s0 ? tmp27697 : tmp27750;
  assign tmp28901 = s1 ? tmp28902 : tmp27750;
  assign tmp28905 = l1 ? 1 : tmp27739;
  assign tmp28904 = s0 ? tmp27750 : tmp28905;
  assign tmp28906 = s0 ? tmp28905 : tmp28820;
  assign tmp28903 = s1 ? tmp28904 : tmp28906;
  assign tmp28900 = ~(s2 ? tmp28901 : tmp28903);
  assign tmp28892 = s3 ? tmp28893 : tmp28900;
  assign tmp28910 = s0 ? tmp28820 : tmp27750;
  assign tmp28911 = s0 ? tmp27750 : tmp28863;
  assign tmp28909 = s1 ? tmp28910 : tmp28911;
  assign tmp28913 = s0 ? tmp27750 : tmp28828;
  assign tmp28912 = s1 ? tmp28913 : tmp28829;
  assign tmp28908 = s2 ? tmp28909 : tmp28912;
  assign tmp28916 = s0 ? tmp28897 : tmp27750;
  assign tmp28917 = s0 ? tmp27750 : tmp28834;
  assign tmp28915 = s1 ? tmp28916 : tmp28917;
  assign tmp28918 = s1 ? tmp28906 : tmp27750;
  assign tmp28914 = s2 ? tmp28915 : tmp28918;
  assign tmp28907 = ~(s3 ? tmp28908 : tmp28914);
  assign tmp28891 = ~(s4 ? tmp28892 : tmp28907);
  assign tmp28864 = s5 ? tmp28865 : tmp28891;
  assign tmp28839 = s6 ? tmp28840 : tmp28864;
  assign tmp28838 = s7 ? tmp28839 : tmp27575;
  assign tmp28837 = s8 ? tmp28735 : tmp28838;
  assign tmp28633 = s9 ? tmp28634 : tmp28837;
  assign tmp28920 = s8 ? tmp28735 : tmp28736;
  assign tmp28919 = s9 ? tmp28920 : tmp27575;
  assign tmp28632 = s10 ? tmp28633 : tmp28919;
  assign tmp28427 = s12 ? tmp28428 : tmp28632;
  assign tmp28930 = l1 ? tmp28643 : tmp27489;
  assign tmp28932 = l1 ? tmp28643 : tmp27820;
  assign tmp28934 = l2 ? tmp27496 : tmp27491;
  assign tmp28933 = ~(l1 ? tmp28934 : tmp27521);
  assign tmp28931 = s0 ? tmp28932 : tmp28933;
  assign tmp28929 = s1 ? tmp28930 : tmp28931;
  assign tmp28938 = l2 ? tmp27496 : tmp27506;
  assign tmp28939 = ~(l1 ? tmp28641 : tmp27729);
  assign tmp28937 = s0 ? tmp28938 : tmp28939;
  assign tmp28941 = l1 ? tmp28938 : tmp27624;
  assign tmp28940 = s0 ? tmp28941 : tmp28939;
  assign tmp28936 = s1 ? tmp28937 : tmp28940;
  assign tmp28943 = s0 ? tmp28941 : tmp27517;
  assign tmp28945 = l1 ? tmp28641 : tmp27729;
  assign tmp28946 = l1 ? tmp28641 : tmp27489;
  assign tmp28944 = ~(s0 ? tmp28945 : tmp28946);
  assign tmp28942 = s1 ? tmp28943 : tmp28944;
  assign tmp28935 = ~(s2 ? tmp28936 : tmp28942);
  assign tmp28928 = s3 ? tmp28929 : tmp28935;
  assign tmp28951 = l1 ? tmp28938 : tmp27521;
  assign tmp28950 = s0 ? tmp28951 : tmp28938;
  assign tmp28952 = ~(s0 ? tmp28946 : tmp28945);
  assign tmp28949 = s1 ? tmp28950 : tmp28952;
  assign tmp28954 = s0 ? tmp28930 : 1;
  assign tmp28956 = l1 ? tmp28643 : tmp27506;
  assign tmp28955 = s0 ? tmp28956 : 1;
  assign tmp28953 = ~(s1 ? tmp28954 : tmp28955);
  assign tmp28948 = s2 ? tmp28949 : tmp28953;
  assign tmp28959 = s0 ? tmp28956 : tmp28932;
  assign tmp28958 = s1 ? tmp28959 : 1;
  assign tmp28962 = l1 ? tmp28678 : tmp27729;
  assign tmp28961 = s0 ? tmp28945 : tmp28962;
  assign tmp28964 = l1 ? tmp28661 : 1;
  assign tmp28963 = s0 ? tmp28964 : tmp28945;
  assign tmp28960 = s1 ? tmp28961 : tmp28963;
  assign tmp28957 = ~(s2 ? tmp28958 : tmp28960);
  assign tmp28947 = ~(s3 ? tmp28948 : tmp28957);
  assign tmp28927 = s4 ? tmp28928 : tmp28947;
  assign tmp28971 = l1 ? tmp28934 : tmp27521;
  assign tmp28970 = s0 ? tmp28971 : tmp27517;
  assign tmp28969 = s1 ? tmp28970 : tmp28938;
  assign tmp28974 = l1 ? tmp28934 : tmp28080;
  assign tmp28973 = s0 ? tmp27517 : tmp28974;
  assign tmp28975 = ~(s0 ? tmp28962 : tmp27960);
  assign tmp28972 = s1 ? tmp28973 : tmp28975;
  assign tmp28968 = s2 ? tmp28969 : tmp28972;
  assign tmp28978 = s0 ? tmp27517 : tmp28941;
  assign tmp28980 = ~(l1 ? tmp28678 : tmp27563);
  assign tmp28979 = s0 ? tmp27517 : tmp28980;
  assign tmp28977 = s1 ? tmp28978 : tmp28979;
  assign tmp28982 = s0 ? tmp28964 : 1;
  assign tmp28984 = l1 ? tmp28641 : tmp27563;
  assign tmp28985 = l1 ? tmp28678 : tmp27563;
  assign tmp28983 = s0 ? tmp28984 : tmp28985;
  assign tmp28981 = ~(s1 ? tmp28982 : tmp28983);
  assign tmp28976 = s2 ? tmp28977 : tmp28981;
  assign tmp28967 = s3 ? tmp28968 : tmp28976;
  assign tmp28990 = l1 ? tmp28641 : tmp27684;
  assign tmp28989 = s0 ? 1 : tmp28990;
  assign tmp28992 = l1 ? tmp28643 : tmp27575;
  assign tmp28991 = s0 ? tmp28992 : tmp27530;
  assign tmp28988 = s1 ? tmp28989 : tmp28991;
  assign tmp28995 = l1 ? tmp28938 : tmp28080;
  assign tmp28996 = ~(l1 ? tmp28643 : tmp27575);
  assign tmp28994 = ~(s0 ? tmp28995 : tmp28996);
  assign tmp28993 = s1 ? tmp28991 : tmp28994;
  assign tmp28987 = s2 ? tmp28988 : tmp28993;
  assign tmp29000 = l1 ? tmp27495 : tmp28080;
  assign tmp29001 = ~(l1 ? tmp28643 : tmp27499);
  assign tmp28999 = s0 ? tmp29000 : tmp29001;
  assign tmp29002 = s0 ? tmp27533 : tmp28980;
  assign tmp28998 = s1 ? tmp28999 : tmp29002;
  assign tmp28997 = ~(s2 ? tmp28998 : 0);
  assign tmp28986 = ~(s3 ? tmp28987 : tmp28997);
  assign tmp28966 = s4 ? tmp28967 : tmp28986;
  assign tmp29007 = s0 ? tmp28985 : 1;
  assign tmp29009 = ~(l1 ? tmp27517 : 0);
  assign tmp29008 = s0 ? 1 : tmp29009;
  assign tmp29006 = s1 ? tmp29007 : tmp29008;
  assign tmp29012 = l1 ? tmp27517 : 0;
  assign tmp29011 = s0 ? tmp29012 : tmp27495;
  assign tmp29010 = ~(s1 ? tmp29011 : tmp27495);
  assign tmp29005 = s2 ? tmp29006 : tmp29010;
  assign tmp29014 = s1 ? tmp27917 : 0;
  assign tmp29017 = ~(l1 ? tmp27495 : tmp27508);
  assign tmp29016 = s0 ? 1 : tmp29017;
  assign tmp29015 = ~(s1 ? 1 : tmp29016);
  assign tmp29013 = ~(s2 ? tmp29014 : tmp29015);
  assign tmp29004 = s3 ? tmp29005 : tmp29013;
  assign tmp29022 = l1 ? tmp27495 : tmp27508;
  assign tmp29021 = s0 ? tmp29022 : tmp29012;
  assign tmp29024 = ~(l1 ? tmp28661 : 1);
  assign tmp29023 = s0 ? tmp29012 : tmp29024;
  assign tmp29020 = s1 ? tmp29021 : tmp29023;
  assign tmp29027 = ~(l1 ? tmp28733 : tmp28080);
  assign tmp29026 = s0 ? 1 : tmp29027;
  assign tmp29025 = ~(s1 ? tmp29026 : tmp27575);
  assign tmp29019 = s2 ? tmp29020 : tmp29025;
  assign tmp29031 = l1 ? tmp28678 : tmp27499;
  assign tmp29030 = ~(s0 ? 1 : tmp29031);
  assign tmp29029 = s1 ? tmp29012 : tmp29030;
  assign tmp29032 = ~(s1 ? tmp29016 : tmp29008);
  assign tmp29028 = s2 ? tmp29029 : tmp29032;
  assign tmp29018 = ~(s3 ? tmp29019 : tmp29028);
  assign tmp29003 = ~(s4 ? tmp29004 : tmp29018);
  assign tmp28965 = ~(s5 ? tmp28966 : tmp29003);
  assign tmp28926 = s6 ? tmp28927 : tmp28965;
  assign tmp28925 = s7 ? tmp28926 : tmp27575;
  assign tmp29038 = l1 ? tmp28643 : tmp28608;
  assign tmp29040 = l1 ? tmp27560 : tmp28525;
  assign tmp29041 = l1 ? tmp28741 : tmp28608;
  assign tmp29039 = s0 ? tmp29040 : tmp29041;
  assign tmp29037 = s1 ? tmp29038 : tmp29039;
  assign tmp29045 = l1 ? tmp28641 : tmp28614;
  assign tmp29044 = s0 ? tmp28263 : tmp29045;
  assign tmp29048 = ~(l2 ? tmp27554 : tmp27506);
  assign tmp29047 = l1 ? tmp27980 : tmp29048;
  assign tmp29046 = s0 ? tmp29047 : tmp29045;
  assign tmp29043 = s1 ? tmp29044 : tmp29046;
  assign tmp29050 = s0 ? tmp29047 : tmp28267;
  assign tmp29052 = l1 ? tmp28641 : tmp28608;
  assign tmp29051 = s0 ? tmp29045 : tmp29052;
  assign tmp29049 = s1 ? tmp29050 : tmp29051;
  assign tmp29042 = s2 ? tmp29043 : tmp29049;
  assign tmp29036 = s3 ? tmp29037 : tmp29042;
  assign tmp29057 = l1 ? tmp27980 : tmp28608;
  assign tmp29056 = s0 ? tmp29057 : tmp28258;
  assign tmp29058 = s0 ? tmp29052 : tmp29045;
  assign tmp29055 = s1 ? tmp29056 : tmp29058;
  assign tmp29060 = s0 ? tmp29038 : 1;
  assign tmp29062 = l1 ? tmp27560 : tmp28324;
  assign tmp29061 = s0 ? tmp29062 : 1;
  assign tmp29059 = s1 ? tmp29060 : tmp29061;
  assign tmp29054 = s2 ? tmp29055 : tmp29059;
  assign tmp29065 = s0 ? tmp29062 : tmp29040;
  assign tmp29064 = s1 ? tmp29065 : 1;
  assign tmp29068 = l1 ? tmp28678 : tmp28614;
  assign tmp29067 = s0 ? tmp29045 : tmp29068;
  assign tmp29070 = l1 ? tmp27891 : tmp27492;
  assign tmp29069 = s0 ? tmp29070 : tmp29045;
  assign tmp29066 = s1 ? tmp29067 : tmp29069;
  assign tmp29063 = s2 ? tmp29064 : tmp29066;
  assign tmp29053 = s3 ? tmp29054 : tmp29063;
  assign tmp29035 = s4 ? tmp29036 : tmp29053;
  assign tmp29076 = s0 ? tmp29041 : tmp27833;
  assign tmp29078 = ~(l1 ? tmp27980 : tmp28226);
  assign tmp29077 = ~(s0 ? tmp27504 : tmp29078);
  assign tmp29075 = s1 ? tmp29076 : tmp29077;
  assign tmp29081 = ~(l1 ? tmp28741 : tmp28324);
  assign tmp29080 = s0 ? tmp27504 : tmp29081;
  assign tmp29082 = ~(s0 ? tmp29068 : tmp28267);
  assign tmp29079 = ~(s1 ? tmp29080 : tmp29082);
  assign tmp29074 = s2 ? tmp29075 : tmp29079;
  assign tmp29085 = s0 ? tmp28267 : tmp29047;
  assign tmp29088 = l2 ? tmp27490 : tmp27492;
  assign tmp29087 = l1 ? tmp29088 : tmp27492;
  assign tmp29086 = s0 ? tmp28267 : tmp29087;
  assign tmp29084 = s1 ? tmp29085 : tmp29086;
  assign tmp29090 = s0 ? tmp29070 : 1;
  assign tmp29092 = l1 ? tmp28641 : tmp27492;
  assign tmp29093 = l1 ? tmp28678 : tmp27492;
  assign tmp29091 = s0 ? tmp29092 : tmp29093;
  assign tmp29089 = s1 ? tmp29090 : tmp29091;
  assign tmp29083 = s2 ? tmp29084 : tmp29089;
  assign tmp29073 = s3 ? tmp29074 : tmp29083;
  assign tmp29098 = l1 ? tmp28641 : tmp28570;
  assign tmp29097 = s0 ? 1 : tmp29098;
  assign tmp29099 = s0 ? tmp28275 : tmp27703;
  assign tmp29096 = s1 ? tmp29097 : tmp29099;
  assign tmp29102 = l1 ? tmp27980 : tmp28324;
  assign tmp29101 = s0 ? tmp29102 : tmp28275;
  assign tmp29100 = s1 ? tmp29099 : tmp29101;
  assign tmp29095 = s2 ? tmp29096 : tmp29100;
  assign tmp29106 = l1 ? 1 : tmp27554;
  assign tmp29107 = ~(l1 ? tmp28643 : tmp27492);
  assign tmp29105 = s0 ? tmp29106 : tmp29107;
  assign tmp29108 = ~(s0 ? tmp27703 : tmp29087);
  assign tmp29104 = s1 ? tmp29105 : tmp29108;
  assign tmp29103 = ~(s2 ? tmp29104 : 0);
  assign tmp29094 = s3 ? tmp29095 : tmp29103;
  assign tmp29072 = s4 ? tmp29073 : tmp29094;
  assign tmp29113 = s0 ? tmp29087 : 1;
  assign tmp29115 = ~(l1 ? tmp27504 : tmp27488);
  assign tmp29114 = s0 ? 1 : tmp29115;
  assign tmp29112 = s1 ? tmp29113 : tmp29114;
  assign tmp29118 = l1 ? tmp27504 : tmp27488;
  assign tmp29117 = s0 ? tmp29118 : 1;
  assign tmp29116 = ~(s1 ? tmp29117 : 1);
  assign tmp29111 = s2 ? tmp29112 : tmp29116;
  assign tmp29120 = s1 ? tmp27999 : 0;
  assign tmp29123 = ~(l1 ? 1 : tmp27488);
  assign tmp29122 = s0 ? 1 : tmp29123;
  assign tmp29121 = ~(s1 ? 1 : tmp29122);
  assign tmp29119 = ~(s2 ? tmp29120 : tmp29121);
  assign tmp29110 = s3 ? tmp29111 : tmp29119;
  assign tmp29127 = s0 ? tmp28812 : tmp27697;
  assign tmp29129 = ~(l1 ? tmp27891 : tmp27492);
  assign tmp29128 = s0 ? tmp27697 : tmp29129;
  assign tmp29126 = s1 ? tmp29127 : tmp29128;
  assign tmp29132 = ~(l1 ? tmp28835 : tmp27554);
  assign tmp29131 = s0 ? 1 : tmp29132;
  assign tmp29130 = ~(s1 ? tmp29131 : 0);
  assign tmp29125 = s2 ? tmp29126 : tmp29130;
  assign tmp29135 = s0 ? tmp29118 : tmp27697;
  assign tmp29137 = l1 ? tmp29088 : tmp27499;
  assign tmp29136 = ~(s0 ? 1 : tmp29137);
  assign tmp29134 = s1 ? tmp29135 : tmp29136;
  assign tmp29139 = s0 ? 1 : tmp28081;
  assign tmp29138 = ~(s1 ? tmp29122 : tmp29139);
  assign tmp29133 = s2 ? tmp29134 : tmp29138;
  assign tmp29124 = ~(s3 ? tmp29125 : tmp29133);
  assign tmp29109 = s4 ? tmp29110 : tmp29124;
  assign tmp29071 = s5 ? tmp29072 : tmp29109;
  assign tmp29034 = s6 ? tmp29035 : tmp29071;
  assign tmp29033 = s7 ? tmp29034 : tmp27575;
  assign tmp28924 = s8 ? tmp28925 : tmp29033;
  assign tmp29147 = l1 ? tmp28741 : tmp27489;
  assign tmp29146 = s0 ? tmp27771 : tmp29147;
  assign tmp29145 = s1 ? tmp28930 : tmp29146;
  assign tmp29151 = l1 ? tmp27980 : tmp27489;
  assign tmp29150 = ~(s0 ? tmp29151 : tmp28945);
  assign tmp29149 = s1 ? tmp28937 : tmp29150;
  assign tmp29154 = ~(l1 ? tmp27497 : tmp27521);
  assign tmp29153 = s0 ? tmp29151 : tmp29154;
  assign tmp29155 = s0 ? tmp28945 : tmp28946;
  assign tmp29152 = ~(s1 ? tmp29153 : tmp29155);
  assign tmp29148 = ~(s2 ? tmp29149 : tmp29152);
  assign tmp29144 = s3 ? tmp29145 : tmp29148;
  assign tmp29160 = l1 ? tmp27560 : tmp27739;
  assign tmp29159 = s0 ? tmp29151 : tmp29160;
  assign tmp29161 = s0 ? tmp28946 : tmp28945;
  assign tmp29158 = s1 ? tmp29159 : tmp29161;
  assign tmp29163 = s0 ? tmp28930 : tmp27750;
  assign tmp29165 = l1 ? tmp27560 : tmp27553;
  assign tmp29164 = s0 ? tmp29165 : tmp27750;
  assign tmp29162 = s1 ? tmp29163 : tmp29164;
  assign tmp29157 = s2 ? tmp29158 : tmp29162;
  assign tmp29168 = s0 ? tmp29165 : tmp27771;
  assign tmp29167 = s1 ? tmp29168 : tmp27750;
  assign tmp29171 = l1 ? tmp27891 : tmp27744;
  assign tmp29170 = s0 ? tmp29171 : tmp28945;
  assign tmp29169 = s1 ? tmp28961 : tmp29170;
  assign tmp29166 = s2 ? tmp29167 : tmp29169;
  assign tmp29156 = s3 ? tmp29157 : tmp29166;
  assign tmp29143 = s4 ? tmp29144 : tmp29156;
  assign tmp29178 = ~(l1 ? tmp27504 : tmp27760);
  assign tmp29177 = s0 ? tmp29147 : tmp29178;
  assign tmp29180 = l1 ? tmp27504 : tmp27760;
  assign tmp29179 = ~(s0 ? tmp29180 : tmp28938);
  assign tmp29176 = s1 ? tmp29177 : tmp29179;
  assign tmp29183 = ~(l1 ? tmp28741 : tmp27489);
  assign tmp29182 = s0 ? tmp29180 : tmp29183;
  assign tmp29184 = ~(s0 ? tmp28962 : tmp27767);
  assign tmp29181 = ~(s1 ? tmp29182 : tmp29184);
  assign tmp29175 = s2 ? tmp29176 : tmp29181;
  assign tmp29187 = s0 ? tmp27767 : tmp29151;
  assign tmp29189 = l1 ? tmp29088 : tmp27729;
  assign tmp29188 = s0 ? tmp27767 : tmp29189;
  assign tmp29186 = s1 ? tmp29187 : tmp29188;
  assign tmp29191 = s0 ? tmp29171 : tmp27750;
  assign tmp29193 = l1 ? tmp28678 : tmp27744;
  assign tmp29192 = s0 ? tmp28945 : tmp29193;
  assign tmp29190 = s1 ? tmp29191 : tmp29192;
  assign tmp29185 = s2 ? tmp29186 : tmp29190;
  assign tmp29174 = s3 ? tmp29175 : tmp29185;
  assign tmp29197 = s0 ? tmp27750 : tmp28946;
  assign tmp29198 = s0 ? tmp28275 : tmp27743;
  assign tmp29196 = s1 ? tmp29197 : tmp29198;
  assign tmp29200 = s0 ? tmp29151 : tmp28275;
  assign tmp29199 = s1 ? tmp29198 : tmp29200;
  assign tmp29195 = s2 ? tmp29196 : tmp29199;
  assign tmp29204 = l1 ? 1 : tmp27521;
  assign tmp29205 = ~(l1 ? tmp28643 : tmp27744);
  assign tmp29203 = s0 ? tmp29204 : tmp29205;
  assign tmp29207 = l1 ? tmp29088 : tmp27744;
  assign tmp29206 = ~(s0 ? tmp27743 : tmp29207);
  assign tmp29202 = s1 ? tmp29203 : tmp29206;
  assign tmp29201 = ~(s2 ? tmp29202 : tmp27791);
  assign tmp29194 = s3 ? tmp29195 : tmp29201;
  assign tmp29173 = s4 ? tmp29174 : tmp29194;
  assign tmp29212 = s0 ? tmp29189 : tmp27750;
  assign tmp29214 = ~(l1 ? tmp27504 : tmp27809);
  assign tmp29213 = s0 ? tmp27750 : tmp29214;
  assign tmp29211 = s1 ? tmp29212 : tmp29213;
  assign tmp29217 = l1 ? tmp27504 : tmp27809;
  assign tmp29218 = l1 ? 1 : tmp28080;
  assign tmp29216 = s0 ? tmp29217 : tmp29218;
  assign tmp29219 = s0 ? 1 : tmp29218;
  assign tmp29215 = ~(s1 ? tmp29216 : tmp29219);
  assign tmp29210 = s2 ? tmp29211 : tmp29215;
  assign tmp29222 = s0 ? 1 : tmp27791;
  assign tmp29221 = s1 ? tmp29222 : tmp27791;
  assign tmp29225 = ~(l1 ? 1 : tmp27809);
  assign tmp29224 = s0 ? tmp27750 : tmp29225;
  assign tmp29223 = ~(s1 ? tmp27750 : tmp29224);
  assign tmp29220 = ~(s2 ? tmp29221 : tmp29223);
  assign tmp29209 = s3 ? tmp29210 : tmp29220;
  assign tmp29230 = l1 ? 1 : tmp27809;
  assign tmp29229 = s0 ? tmp29230 : tmp29217;
  assign tmp29232 = ~(l1 ? tmp27891 : tmp27744);
  assign tmp29231 = s0 ? tmp29217 : tmp29232;
  assign tmp29228 = s1 ? tmp29229 : tmp29231;
  assign tmp29235 = ~(l1 ? tmp28835 : tmp27521);
  assign tmp29234 = s0 ? tmp27750 : tmp29235;
  assign tmp29236 = ~(s0 ? tmp29218 : 1);
  assign tmp29233 = ~(s1 ? tmp29234 : tmp29236);
  assign tmp29227 = s2 ? tmp29228 : tmp29233;
  assign tmp29239 = ~(s0 ? tmp27750 : tmp29207);
  assign tmp29238 = s1 ? tmp29217 : tmp29239;
  assign tmp29240 = ~(s1 ? tmp29224 : tmp29213);
  assign tmp29237 = s2 ? tmp29238 : tmp29240;
  assign tmp29226 = ~(s3 ? tmp29227 : tmp29237);
  assign tmp29208 = s4 ? tmp29209 : tmp29226;
  assign tmp29172 = s5 ? tmp29173 : tmp29208;
  assign tmp29142 = s6 ? tmp29143 : tmp29172;
  assign tmp29141 = s7 ? tmp29142 : tmp27575;
  assign tmp29140 = s8 ? tmp29033 : tmp29141;
  assign tmp28923 = s9 ? tmp28924 : tmp29140;
  assign tmp29249 = l1 ? tmp27560 : tmp27820;
  assign tmp29248 = s0 ? tmp29249 : tmp29147;
  assign tmp29247 = s1 ? tmp28930 : tmp29248;
  assign tmp29253 = l1 ? tmp27980 : tmp27513;
  assign tmp29252 = ~(s0 ? tmp29253 : tmp28945);
  assign tmp29251 = s1 ? tmp28937 : tmp29252;
  assign tmp29255 = s0 ? tmp29253 : tmp27820;
  assign tmp29254 = ~(s1 ? tmp29255 : tmp29155);
  assign tmp29250 = ~(s2 ? tmp29251 : tmp29254);
  assign tmp29246 = s3 ? tmp29247 : tmp29250;
  assign tmp29259 = s0 ? tmp29151 : tmp28258;
  assign tmp29258 = s1 ? tmp29259 : tmp29161;
  assign tmp29262 = l1 ? tmp27560 : tmp27506;
  assign tmp29261 = s0 ? tmp29262 : 1;
  assign tmp29260 = s1 ? tmp28954 : tmp29261;
  assign tmp29257 = s2 ? tmp29258 : tmp29260;
  assign tmp29265 = s0 ? tmp29262 : tmp29249;
  assign tmp29264 = s1 ? tmp29265 : 1;
  assign tmp29268 = l1 ? tmp27891 : 1;
  assign tmp29267 = s0 ? tmp29268 : tmp28945;
  assign tmp29266 = s1 ? tmp28961 : tmp29267;
  assign tmp29263 = s2 ? tmp29264 : tmp29266;
  assign tmp29256 = s3 ? tmp29257 : tmp29263;
  assign tmp29245 = s4 ? tmp29246 : tmp29256;
  assign tmp29274 = s0 ? tmp29147 : tmp27833;
  assign tmp29275 = ~(s0 ? tmp27504 : tmp28938);
  assign tmp29273 = s1 ? tmp29274 : tmp29275;
  assign tmp29278 = ~(l1 ? tmp28741 : tmp27684);
  assign tmp29277 = s0 ? tmp27504 : tmp29278;
  assign tmp29279 = ~(s0 ? tmp28962 : tmp27858);
  assign tmp29276 = ~(s1 ? tmp29277 : tmp29279);
  assign tmp29272 = s2 ? tmp29273 : tmp29276;
  assign tmp29282 = s0 ? tmp27858 : tmp29253;
  assign tmp29284 = l1 ? tmp29088 : tmp27563;
  assign tmp29283 = s0 ? tmp27858 : tmp29284;
  assign tmp29281 = s1 ? tmp29282 : tmp29283;
  assign tmp29286 = s0 ? tmp29268 : 1;
  assign tmp29287 = s0 ? tmp28984 : tmp29031;
  assign tmp29285 = s1 ? tmp29286 : tmp29287;
  assign tmp29280 = s2 ? tmp29281 : tmp29285;
  assign tmp29271 = s3 ? tmp29272 : tmp29280;
  assign tmp29291 = s0 ? tmp28275 : tmp27836;
  assign tmp29290 = s1 ? tmp28989 : tmp29291;
  assign tmp29294 = l1 ? tmp27980 : tmp27684;
  assign tmp29293 = s0 ? tmp29294 : tmp28275;
  assign tmp29292 = s1 ? tmp29291 : tmp29293;
  assign tmp29289 = s2 ? tmp29290 : tmp29292;
  assign tmp29298 = l1 ? 1 : tmp27569;
  assign tmp29297 = s0 ? tmp29298 : tmp29001;
  assign tmp29299 = ~(s0 ? tmp27836 : tmp29087);
  assign tmp29296 = s1 ? tmp29297 : tmp29299;
  assign tmp29295 = ~(s2 ? tmp29296 : 0);
  assign tmp29288 = s3 ? tmp29289 : tmp29295;
  assign tmp29270 = s4 ? tmp29271 : tmp29288;
  assign tmp29304 = s0 ? tmp29284 : 1;
  assign tmp29303 = s1 ? tmp29304 : tmp29139;
  assign tmp29306 = s0 ? tmp27697 : tmp27985;
  assign tmp29307 = s0 ? 1 : tmp27985;
  assign tmp29305 = ~(s1 ? tmp29306 : tmp29307);
  assign tmp29302 = s2 ? tmp29303 : tmp29305;
  assign tmp29301 = s3 ? tmp29302 : tmp29119;
  assign tmp29312 = ~(l1 ? tmp27891 : 1);
  assign tmp29311 = s0 ? tmp27697 : tmp29312;
  assign tmp29310 = s1 ? tmp29127 : tmp29311;
  assign tmp29315 = ~(l1 ? tmp28835 : tmp27569);
  assign tmp29314 = s0 ? 1 : tmp29315;
  assign tmp29316 = ~(s0 ? tmp27985 : 1);
  assign tmp29313 = ~(s1 ? tmp29314 : tmp29316);
  assign tmp29309 = s2 ? tmp29310 : tmp29313;
  assign tmp29318 = s1 ? tmp27697 : tmp29136;
  assign tmp29317 = s2 ? tmp29318 : tmp29138;
  assign tmp29308 = ~(s3 ? tmp29309 : tmp29317);
  assign tmp29300 = s4 ? tmp29301 : tmp29308;
  assign tmp29269 = s5 ? tmp29270 : tmp29300;
  assign tmp29244 = s6 ? tmp29245 : tmp29269;
  assign tmp29243 = s7 ? tmp29244 : tmp27575;
  assign tmp29242 = s8 ? tmp29243 : tmp29244;
  assign tmp29241 = s9 ? tmp29242 : tmp27575;
  assign tmp28922 = s10 ? tmp28923 : tmp29241;
  assign tmp29327 = l1 ? tmp28643 : tmp27744;
  assign tmp29329 = ~(l1 ? tmp28934 : tmp27809);
  assign tmp29328 = s0 ? tmp28654 : tmp29329;
  assign tmp29326 = s1 ? tmp29327 : tmp29328;
  assign tmp29333 = l1 ? tmp28938 : tmp28490;
  assign tmp29334 = ~(l1 ? tmp28641 : tmp27744);
  assign tmp29332 = s0 ? tmp29333 : tmp29334;
  assign tmp29336 = l1 ? tmp28938 : tmp28495;
  assign tmp29335 = s0 ? tmp29336 : tmp29334;
  assign tmp29331 = s1 ? tmp29332 : tmp29335;
  assign tmp29338 = s0 ? tmp29336 : 0;
  assign tmp29337 = s1 ? tmp29338 : tmp29334;
  assign tmp29330 = ~(s2 ? tmp29331 : tmp29337);
  assign tmp29325 = s3 ? tmp29326 : tmp29330;
  assign tmp29343 = l1 ? tmp28938 : tmp27809;
  assign tmp29344 = ~(l1 ? tmp28643 : 1);
  assign tmp29342 = s0 ? tmp29343 : tmp29344;
  assign tmp29341 = s1 ? tmp29342 : tmp29334;
  assign tmp29346 = s0 ? tmp29327 : 1;
  assign tmp29347 = s0 ? tmp28654 : 1;
  assign tmp29345 = ~(s1 ? tmp29346 : tmp29347);
  assign tmp29340 = s2 ? tmp29341 : tmp29345;
  assign tmp29349 = s1 ? tmp28654 : 1;
  assign tmp29352 = l1 ? tmp28641 : tmp27744;
  assign tmp29351 = s0 ? tmp29352 : tmp29193;
  assign tmp29353 = s0 ? tmp28964 : tmp29352;
  assign tmp29350 = s1 ? tmp29351 : tmp29353;
  assign tmp29348 = ~(s2 ? tmp29349 : tmp29350);
  assign tmp29339 = ~(s3 ? tmp29340 : tmp29348);
  assign tmp29324 = s4 ? tmp29325 : tmp29339;
  assign tmp29360 = l1 ? tmp28934 : tmp27809;
  assign tmp29359 = s0 ? tmp29360 : 0;
  assign tmp29358 = s1 ? tmp29359 : tmp29333;
  assign tmp29363 = ~(l1 ? tmp28934 : tmp27606);
  assign tmp29362 = s0 ? 1 : tmp29363;
  assign tmp29364 = s0 ? tmp29193 : 1;
  assign tmp29361 = ~(s1 ? tmp29362 : tmp29364);
  assign tmp29357 = s2 ? tmp29358 : tmp29361;
  assign tmp29368 = ~(l1 ? tmp28938 : tmp28495);
  assign tmp29367 = s0 ? 1 : tmp29368;
  assign tmp29369 = s0 ? 1 : tmp29031;
  assign tmp29366 = s1 ? tmp29367 : tmp29369;
  assign tmp29372 = l1 ? tmp28641 : tmp27499;
  assign tmp29371 = s0 ? tmp29372 : tmp28985;
  assign tmp29370 = s1 ? tmp28982 : tmp29371;
  assign tmp29365 = ~(s2 ? tmp29366 : tmp29370);
  assign tmp29356 = s3 ? tmp29357 : tmp29365;
  assign tmp29376 = s0 ? 1 : tmp29372;
  assign tmp29377 = s0 ? tmp28654 : tmp27530;
  assign tmp29375 = s1 ? tmp29376 : tmp29377;
  assign tmp29380 = l1 ? tmp28938 : tmp27606;
  assign tmp29379 = ~(s0 ? tmp29380 : tmp29344);
  assign tmp29378 = s1 ? tmp29377 : tmp29379;
  assign tmp29374 = s2 ? tmp29375 : tmp29378;
  assign tmp29384 = l1 ? tmp27495 : tmp27606;
  assign tmp29383 = s0 ? tmp29384 : tmp29001;
  assign tmp29382 = s1 ? tmp29383 : tmp29002;
  assign tmp29381 = ~(s2 ? tmp29382 : 0);
  assign tmp29373 = ~(s3 ? tmp29374 : tmp29381);
  assign tmp29355 = s4 ? tmp29356 : tmp29373;
  assign tmp29389 = s0 ? tmp29031 : 1;
  assign tmp29388 = s1 ? tmp29389 : tmp29008;
  assign tmp29391 = s0 ? tmp29012 : tmp28225;
  assign tmp29392 = s0 ? tmp27495 : tmp28225;
  assign tmp29390 = ~(s1 ? tmp29391 : tmp29392);
  assign tmp29387 = s2 ? tmp29388 : tmp29390;
  assign tmp29386 = s3 ? tmp29387 : tmp29013;
  assign tmp29397 = ~(l1 ? tmp28733 : tmp27606);
  assign tmp29396 = s0 ? 1 : tmp29397;
  assign tmp29398 = ~(s0 ? tmp28225 : tmp27495);
  assign tmp29395 = ~(s1 ? tmp29396 : tmp29398);
  assign tmp29394 = s2 ? tmp29020 : tmp29395;
  assign tmp29393 = ~(s3 ? tmp29394 : tmp29028);
  assign tmp29385 = ~(s4 ? tmp29386 : tmp29393);
  assign tmp29354 = ~(s5 ? tmp29355 : tmp29385);
  assign tmp29323 = s6 ? tmp29324 : tmp29354;
  assign tmp29322 = s7 ? tmp29323 : tmp27575;
  assign tmp29404 = l1 ? tmp28643 : tmp27496;
  assign tmp29406 = l1 ? tmp27560 : tmp27495;
  assign tmp29407 = l1 ? tmp28741 : tmp27496;
  assign tmp29405 = s0 ? tmp29406 : tmp29407;
  assign tmp29403 = s1 ? tmp29404 : tmp29405;
  assign tmp29411 = l1 ? tmp28641 : tmp27496;
  assign tmp29410 = s0 ? tmp27979 : tmp29411;
  assign tmp29414 = l2 ? tmp27496 : tmp27490;
  assign tmp29413 = l1 ? tmp27980 : tmp29414;
  assign tmp29412 = s0 ? tmp29413 : tmp29411;
  assign tmp29409 = s1 ? tmp29410 : tmp29412;
  assign tmp29416 = s0 ? tmp29413 : tmp27642;
  assign tmp29415 = s1 ? tmp29416 : tmp29411;
  assign tmp29408 = s2 ? tmp29409 : tmp29415;
  assign tmp29402 = s3 ? tmp29403 : tmp29408;
  assign tmp29421 = l1 ? tmp27980 : tmp27496;
  assign tmp29420 = s0 ? tmp29421 : tmp27991;
  assign tmp29419 = s1 ? tmp29420 : tmp29411;
  assign tmp29423 = s0 ? tmp29404 : 1;
  assign tmp29425 = l1 ? tmp27560 : tmp27496;
  assign tmp29424 = s0 ? tmp29425 : 1;
  assign tmp29422 = s1 ? tmp29423 : tmp29424;
  assign tmp29418 = s2 ? tmp29419 : tmp29422;
  assign tmp29428 = s0 ? tmp29425 : tmp29406;
  assign tmp29427 = s1 ? tmp29428 : 1;
  assign tmp29431 = l1 ? tmp28678 : tmp27496;
  assign tmp29430 = s0 ? tmp29411 : tmp29431;
  assign tmp29432 = s0 ? tmp29070 : tmp29411;
  assign tmp29429 = s1 ? tmp29430 : tmp29432;
  assign tmp29426 = s2 ? tmp29427 : tmp29429;
  assign tmp29417 = s3 ? tmp29418 : tmp29426;
  assign tmp29401 = s4 ? tmp29402 : tmp29417;
  assign tmp29438 = s0 ? tmp29407 : 1;
  assign tmp29437 = s1 ? tmp29438 : tmp28009;
  assign tmp29442 = l2 ? tmp27496 : tmp27492;
  assign tmp29441 = l1 ? tmp28741 : tmp29442;
  assign tmp29440 = s0 ? 1 : tmp29441;
  assign tmp29443 = s0 ? tmp29431 : tmp27642;
  assign tmp29439 = s1 ? tmp29440 : tmp29443;
  assign tmp29436 = s2 ? tmp29437 : tmp29439;
  assign tmp29446 = s0 ? tmp27642 : tmp29413;
  assign tmp29448 = l1 ? tmp29088 : tmp29442;
  assign tmp29447 = s0 ? tmp27642 : tmp29448;
  assign tmp29445 = s1 ? tmp29446 : tmp29447;
  assign tmp29451 = l1 ? tmp28641 : tmp29442;
  assign tmp29450 = s0 ? tmp29451 : tmp29093;
  assign tmp29449 = s1 ? tmp29090 : tmp29450;
  assign tmp29444 = s2 ? tmp29445 : tmp29449;
  assign tmp29435 = s3 ? tmp29436 : tmp29444;
  assign tmp29455 = s0 ? 1 : tmp29451;
  assign tmp29456 = s0 ? tmp27991 : tmp27703;
  assign tmp29454 = s1 ? tmp29455 : tmp29456;
  assign tmp29459 = l1 ? tmp27980 : tmp29442;
  assign tmp29458 = s0 ? tmp29459 : tmp27991;
  assign tmp29457 = s1 ? tmp29456 : tmp29458;
  assign tmp29453 = s2 ? tmp29454 : tmp29457;
  assign tmp29464 = ~(l2 ? tmp27496 : tmp27492);
  assign tmp29463 = l1 ? 1 : tmp29464;
  assign tmp29462 = s0 ? tmp29463 : tmp29107;
  assign tmp29461 = s1 ? tmp29462 : tmp29108;
  assign tmp29460 = ~(s2 ? tmp29461 : 0);
  assign tmp29452 = s3 ? tmp29453 : tmp29460;
  assign tmp29434 = s4 ? tmp29435 : tmp29452;
  assign tmp29469 = s0 ? tmp29448 : 1;
  assign tmp29468 = s1 ? tmp29469 : tmp29114;
  assign tmp29471 = s0 ? tmp29118 : tmp27858;
  assign tmp29470 = ~(s1 ? tmp29471 : tmp27964);
  assign tmp29467 = s2 ? tmp29468 : tmp29470;
  assign tmp29466 = s3 ? tmp29467 : tmp29119;
  assign tmp29476 = ~(l1 ? tmp28835 : tmp29464);
  assign tmp29475 = s0 ? 1 : tmp29476;
  assign tmp29477 = ~(s0 ? tmp27858 : 1);
  assign tmp29474 = ~(s1 ? tmp29475 : tmp29477);
  assign tmp29473 = s2 ? tmp29126 : tmp29474;
  assign tmp29472 = ~(s3 ? tmp29473 : tmp29133);
  assign tmp29465 = s4 ? tmp29466 : tmp29472;
  assign tmp29433 = s5 ? tmp29434 : tmp29465;
  assign tmp29400 = s6 ? tmp29401 : tmp29433;
  assign tmp29399 = s7 ? tmp29400 : tmp27575;
  assign tmp29321 = s8 ? tmp29322 : tmp29399;
  assign tmp29485 = l1 ? tmp28741 : tmp27744;
  assign tmp29484 = s0 ? tmp27784 : tmp29485;
  assign tmp29483 = s1 ? tmp29327 : tmp29484;
  assign tmp29488 = l1 ? tmp27980 : tmp27744;
  assign tmp29487 = s0 ? tmp29488 : tmp29352;
  assign tmp29490 = s0 ? tmp29488 : tmp27750;
  assign tmp29489 = s1 ? tmp29490 : tmp29352;
  assign tmp29486 = s2 ? tmp29487 : tmp29489;
  assign tmp29482 = s3 ? tmp29483 : tmp29486;
  assign tmp29494 = s0 ? tmp29488 : tmp27784;
  assign tmp29493 = s1 ? tmp29494 : tmp29352;
  assign tmp29496 = s0 ? tmp29327 : tmp27750;
  assign tmp29497 = s0 ? tmp27784 : tmp27750;
  assign tmp29495 = s1 ? tmp29496 : tmp29497;
  assign tmp29492 = s2 ? tmp29493 : tmp29495;
  assign tmp29499 = s1 ? tmp27784 : tmp27750;
  assign tmp29501 = s0 ? tmp29171 : tmp29352;
  assign tmp29500 = s1 ? tmp29351 : tmp29501;
  assign tmp29498 = s2 ? tmp29499 : tmp29500;
  assign tmp29491 = s3 ? tmp29492 : tmp29498;
  assign tmp29481 = s4 ? tmp29482 : tmp29491;
  assign tmp29507 = s0 ? tmp29485 : tmp27750;
  assign tmp29508 = s0 ? tmp27750 : tmp29488;
  assign tmp29506 = s1 ? tmp29507 : tmp29508;
  assign tmp29510 = s0 ? tmp27750 : tmp29485;
  assign tmp29511 = s0 ? tmp29193 : tmp27750;
  assign tmp29509 = s1 ? tmp29510 : tmp29511;
  assign tmp29505 = s2 ? tmp29506 : tmp29509;
  assign tmp29514 = s0 ? tmp27750 : tmp29207;
  assign tmp29513 = s1 ? tmp29508 : tmp29514;
  assign tmp29515 = s1 ? tmp29191 : tmp29351;
  assign tmp29512 = s2 ? tmp29513 : tmp29515;
  assign tmp29504 = s3 ? tmp29505 : tmp29512;
  assign tmp29519 = s0 ? tmp27750 : tmp29352;
  assign tmp29520 = s0 ? tmp27784 : tmp27743;
  assign tmp29518 = s1 ? tmp29519 : tmp29520;
  assign tmp29521 = s1 ? tmp29520 : tmp29494;
  assign tmp29517 = s2 ? tmp29518 : tmp29521;
  assign tmp29524 = s0 ? tmp29230 : tmp29205;
  assign tmp29523 = s1 ? tmp29524 : tmp29206;
  assign tmp29522 = ~(s2 ? tmp29523 : tmp27791);
  assign tmp29516 = s3 ? tmp29517 : tmp29522;
  assign tmp29503 = s4 ? tmp29504 : tmp29516;
  assign tmp29529 = s0 ? tmp29207 : tmp27750;
  assign tmp29528 = s1 ? tmp29529 : tmp29213;
  assign tmp29531 = s0 ? tmp29217 : tmp29230;
  assign tmp29532 = s0 ? 1 : tmp29230;
  assign tmp29530 = ~(s1 ? tmp29531 : tmp29532);
  assign tmp29527 = s2 ? tmp29528 : tmp29530;
  assign tmp29526 = s3 ? tmp29527 : tmp29220;
  assign tmp29537 = ~(l1 ? tmp28835 : tmp27809);
  assign tmp29536 = s0 ? tmp27750 : tmp29537;
  assign tmp29538 = ~(s0 ? tmp29230 : 1);
  assign tmp29535 = ~(s1 ? tmp29536 : tmp29538);
  assign tmp29534 = s2 ? tmp29228 : tmp29535;
  assign tmp29533 = ~(s3 ? tmp29534 : tmp29237);
  assign tmp29525 = s4 ? tmp29526 : tmp29533;
  assign tmp29502 = s5 ? tmp29503 : tmp29525;
  assign tmp29480 = s6 ? tmp29481 : tmp29502;
  assign tmp29479 = s7 ? tmp29480 : tmp27575;
  assign tmp29478 = s8 ? tmp29399 : tmp29479;
  assign tmp29320 = s9 ? tmp29321 : tmp29478;
  assign tmp29546 = s0 ? tmp27991 : tmp29485;
  assign tmp29545 = s1 ? tmp29327 : tmp29546;
  assign tmp29549 = l1 ? tmp27980 : tmp27560;
  assign tmp29548 = s0 ? tmp29549 : tmp29352;
  assign tmp29551 = s0 ? tmp29549 : 1;
  assign tmp29550 = s1 ? tmp29551 : tmp29352;
  assign tmp29547 = s2 ? tmp29548 : tmp29550;
  assign tmp29544 = s3 ? tmp29545 : tmp29547;
  assign tmp29555 = s0 ? tmp29488 : tmp27991;
  assign tmp29554 = s1 ? tmp29555 : tmp29352;
  assign tmp29557 = s0 ? tmp27991 : 1;
  assign tmp29556 = s1 ? tmp29346 : tmp29557;
  assign tmp29553 = s2 ? tmp29554 : tmp29556;
  assign tmp29559 = s1 ? tmp27991 : 1;
  assign tmp29561 = s0 ? tmp29268 : tmp29352;
  assign tmp29560 = s1 ? tmp29351 : tmp29561;
  assign tmp29558 = s2 ? tmp29559 : tmp29560;
  assign tmp29552 = s3 ? tmp29553 : tmp29558;
  assign tmp29543 = s4 ? tmp29544 : tmp29552;
  assign tmp29567 = s0 ? tmp29485 : 1;
  assign tmp29568 = s0 ? 1 : tmp29549;
  assign tmp29566 = s1 ? tmp29567 : tmp29568;
  assign tmp29571 = l1 ? tmp28741 : tmp27499;
  assign tmp29570 = s0 ? 1 : tmp29571;
  assign tmp29569 = s1 ? tmp29570 : tmp29364;
  assign tmp29565 = s2 ? tmp29566 : tmp29569;
  assign tmp29574 = s0 ? 1 : tmp29137;
  assign tmp29573 = s1 ? tmp29568 : tmp29574;
  assign tmp29576 = s0 ? tmp29372 : tmp29031;
  assign tmp29575 = s1 ? tmp29286 : tmp29576;
  assign tmp29572 = s2 ? tmp29573 : tmp29575;
  assign tmp29564 = s3 ? tmp29565 : tmp29572;
  assign tmp29580 = s0 ? tmp27991 : tmp27836;
  assign tmp29579 = s1 ? tmp29376 : tmp29580;
  assign tmp29583 = l1 ? tmp27980 : tmp27499;
  assign tmp29582 = s0 ? tmp29583 : tmp27991;
  assign tmp29581 = s1 ? tmp29580 : tmp29582;
  assign tmp29578 = s2 ? tmp29579 : tmp29581;
  assign tmp29587 = l1 ? 1 : tmp27606;
  assign tmp29586 = s0 ? tmp29587 : tmp29001;
  assign tmp29585 = s1 ? tmp29586 : tmp29299;
  assign tmp29584 = ~(s2 ? tmp29585 : 0);
  assign tmp29577 = s3 ? tmp29578 : tmp29584;
  assign tmp29563 = s4 ? tmp29564 : tmp29577;
  assign tmp29592 = s0 ? tmp29137 : 1;
  assign tmp29591 = s1 ? tmp29592 : tmp29139;
  assign tmp29594 = s0 ? tmp27697 : tmp28267;
  assign tmp29593 = ~(s1 ? tmp29594 : tmp28818);
  assign tmp29590 = s2 ? tmp29591 : tmp29593;
  assign tmp29589 = s3 ? tmp29590 : tmp29119;
  assign tmp29599 = ~(l1 ? tmp28835 : tmp27606);
  assign tmp29598 = s0 ? 1 : tmp29599;
  assign tmp29600 = ~(s0 ? tmp28267 : 1);
  assign tmp29597 = ~(s1 ? tmp29598 : tmp29600);
  assign tmp29596 = s2 ? tmp29310 : tmp29597;
  assign tmp29595 = ~(s3 ? tmp29596 : tmp29317);
  assign tmp29588 = s4 ? tmp29589 : tmp29595;
  assign tmp29562 = s5 ? tmp29563 : tmp29588;
  assign tmp29542 = s6 ? tmp29543 : tmp29562;
  assign tmp29541 = s7 ? tmp29542 : tmp27575;
  assign tmp29540 = s8 ? tmp29541 : tmp29542;
  assign tmp29539 = s9 ? tmp29540 : tmp27575;
  assign tmp29319 = s10 ? tmp29320 : tmp29539;
  assign tmp28921 = s12 ? tmp28922 : tmp29319;
  assign tmp28426 = s13 ? tmp28427 : tmp28921;
  assign tmp27475 = s14 ? tmp27476 : tmp28426;
  assign tmp29612 = l1 ? tmp29088 : 0;
  assign tmp29615 = l2 ? 1 : tmp27615;
  assign tmp29614 = l1 ? tmp29615 : 1;
  assign tmp29613 = ~(s0 ? 1 : tmp29614);
  assign tmp29611 = s1 ? tmp29612 : tmp29613;
  assign tmp29620 = l2 ? tmp27490 : tmp27487;
  assign tmp29621 = ~(l2 ? tmp27615 : 1);
  assign tmp29619 = ~(l1 ? tmp29620 : tmp29621);
  assign tmp29618 = s0 ? 1 : tmp29619;
  assign tmp29623 = l1 ? tmp28835 : 1;
  assign tmp29622 = s0 ? tmp29623 : tmp29619;
  assign tmp29617 = s1 ? tmp29618 : tmp29622;
  assign tmp29625 = s0 ? tmp29623 : 1;
  assign tmp29624 = s1 ? tmp29625 : tmp29619;
  assign tmp29616 = ~(s2 ? tmp29617 : tmp29624);
  assign tmp29610 = s3 ? tmp29611 : tmp29616;
  assign tmp29628 = s1 ? 1 : tmp29619;
  assign tmp29630 = s0 ? tmp29612 : 0;
  assign tmp29629 = ~(s1 ? tmp29630 : 0);
  assign tmp29627 = s2 ? tmp29628 : tmp29629;
  assign tmp29634 = ~(l1 ? tmp29414 : tmp27497);
  assign tmp29633 = s0 ? 1 : tmp29634;
  assign tmp29632 = s1 ? 1 : tmp29633;
  assign tmp29637 = l1 ? tmp29620 : tmp29621;
  assign tmp29638 = l1 ? tmp27490 : tmp29621;
  assign tmp29636 = s0 ? tmp29637 : tmp29638;
  assign tmp29640 = l1 ? tmp27490 : tmp27497;
  assign tmp29639 = s0 ? tmp29640 : tmp29637;
  assign tmp29635 = ~(s1 ? tmp29636 : tmp29639);
  assign tmp29631 = s2 ? tmp29632 : tmp29635;
  assign tmp29626 = ~(s3 ? tmp29627 : tmp29631);
  assign tmp29609 = s4 ? tmp29610 : tmp29626;
  assign tmp29646 = s0 ? tmp29614 : 1;
  assign tmp29645 = s1 ? tmp29646 : 1;
  assign tmp29648 = s0 ? 1 : tmp29614;
  assign tmp29649 = ~(s0 ? tmp29638 : 0);
  assign tmp29647 = s1 ? tmp29648 : tmp29649;
  assign tmp29644 = s2 ? tmp29645 : tmp29647;
  assign tmp29652 = s0 ? 1 : tmp28248;
  assign tmp29654 = ~(l1 ? tmp27490 : tmp29621);
  assign tmp29653 = s0 ? 1 : tmp29654;
  assign tmp29651 = s1 ? tmp29652 : tmp29653;
  assign tmp29657 = l1 ? tmp29414 : tmp27517;
  assign tmp29656 = s0 ? tmp29640 : tmp29657;
  assign tmp29658 = s0 ? tmp29637 : tmp29640;
  assign tmp29655 = ~(s1 ? tmp29656 : tmp29658);
  assign tmp29650 = s2 ? tmp29651 : tmp29655;
  assign tmp29643 = s3 ? tmp29644 : tmp29650;
  assign tmp29663 = l1 ? tmp29620 : 0;
  assign tmp29662 = s0 ? tmp27494 : tmp29663;
  assign tmp29661 = s1 ? tmp29662 : 0;
  assign tmp29660 = s2 ? tmp29661 : 0;
  assign tmp29666 = s0 ? 1 : tmp28249;
  assign tmp29668 = ~(l1 ? tmp27490 : tmp27497);
  assign tmp29667 = s0 ? 1 : tmp29668;
  assign tmp29665 = s1 ? tmp29666 : tmp29667;
  assign tmp29671 = l1 ? tmp29414 : tmp27497;
  assign tmp29670 = s0 ? tmp29671 : tmp27548;
  assign tmp29669 = ~(s1 ? tmp27548 : tmp29670);
  assign tmp29664 = ~(s2 ? tmp29665 : tmp29669);
  assign tmp29659 = ~(s3 ? tmp29660 : tmp29664);
  assign tmp29642 = s4 ? tmp29643 : tmp29659;
  assign tmp29676 = s0 ? tmp29638 : tmp27495;
  assign tmp29677 = s0 ? tmp27495 : tmp27833;
  assign tmp29675 = s1 ? tmp29676 : tmp29677;
  assign tmp29678 = ~(s1 ? tmp28236 : 1);
  assign tmp29674 = s2 ? tmp29675 : tmp29678;
  assign tmp29682 = ~(l1 ? tmp27490 : tmp27517);
  assign tmp29681 = s0 ? 1 : tmp29682;
  assign tmp29680 = s1 ? 1 : tmp29681;
  assign tmp29685 = l1 ? tmp27490 : tmp27517;
  assign tmp29684 = s0 ? tmp29685 : tmp27533;
  assign tmp29683 = ~(s1 ? tmp29684 : tmp27537);
  assign tmp29679 = ~(s2 ? tmp29680 : tmp29683);
  assign tmp29673 = s3 ? tmp29674 : tmp29679;
  assign tmp29689 = ~(s0 ? tmp28214 : tmp29640);
  assign tmp29688 = s1 ? tmp29666 : tmp29689;
  assign tmp29692 = ~(l1 ? tmp27897 : 1);
  assign tmp29691 = s0 ? tmp27495 : tmp29692;
  assign tmp29690 = ~(s1 ? tmp29691 : 0);
  assign tmp29687 = s2 ? tmp29688 : tmp29690;
  assign tmp29695 = s0 ? tmp27504 : tmp29682;
  assign tmp29696 = ~(s0 ? tmp29685 : tmp28214);
  assign tmp29694 = s1 ? tmp29695 : tmp29696;
  assign tmp29698 = ~(s0 ? 1 : tmp28249);
  assign tmp29697 = ~(s1 ? tmp27537 : tmp29698);
  assign tmp29693 = s2 ? tmp29694 : tmp29697;
  assign tmp29686 = ~(s3 ? tmp29687 : tmp29693);
  assign tmp29672 = ~(s4 ? tmp29673 : tmp29686);
  assign tmp29641 = ~(s5 ? tmp29642 : tmp29672);
  assign tmp29608 = s6 ? tmp29609 : tmp29641;
  assign tmp29607 = s7 ? tmp29608 : tmp27495;
  assign tmp29706 = ~(l1 ? tmp27560 : tmp27497);
  assign tmp29705 = s0 ? 1 : tmp29706;
  assign tmp29704 = s1 ? 1 : tmp29705;
  assign tmp29703 = s2 ? tmp29704 : tmp29635;
  assign tmp29702 = ~(s3 ? tmp29627 : tmp29703);
  assign tmp29701 = s4 ? tmp29610 : tmp29702;
  assign tmp29713 = l1 ? tmp27560 : tmp27504;
  assign tmp29712 = s0 ? tmp29640 : tmp29713;
  assign tmp29711 = ~(s1 ? tmp29712 : tmp29658);
  assign tmp29710 = s2 ? tmp29651 : tmp29711;
  assign tmp29709 = s3 ? tmp29644 : tmp29710;
  assign tmp29717 = s0 ? tmp27617 : tmp29663;
  assign tmp29716 = s1 ? tmp29717 : 0;
  assign tmp29715 = s2 ? tmp29716 : 0;
  assign tmp29721 = l1 ? tmp27560 : tmp27497;
  assign tmp29720 = s0 ? tmp29721 : tmp27636;
  assign tmp29719 = ~(s1 ? tmp27636 : tmp29720);
  assign tmp29718 = ~(s2 ? tmp29665 : tmp29719);
  assign tmp29714 = ~(s3 ? tmp29715 : tmp29718);
  assign tmp29708 = s4 ? tmp29709 : tmp29714;
  assign tmp29726 = s0 ? tmp29638 : 1;
  assign tmp29728 = ~(l1 ? tmp27504 : 1);
  assign tmp29727 = s0 ? 1 : tmp29728;
  assign tmp29725 = s1 ? tmp29726 : tmp29727;
  assign tmp29729 = ~(s1 ? tmp27842 : 1);
  assign tmp29724 = s2 ? tmp29725 : tmp29729;
  assign tmp29733 = ~(l1 ? tmp27490 : tmp27504);
  assign tmp29732 = s0 ? 1 : tmp29733;
  assign tmp29731 = s1 ? 1 : tmp29732;
  assign tmp29736 = l1 ? tmp27490 : tmp27504;
  assign tmp29735 = s0 ? tmp29736 : tmp27640;
  assign tmp29734 = ~(s1 ? tmp29735 : tmp27646);
  assign tmp29730 = ~(s2 ? tmp29731 : tmp29734);
  assign tmp29723 = s3 ? tmp29724 : tmp29730;
  assign tmp29740 = s0 ? 1 : tmp29692;
  assign tmp29739 = ~(s1 ? tmp29740 : 0);
  assign tmp29738 = s2 ? tmp29688 : tmp29739;
  assign tmp29743 = s0 ? tmp27836 : tmp29733;
  assign tmp29744 = ~(s0 ? tmp29736 : tmp28214);
  assign tmp29742 = s1 ? tmp29743 : tmp29744;
  assign tmp29745 = ~(s1 ? tmp27646 : tmp29698);
  assign tmp29741 = s2 ? tmp29742 : tmp29745;
  assign tmp29737 = ~(s3 ? tmp29738 : tmp29741);
  assign tmp29722 = ~(s4 ? tmp29723 : tmp29737);
  assign tmp29707 = ~(s5 ? tmp29708 : tmp29722);
  assign tmp29700 = s6 ? tmp29701 : tmp29707;
  assign tmp29699 = s7 ? tmp29700 : tmp27495;
  assign tmp29606 = s8 ? tmp29607 : tmp29699;
  assign tmp29752 = l1 ? tmp29088 : tmp27809;
  assign tmp29754 = l1 ? tmp29615 : tmp27744;
  assign tmp29753 = ~(s0 ? tmp27750 : tmp29754);
  assign tmp29751 = s1 ? tmp29752 : tmp29753;
  assign tmp29759 = ~(l2 ? tmp27615 : tmp27496);
  assign tmp29758 = ~(l1 ? tmp29620 : tmp29759);
  assign tmp29757 = s0 ? tmp27750 : tmp29758;
  assign tmp29761 = l1 ? tmp28835 : tmp27744;
  assign tmp29760 = s0 ? tmp29761 : tmp29758;
  assign tmp29756 = s1 ? tmp29757 : tmp29760;
  assign tmp29763 = s0 ? tmp29761 : tmp27750;
  assign tmp29762 = s1 ? tmp29763 : tmp29758;
  assign tmp29755 = ~(s2 ? tmp29756 : tmp29762);
  assign tmp29750 = s3 ? tmp29751 : tmp29755;
  assign tmp29766 = s1 ? tmp27750 : tmp29758;
  assign tmp29768 = s0 ? tmp29752 : tmp27791;
  assign tmp29767 = ~(s1 ? tmp29768 : tmp27791);
  assign tmp29765 = s2 ? tmp29766 : tmp29767;
  assign tmp29772 = ~(l1 ? tmp27560 : tmp27521);
  assign tmp29771 = s0 ? tmp27750 : tmp29772;
  assign tmp29770 = s1 ? tmp27750 : tmp29771;
  assign tmp29775 = l1 ? tmp29620 : tmp29759;
  assign tmp29776 = l1 ? tmp27490 : tmp29759;
  assign tmp29774 = s0 ? tmp29775 : tmp29776;
  assign tmp29778 = l1 ? tmp27490 : tmp27521;
  assign tmp29777 = s0 ? tmp29778 : tmp29775;
  assign tmp29773 = ~(s1 ? tmp29774 : tmp29777);
  assign tmp29769 = s2 ? tmp29770 : tmp29773;
  assign tmp29764 = ~(s3 ? tmp29765 : tmp29769);
  assign tmp29749 = s4 ? tmp29750 : tmp29764;
  assign tmp29784 = s0 ? tmp29754 : tmp27750;
  assign tmp29783 = s1 ? tmp29784 : tmp27750;
  assign tmp29786 = s0 ? tmp27750 : tmp29754;
  assign tmp29787 = ~(s0 ? tmp29776 : tmp27791);
  assign tmp29785 = s1 ? tmp29786 : tmp29787;
  assign tmp29782 = s2 ? tmp29783 : tmp29785;
  assign tmp29790 = s0 ? tmp27750 : tmp28378;
  assign tmp29792 = ~(l1 ? tmp27490 : tmp29759);
  assign tmp29791 = s0 ? tmp27750 : tmp29792;
  assign tmp29789 = s1 ? tmp29790 : tmp29791;
  assign tmp29795 = l1 ? tmp27560 : tmp27760;
  assign tmp29794 = s0 ? tmp29778 : tmp29795;
  assign tmp29796 = s0 ? tmp29775 : tmp29778;
  assign tmp29793 = ~(s1 ? tmp29794 : tmp29796);
  assign tmp29788 = s2 ? tmp29789 : tmp29793;
  assign tmp29781 = s3 ? tmp29782 : tmp29788;
  assign tmp29801 = l1 ? tmp29620 : tmp27809;
  assign tmp29800 = s0 ? tmp29204 : tmp29801;
  assign tmp29799 = s1 ? tmp29800 : tmp27791;
  assign tmp29798 = s2 ? tmp29799 : tmp27791;
  assign tmp29804 = s0 ? tmp27750 : tmp28379;
  assign tmp29806 = ~(l1 ? tmp27490 : tmp27521);
  assign tmp29805 = s0 ? tmp27750 : tmp29806;
  assign tmp29803 = s1 ? tmp29804 : tmp29805;
  assign tmp29809 = l1 ? tmp27560 : tmp27521;
  assign tmp29808 = s0 ? tmp29809 : tmp27762;
  assign tmp29807 = ~(s1 ? tmp27762 : tmp29808);
  assign tmp29802 = ~(s2 ? tmp29803 : tmp29807);
  assign tmp29797 = ~(s3 ? tmp29798 : tmp29802);
  assign tmp29780 = s4 ? tmp29781 : tmp29797;
  assign tmp29814 = s0 ? tmp29776 : 1;
  assign tmp29816 = ~(l1 ? tmp27504 : tmp27744);
  assign tmp29815 = s0 ? 1 : tmp29816;
  assign tmp29813 = s1 ? tmp29814 : tmp29815;
  assign tmp29817 = ~(s1 ? tmp27749 : tmp27750);
  assign tmp29812 = s2 ? tmp29813 : tmp29817;
  assign tmp29821 = ~(l1 ? tmp27490 : tmp27760);
  assign tmp29820 = s0 ? tmp27750 : tmp29821;
  assign tmp29819 = s1 ? tmp27750 : tmp29820;
  assign tmp29824 = l1 ? tmp27490 : tmp27760;
  assign tmp29823 = s0 ? tmp29824 : tmp29230;
  assign tmp29825 = s0 ? tmp29230 : tmp27791;
  assign tmp29822 = ~(s1 ? tmp29823 : tmp29825);
  assign tmp29818 = ~(s2 ? tmp29819 : tmp29822);
  assign tmp29811 = s3 ? tmp29812 : tmp29818;
  assign tmp29829 = ~(s0 ? tmp28342 : tmp29778);
  assign tmp29828 = s1 ? tmp29804 : tmp29829;
  assign tmp29832 = ~(l1 ? tmp27897 : tmp27744);
  assign tmp29831 = s0 ? 1 : tmp29832;
  assign tmp29830 = ~(s1 ? tmp29831 : tmp27791);
  assign tmp29827 = s2 ? tmp29828 : tmp29830;
  assign tmp29835 = s0 ? tmp27743 : tmp29821;
  assign tmp29836 = ~(s0 ? tmp29824 : tmp28342);
  assign tmp29834 = s1 ? tmp29835 : tmp29836;
  assign tmp29838 = ~(s0 ? tmp27750 : tmp28379);
  assign tmp29837 = ~(s1 ? tmp29825 : tmp29838);
  assign tmp29833 = s2 ? tmp29834 : tmp29837;
  assign tmp29826 = ~(s3 ? tmp29827 : tmp29833);
  assign tmp29810 = ~(s4 ? tmp29811 : tmp29826);
  assign tmp29779 = ~(s5 ? tmp29780 : tmp29810);
  assign tmp29748 = s6 ? tmp29749 : tmp29779;
  assign tmp29747 = s7 ? tmp29748 : tmp27495;
  assign tmp29746 = s8 ? tmp29699 : tmp29747;
  assign tmp29605 = s9 ? tmp29606 : tmp29746;
  assign tmp29840 = s8 ? tmp29699 : tmp29700;
  assign tmp29839 = s9 ? tmp29840 : tmp27495;
  assign tmp29604 = s10 ? tmp29605 : tmp29839;
  assign tmp29850 = ~(l2 ? 1 : tmp27615);
  assign tmp29849 = l1 ? tmp27497 : tmp29850;
  assign tmp29848 = s1 ? tmp29849 : 0;
  assign tmp29853 = ~(l1 ? tmp27497 : tmp27487);
  assign tmp29852 = s0 ? 1 : tmp29853;
  assign tmp29854 = s1 ? 1 : tmp29853;
  assign tmp29851 = ~(s2 ? tmp29852 : tmp29854);
  assign tmp29847 = s3 ? tmp29848 : tmp29851;
  assign tmp29858 = s0 ? tmp29849 : 0;
  assign tmp29857 = ~(s1 ? tmp29858 : 0);
  assign tmp29856 = s2 ? tmp29854 : tmp29857;
  assign tmp29862 = ~(l1 ? tmp27517 : tmp27490);
  assign tmp29861 = s0 ? 1 : tmp29862;
  assign tmp29860 = s1 ? 1 : tmp29861;
  assign tmp29864 = l1 ? tmp27497 : tmp27487;
  assign tmp29866 = l1 ? tmp27497 : tmp27490;
  assign tmp29865 = s0 ? tmp29866 : tmp29864;
  assign tmp29863 = ~(s1 ? tmp29864 : tmp29865);
  assign tmp29859 = s2 ? tmp29860 : tmp29863;
  assign tmp29855 = ~(s3 ? tmp29856 : tmp29859);
  assign tmp29846 = s4 ? tmp29847 : tmp29855;
  assign tmp29872 = ~(s0 ? tmp29864 : 0);
  assign tmp29871 = s1 ? 1 : tmp29872;
  assign tmp29870 = s2 ? 1 : tmp29871;
  assign tmp29877 = ~(l2 ? tmp27615 : tmp27506);
  assign tmp29876 = ~(l1 ? tmp27497 : tmp29877);
  assign tmp29875 = s0 ? 1 : tmp29876;
  assign tmp29874 = s1 ? 1 : tmp29875;
  assign tmp29880 = l1 ? tmp27517 : tmp27495;
  assign tmp29879 = s0 ? tmp29866 : tmp29880;
  assign tmp29882 = l1 ? tmp27497 : tmp29877;
  assign tmp29881 = s0 ? tmp29882 : tmp29866;
  assign tmp29878 = ~(s1 ? tmp29879 : tmp29881);
  assign tmp29873 = s2 ? tmp29874 : tmp29878;
  assign tmp29869 = s3 ? tmp29870 : tmp29873;
  assign tmp29887 = l1 ? tmp27517 : tmp27490;
  assign tmp29888 = l1 ? tmp27497 : tmp28226;
  assign tmp29886 = s0 ? tmp29887 : tmp29888;
  assign tmp29885 = s1 ? tmp29886 : 0;
  assign tmp29884 = s2 ? tmp29885 : 0;
  assign tmp29892 = ~(l1 ? tmp27497 : tmp28226);
  assign tmp29891 = s0 ? 1 : tmp29892;
  assign tmp29894 = ~(l1 ? tmp27497 : tmp27490);
  assign tmp29893 = s0 ? 1 : tmp29894;
  assign tmp29890 = s1 ? tmp29891 : tmp29893;
  assign tmp29896 = s0 ? tmp29887 : tmp27495;
  assign tmp29895 = ~(s1 ? tmp27495 : tmp29896);
  assign tmp29889 = ~(s2 ? tmp29890 : tmp29895);
  assign tmp29883 = ~(s3 ? tmp29884 : tmp29889);
  assign tmp29868 = s4 ? tmp29869 : tmp29883;
  assign tmp29901 = s0 ? tmp29882 : tmp29880;
  assign tmp29902 = s0 ? tmp29880 : 0;
  assign tmp29900 = s1 ? tmp29901 : tmp29902;
  assign tmp29899 = s2 ? tmp29900 : 0;
  assign tmp29905 = s0 ? 1 : tmp27506;
  assign tmp29907 = ~(l1 ? 1 : tmp27575);
  assign tmp29906 = ~(s0 ? tmp27490 : tmp29907);
  assign tmp29904 = s1 ? tmp29905 : tmp29906;
  assign tmp29909 = s0 ? tmp28446 : tmp29862;
  assign tmp29910 = ~(s0 ? tmp29887 : 0);
  assign tmp29908 = s1 ? tmp29909 : tmp29910;
  assign tmp29903 = ~(s2 ? tmp29904 : tmp29908);
  assign tmp29898 = s3 ? tmp29899 : tmp29903;
  assign tmp29913 = s1 ? 1 : tmp29893;
  assign tmp29914 = ~(s1 ? tmp29902 : 0);
  assign tmp29912 = s2 ? tmp29913 : tmp29914;
  assign tmp29917 = s0 ? 1 : tmp28442;
  assign tmp29918 = s0 ? tmp28446 : tmp29892;
  assign tmp29916 = s1 ? tmp29917 : tmp29918;
  assign tmp29920 = s0 ? tmp29887 : 0;
  assign tmp29921 = s0 ? tmp27490 : 0;
  assign tmp29919 = ~(s1 ? tmp29920 : tmp29921);
  assign tmp29915 = s2 ? tmp29916 : tmp29919;
  assign tmp29911 = ~(s3 ? tmp29912 : tmp29915);
  assign tmp29897 = ~(s4 ? tmp29898 : tmp29911);
  assign tmp29867 = ~(s5 ? tmp29868 : tmp29897);
  assign tmp29845 = s6 ? tmp29846 : tmp29867;
  assign tmp29844 = s7 ? tmp29845 : tmp27495;
  assign tmp29926 = s1 ? tmp29864 : 0;
  assign tmp29925 = s3 ? tmp29926 : tmp29851;
  assign tmp29930 = s0 ? tmp29864 : 0;
  assign tmp29929 = ~(s1 ? tmp29930 : 0);
  assign tmp29928 = s2 ? tmp29854 : tmp29929;
  assign tmp29934 = ~(l1 ? tmp27504 : tmp27490);
  assign tmp29933 = s0 ? 1 : tmp29934;
  assign tmp29932 = s1 ? 1 : tmp29933;
  assign tmp29931 = s2 ? tmp29932 : tmp29863;
  assign tmp29927 = ~(s3 ? tmp29928 : tmp29931);
  assign tmp29924 = s4 ? tmp29925 : tmp29927;
  assign tmp29940 = s0 ? tmp29866 : tmp27836;
  assign tmp29939 = ~(s1 ? tmp29940 : tmp29881);
  assign tmp29938 = s2 ? tmp29874 : tmp29939;
  assign tmp29937 = s3 ? tmp29870 : tmp29938;
  assign tmp29945 = l1 ? tmp27504 : tmp27490;
  assign tmp29944 = s0 ? tmp29945 : tmp29888;
  assign tmp29943 = s1 ? tmp29944 : 0;
  assign tmp29942 = s2 ? tmp29943 : 0;
  assign tmp29948 = s0 ? tmp29945 : 1;
  assign tmp29947 = ~(s1 ? 1 : tmp29948);
  assign tmp29946 = ~(s2 ? tmp29893 : tmp29947);
  assign tmp29941 = ~(s3 ? tmp29942 : tmp29946);
  assign tmp29936 = s4 ? tmp29937 : tmp29941;
  assign tmp29953 = s0 ? tmp29882 : tmp27836;
  assign tmp29954 = s0 ? tmp27836 : 0;
  assign tmp29952 = s1 ? tmp29953 : tmp29954;
  assign tmp29951 = s2 ? tmp29952 : 0;
  assign tmp29958 = ~(l1 ? 1 : 0);
  assign tmp29957 = ~(s0 ? tmp27490 : tmp29958);
  assign tmp29956 = s1 ? tmp29905 : tmp29957;
  assign tmp29960 = s0 ? tmp27640 : tmp29934;
  assign tmp29961 = ~(s0 ? tmp29945 : 0);
  assign tmp29959 = s1 ? tmp29960 : tmp29961;
  assign tmp29955 = ~(s2 ? tmp29956 : tmp29959);
  assign tmp29950 = s3 ? tmp29951 : tmp29955;
  assign tmp29964 = ~(s1 ? tmp29954 : 0);
  assign tmp29963 = s2 ? tmp29913 : tmp29964;
  assign tmp29967 = s0 ? 1 : tmp28494;
  assign tmp29968 = s0 ? tmp27640 : tmp29892;
  assign tmp29966 = s1 ? tmp29967 : tmp29968;
  assign tmp29970 = s0 ? tmp29945 : 0;
  assign tmp29969 = ~(s1 ? tmp29970 : tmp29921);
  assign tmp29965 = s2 ? tmp29966 : tmp29969;
  assign tmp29962 = ~(s3 ? tmp29963 : tmp29965);
  assign tmp29949 = ~(s4 ? tmp29950 : tmp29962);
  assign tmp29935 = ~(s5 ? tmp29936 : tmp29949);
  assign tmp29923 = s6 ? tmp29924 : tmp29935;
  assign tmp29922 = s7 ? tmp29923 : tmp27495;
  assign tmp29843 = s8 ? tmp29844 : tmp29922;
  assign tmp29979 = l3 ? tmp27488 : tmp27492;
  assign tmp29978 = ~(l2 ? 1 : tmp29979);
  assign tmp29977 = l1 ? tmp27497 : tmp29978;
  assign tmp29976 = s1 ? tmp29977 : tmp27791;
  assign tmp29983 = ~(l2 ? tmp27615 : tmp29979);
  assign tmp29982 = ~(l1 ? tmp27497 : tmp29983);
  assign tmp29981 = s0 ? tmp27750 : tmp29982;
  assign tmp29984 = s1 ? tmp27750 : tmp29982;
  assign tmp29980 = ~(s2 ? tmp29981 : tmp29984);
  assign tmp29975 = s3 ? tmp29976 : tmp29980;
  assign tmp29988 = s0 ? tmp29977 : tmp27791;
  assign tmp29987 = ~(s1 ? tmp29988 : tmp27791);
  assign tmp29986 = s2 ? tmp29984 : tmp29987;
  assign tmp29992 = ~(l1 ? tmp27504 : tmp28080);
  assign tmp29991 = s0 ? tmp27750 : tmp29992;
  assign tmp29990 = s1 ? tmp27750 : tmp29991;
  assign tmp29994 = l1 ? tmp27497 : tmp29983;
  assign tmp29996 = l1 ? tmp27497 : tmp28080;
  assign tmp29995 = s0 ? tmp29996 : tmp29994;
  assign tmp29993 = ~(s1 ? tmp29994 : tmp29995);
  assign tmp29989 = s2 ? tmp29990 : tmp29993;
  assign tmp29985 = ~(s3 ? tmp29986 : tmp29989);
  assign tmp29974 = s4 ? tmp29975 : tmp29985;
  assign tmp30002 = ~(s0 ? tmp29994 : tmp27791);
  assign tmp30001 = s1 ? tmp27750 : tmp30002;
  assign tmp30000 = s2 ? tmp27750 : tmp30001;
  assign tmp30007 = ~(l2 ? tmp27615 : tmp28324);
  assign tmp30006 = ~(l1 ? tmp27497 : tmp30007);
  assign tmp30005 = s0 ? tmp27750 : tmp30006;
  assign tmp30004 = s1 ? tmp27750 : tmp30005;
  assign tmp30009 = s0 ? tmp29996 : tmp27836;
  assign tmp30011 = l1 ? tmp27497 : tmp30007;
  assign tmp30010 = s0 ? tmp30011 : tmp29996;
  assign tmp30008 = ~(s1 ? tmp30009 : tmp30010);
  assign tmp30003 = s2 ? tmp30004 : tmp30008;
  assign tmp29999 = s3 ? tmp30000 : tmp30003;
  assign tmp30016 = l1 ? tmp27504 : tmp28080;
  assign tmp30018 = ~(l2 ? 1 : tmp28324);
  assign tmp30017 = l1 ? tmp27497 : tmp30018;
  assign tmp30015 = s0 ? tmp30016 : tmp30017;
  assign tmp30014 = s1 ? tmp30015 : tmp27791;
  assign tmp30013 = s2 ? tmp30014 : tmp27791;
  assign tmp30022 = ~(l1 ? tmp27497 : tmp30018);
  assign tmp30021 = s0 ? tmp27750 : tmp30022;
  assign tmp30024 = ~(l1 ? tmp27497 : tmp28080);
  assign tmp30023 = s0 ? tmp27750 : tmp30024;
  assign tmp30020 = s1 ? tmp30021 : tmp30023;
  assign tmp30026 = s0 ? tmp30016 : 1;
  assign tmp30025 = ~(s1 ? 1 : tmp30026);
  assign tmp30019 = ~(s2 ? tmp30020 : tmp30025);
  assign tmp30012 = ~(s3 ? tmp30013 : tmp30019);
  assign tmp29998 = s4 ? tmp29999 : tmp30012;
  assign tmp30031 = s0 ? tmp30011 : tmp27836;
  assign tmp30032 = s0 ? tmp27836 : tmp27791;
  assign tmp30030 = s1 ? tmp30031 : tmp30032;
  assign tmp30029 = s2 ? tmp30030 : tmp27791;
  assign tmp30036 = ~(l1 ? tmp27490 : tmp28080);
  assign tmp30035 = s0 ? tmp27750 : tmp30036;
  assign tmp30037 = ~(s0 ? tmp28079 : tmp29958);
  assign tmp30034 = s1 ? tmp30035 : tmp30037;
  assign tmp30039 = s0 ? tmp27640 : tmp29992;
  assign tmp30040 = ~(s0 ? tmp30016 : tmp27791);
  assign tmp30038 = s1 ? tmp30039 : tmp30040;
  assign tmp30033 = ~(s2 ? tmp30034 : tmp30038);
  assign tmp30028 = s3 ? tmp30029 : tmp30033;
  assign tmp30043 = s1 ? tmp27750 : tmp30023;
  assign tmp30044 = ~(s1 ? tmp30032 : tmp27791);
  assign tmp30042 = s2 ? tmp30043 : tmp30044;
  assign tmp30049 = ~(l2 ? 1 : tmp27554);
  assign tmp30048 = l1 ? 1 : tmp30049;
  assign tmp30047 = s0 ? tmp27750 : tmp30048;
  assign tmp30050 = s0 ? tmp27640 : tmp30024;
  assign tmp30046 = s1 ? tmp30047 : tmp30050;
  assign tmp30052 = s0 ? tmp30016 : tmp27791;
  assign tmp30053 = s0 ? tmp28079 : tmp27791;
  assign tmp30051 = ~(s1 ? tmp30052 : tmp30053);
  assign tmp30045 = s2 ? tmp30046 : tmp30051;
  assign tmp30041 = ~(s3 ? tmp30042 : tmp30045);
  assign tmp30027 = ~(s4 ? tmp30028 : tmp30041);
  assign tmp29997 = ~(s5 ? tmp29998 : tmp30027);
  assign tmp29973 = s6 ? tmp29974 : tmp29997;
  assign tmp29972 = s7 ? tmp29973 : tmp27495;
  assign tmp29971 = s8 ? tmp29922 : tmp29972;
  assign tmp29842 = s9 ? tmp29843 : tmp29971;
  assign tmp30055 = s8 ? tmp29922 : tmp29923;
  assign tmp30054 = s9 ? tmp30055 : tmp27495;
  assign tmp29841 = s10 ? tmp29842 : tmp30054;
  assign tmp29603 = s12 ? tmp29604 : tmp29841;
  assign tmp30065 = l1 ? tmp29088 : tmp28570;
  assign tmp30067 = l1 ? 1 : tmp28643;
  assign tmp30069 = l2 ? tmp27554 : tmp27488;
  assign tmp30068 = l1 ? tmp29615 : tmp30069;
  assign tmp30066 = ~(s0 ? tmp30067 : tmp30068);
  assign tmp30064 = s1 ? tmp30065 : tmp30066;
  assign tmp30072 = l1 ? tmp28835 : tmp28661;
  assign tmp30073 = ~(l1 ? tmp29620 : tmp28570);
  assign tmp30071 = s0 ? tmp30072 : tmp30073;
  assign tmp30075 = s0 ? tmp30072 : 1;
  assign tmp30074 = s1 ? tmp30075 : tmp30073;
  assign tmp30070 = ~(s2 ? tmp30071 : tmp30074);
  assign tmp30063 = s3 ? tmp30064 : tmp30070;
  assign tmp30080 = l1 ? 1 : tmp30069;
  assign tmp30079 = s0 ? tmp30080 : 1;
  assign tmp30078 = s1 ? tmp30079 : tmp30073;
  assign tmp30082 = s0 ? tmp30065 : 0;
  assign tmp30083 = ~(s0 ? tmp30067 : 1);
  assign tmp30081 = ~(s1 ? tmp30082 : tmp30083);
  assign tmp30077 = s2 ? tmp30078 : tmp30081;
  assign tmp30087 = ~(l1 ? tmp29414 : tmp28525);
  assign tmp30086 = s0 ? 1 : tmp30087;
  assign tmp30085 = s1 ? tmp30067 : tmp30086;
  assign tmp30090 = l1 ? tmp29620 : tmp28570;
  assign tmp30091 = l1 ? tmp27490 : tmp28570;
  assign tmp30089 = s0 ? tmp30090 : tmp30091;
  assign tmp30093 = l1 ? tmp27490 : tmp28525;
  assign tmp30092 = s0 ? tmp30093 : tmp30090;
  assign tmp30088 = ~(s1 ? tmp30089 : tmp30092);
  assign tmp30084 = s2 ? tmp30085 : tmp30088;
  assign tmp30076 = ~(s3 ? tmp30077 : tmp30084);
  assign tmp30062 = s4 ? tmp30063 : tmp30076;
  assign tmp30099 = s0 ? tmp30068 : 1;
  assign tmp30098 = s1 ? tmp30099 : 1;
  assign tmp30101 = s0 ? 1 : tmp30068;
  assign tmp30102 = ~(s0 ? tmp30091 : 0);
  assign tmp30100 = s1 ? tmp30101 : tmp30102;
  assign tmp30097 = s2 ? tmp30098 : tmp30100;
  assign tmp30106 = l1 ? tmp27897 : tmp28661;
  assign tmp30105 = s0 ? 1 : tmp30106;
  assign tmp30108 = ~(l1 ? tmp27490 : tmp28608);
  assign tmp30107 = s0 ? 1 : tmp30108;
  assign tmp30104 = s1 ? tmp30105 : tmp30107;
  assign tmp30111 = l1 ? tmp29414 : tmp27833;
  assign tmp30110 = s0 ? tmp30093 : tmp30111;
  assign tmp30113 = l1 ? tmp29620 : tmp28608;
  assign tmp30114 = l1 ? tmp27490 : tmp28608;
  assign tmp30112 = s0 ? tmp30113 : tmp30114;
  assign tmp30109 = ~(s1 ? tmp30110 : tmp30112);
  assign tmp30103 = s2 ? tmp30104 : tmp30109;
  assign tmp30096 = s3 ? tmp30097 : tmp30103;
  assign tmp30119 = l1 ? tmp27495 : tmp28525;
  assign tmp30118 = s0 ? tmp30119 : tmp30113;
  assign tmp30117 = s1 ? tmp30118 : tmp28712;
  assign tmp30121 = s0 ? 1 : tmp28446;
  assign tmp30120 = ~(s1 ? tmp30121 : tmp30079);
  assign tmp30116 = s2 ? tmp30117 : tmp30120;
  assign tmp30125 = ~(l1 ? tmp27490 : tmp27496);
  assign tmp30124 = s0 ? tmp30080 : tmp30125;
  assign tmp30126 = s0 ? tmp28446 : tmp30108;
  assign tmp30123 = s1 ? tmp30124 : tmp30126;
  assign tmp30129 = l1 ? tmp29414 : tmp28525;
  assign tmp30128 = s0 ? tmp30129 : tmp28225;
  assign tmp30127 = ~(s1 ? tmp28225 : tmp30128);
  assign tmp30122 = ~(s2 ? tmp30123 : tmp30127);
  assign tmp30115 = ~(s3 ? tmp30116 : tmp30122);
  assign tmp30095 = s4 ? tmp30096 : tmp30115;
  assign tmp30134 = s0 ? tmp30114 : tmp27533;
  assign tmp30136 = ~(l1 ? tmp27504 : tmp27575);
  assign tmp30135 = s0 ? tmp27533 : tmp30136;
  assign tmp30133 = s1 ? tmp30134 : tmp30135;
  assign tmp30137 = ~(s1 ? tmp27591 : 1);
  assign tmp30132 = s2 ? tmp30133 : tmp30137;
  assign tmp30140 = s0 ? tmp28446 : tmp28210;
  assign tmp30139 = s1 ? tmp30121 : tmp30140;
  assign tmp30142 = s0 ? tmp28196 : tmp27495;
  assign tmp30144 = ~(l1 ? 1 : tmp29464);
  assign tmp30143 = s0 ? tmp27495 : tmp30144;
  assign tmp30141 = ~(s1 ? tmp30142 : tmp30143);
  assign tmp30138 = ~(s2 ? tmp30139 : tmp30141);
  assign tmp30131 = s3 ? tmp30132 : tmp30138;
  assign tmp30148 = s0 ? tmp29463 : tmp27910;
  assign tmp30149 = ~(s0 ? tmp27944 : tmp30093);
  assign tmp30147 = s1 ? tmp30148 : tmp30149;
  assign tmp30152 = ~(l1 ? tmp27897 : tmp30069);
  assign tmp30151 = s0 ? tmp27533 : tmp30152;
  assign tmp30150 = ~(s1 ? tmp30151 : 0);
  assign tmp30146 = s2 ? tmp30147 : tmp30150;
  assign tmp30155 = s0 ? tmp27588 : tmp28210;
  assign tmp30157 = l1 ? tmp27490 : tmp27496;
  assign tmp30156 = ~(s0 ? tmp28196 : tmp30157);
  assign tmp30154 = s1 ? tmp30155 : tmp30156;
  assign tmp30159 = ~(s0 ? tmp28446 : tmp27910);
  assign tmp30158 = ~(s1 ? tmp30143 : tmp30159);
  assign tmp30153 = s2 ? tmp30154 : tmp30158;
  assign tmp30145 = ~(s3 ? tmp30146 : tmp30153);
  assign tmp30130 = ~(s4 ? tmp30131 : tmp30145);
  assign tmp30094 = ~(s5 ? tmp30095 : tmp30130);
  assign tmp30061 = s6 ? tmp30062 : tmp30094;
  assign tmp30060 = s7 ? tmp30061 : tmp27495;
  assign tmp30166 = l1 ? 1 : tmp27623;
  assign tmp30167 = l1 ? tmp29615 : tmp27488;
  assign tmp30165 = ~(s0 ? tmp30166 : tmp30167);
  assign tmp30164 = s1 ? tmp29087 : tmp30165;
  assign tmp30170 = l1 ? tmp28835 : tmp27488;
  assign tmp30169 = s0 ? tmp30170 : tmp30073;
  assign tmp30172 = s0 ? tmp30170 : 1;
  assign tmp30174 = l1 ? tmp29620 : tmp27492;
  assign tmp30173 = ~(s0 ? tmp30090 : tmp30174);
  assign tmp30171 = s1 ? tmp30172 : tmp30173;
  assign tmp30168 = ~(s2 ? tmp30169 : tmp30171);
  assign tmp30163 = s3 ? tmp30164 : tmp30168;
  assign tmp30178 = ~(s0 ? tmp30174 : tmp30090);
  assign tmp30177 = s1 ? tmp28832 : tmp30178;
  assign tmp30180 = s0 ? tmp29087 : 0;
  assign tmp30181 = ~(s0 ? tmp28812 : 1);
  assign tmp30179 = ~(s1 ? tmp30180 : tmp30181);
  assign tmp30176 = s2 ? tmp30177 : tmp30179;
  assign tmp30184 = s0 ? tmp28812 : tmp30166;
  assign tmp30186 = ~(l1 ? tmp27560 : tmp27820);
  assign tmp30185 = s0 ? 1 : tmp30186;
  assign tmp30183 = s1 ? tmp30184 : tmp30185;
  assign tmp30182 = s2 ? tmp30183 : tmp30088;
  assign tmp30175 = ~(s3 ? tmp30176 : tmp30182);
  assign tmp30162 = s4 ? tmp30163 : tmp30175;
  assign tmp30192 = s0 ? tmp30167 : 1;
  assign tmp30191 = s1 ? tmp30192 : 1;
  assign tmp30194 = s0 ? 1 : tmp30167;
  assign tmp30193 = s1 ? tmp30194 : tmp30102;
  assign tmp30190 = s2 ? tmp30191 : tmp30193;
  assign tmp30198 = l1 ? tmp27897 : tmp27488;
  assign tmp30197 = s0 ? 1 : tmp30198;
  assign tmp30196 = s1 ? tmp30197 : tmp30107;
  assign tmp30200 = s0 ? tmp30093 : tmp28258;
  assign tmp30199 = ~(s1 ? tmp30200 : tmp30112);
  assign tmp30195 = s2 ? tmp30196 : tmp30199;
  assign tmp30189 = s3 ? tmp30190 : tmp30195;
  assign tmp30205 = l1 ? tmp29620 : tmp28614;
  assign tmp30204 = s0 ? tmp27858 : tmp30205;
  assign tmp30203 = s1 ? tmp30204 : tmp28811;
  assign tmp30207 = s0 ? 1 : tmp28812;
  assign tmp30206 = ~(s1 ? tmp30207 : tmp28832);
  assign tmp30202 = s2 ? tmp30203 : tmp30206;
  assign tmp30210 = s0 ? tmp28812 : tmp30125;
  assign tmp30212 = ~(l1 ? tmp27490 : tmp27489);
  assign tmp30211 = s0 ? tmp28812 : tmp30212;
  assign tmp30209 = s1 ? tmp30210 : tmp30211;
  assign tmp30214 = s0 ? tmp29249 : tmp28267;
  assign tmp30213 = ~(s1 ? tmp28267 : tmp30214);
  assign tmp30208 = ~(s2 ? tmp30209 : tmp30213);
  assign tmp30201 = ~(s3 ? tmp30202 : tmp30208);
  assign tmp30188 = s4 ? tmp30189 : tmp30201;
  assign tmp30219 = s0 ? tmp30114 : tmp27640;
  assign tmp30220 = s0 ? tmp27640 : tmp29115;
  assign tmp30218 = s1 ? tmp30219 : tmp30220;
  assign tmp30217 = s2 ? tmp30218 : tmp29116;
  assign tmp30223 = s0 ? tmp27640 : tmp28210;
  assign tmp30222 = s1 ? tmp27677 : tmp30223;
  assign tmp30225 = s0 ? tmp28196 : 1;
  assign tmp30227 = ~(l1 ? 1 : tmp27606);
  assign tmp30226 = s0 ? 1 : tmp30227;
  assign tmp30224 = ~(s1 ? tmp30225 : tmp30226);
  assign tmp30221 = ~(s2 ? tmp30222 : tmp30224);
  assign tmp30216 = s3 ? tmp30217 : tmp30221;
  assign tmp30231 = s0 ? tmp29587 : tmp28074;
  assign tmp30232 = ~(s0 ? tmp28115 : tmp30093);
  assign tmp30230 = s1 ? tmp30231 : tmp30232;
  assign tmp30235 = ~(l1 ? tmp27897 : tmp27488);
  assign tmp30234 = s0 ? tmp27640 : tmp30235;
  assign tmp30233 = ~(s1 ? tmp30234 : 0);
  assign tmp30229 = s2 ? tmp30230 : tmp30233;
  assign tmp30238 = s0 ? tmp29118 : tmp28210;
  assign tmp30240 = l1 ? tmp27490 : tmp27744;
  assign tmp30239 = ~(s0 ? tmp28196 : tmp30240);
  assign tmp30237 = s1 ? tmp30238 : tmp30239;
  assign tmp30242 = ~(s0 ? tmp27640 : tmp28074);
  assign tmp30241 = ~(s1 ? tmp30226 : tmp30242);
  assign tmp30236 = s2 ? tmp30237 : tmp30241;
  assign tmp30228 = ~(s3 ? tmp30229 : tmp30236);
  assign tmp30215 = ~(s4 ? tmp30216 : tmp30228);
  assign tmp30187 = ~(s5 ? tmp30188 : tmp30215);
  assign tmp30161 = s6 ? tmp30162 : tmp30187;
  assign tmp30160 = s7 ? tmp30161 : tmp27495;
  assign tmp30059 = s8 ? tmp30060 : tmp30160;
  assign tmp30249 = l1 ? tmp29088 : tmp28497;
  assign tmp30251 = l1 ? 1 : tmp28741;
  assign tmp30252 = l1 ? tmp29615 : tmp27980;
  assign tmp30250 = ~(s0 ? tmp30251 : tmp30252);
  assign tmp30248 = s1 ? tmp30249 : tmp30250;
  assign tmp30255 = l1 ? tmp28835 : tmp28741;
  assign tmp30256 = ~(l1 ? tmp29620 : tmp28485);
  assign tmp30254 = s0 ? tmp30255 : tmp30256;
  assign tmp30258 = s0 ? tmp30255 : tmp27750;
  assign tmp30260 = l1 ? tmp29620 : tmp28485;
  assign tmp30261 = l1 ? tmp29620 : tmp28497;
  assign tmp30259 = ~(s0 ? tmp30260 : tmp30261);
  assign tmp30257 = s1 ? tmp30258 : tmp30259;
  assign tmp30253 = ~(s2 ? tmp30254 : tmp30257);
  assign tmp30247 = s3 ? tmp30248 : tmp30253;
  assign tmp30266 = l1 ? 1 : tmp27980;
  assign tmp30265 = s0 ? tmp30266 : tmp27750;
  assign tmp30267 = ~(s0 ? tmp30261 : tmp30260);
  assign tmp30264 = s1 ? tmp30265 : tmp30267;
  assign tmp30269 = s0 ? tmp30249 : tmp27791;
  assign tmp30270 = ~(s0 ? tmp28897 : tmp27750);
  assign tmp30268 = ~(s1 ? tmp30269 : tmp30270);
  assign tmp30263 = s2 ? tmp30264 : tmp30268;
  assign tmp30273 = s0 ? tmp28897 : tmp30251;
  assign tmp30274 = s0 ? tmp27750 : tmp30186;
  assign tmp30272 = s1 ? tmp30273 : tmp30274;
  assign tmp30277 = l1 ? tmp27490 : tmp28485;
  assign tmp30276 = s0 ? tmp30260 : tmp30277;
  assign tmp30278 = s0 ? tmp30093 : tmp30260;
  assign tmp30275 = ~(s1 ? tmp30276 : tmp30278);
  assign tmp30271 = s2 ? tmp30272 : tmp30275;
  assign tmp30262 = ~(s3 ? tmp30263 : tmp30271);
  assign tmp30246 = s4 ? tmp30247 : tmp30262;
  assign tmp30284 = s0 ? tmp30252 : tmp27750;
  assign tmp30283 = s1 ? tmp30284 : tmp27750;
  assign tmp30287 = l1 ? tmp29615 : tmp28014;
  assign tmp30286 = s0 ? tmp27750 : tmp30287;
  assign tmp30288 = ~(s0 ? tmp30277 : tmp27791);
  assign tmp30285 = s1 ? tmp30286 : tmp30288;
  assign tmp30282 = s2 ? tmp30283 : tmp30285;
  assign tmp30292 = l1 ? tmp27897 : tmp28741;
  assign tmp30291 = s0 ? tmp27750 : tmp30292;
  assign tmp30294 = ~(l1 ? tmp27490 : tmp28525);
  assign tmp30293 = s0 ? tmp27750 : tmp30294;
  assign tmp30290 = s1 ? tmp30291 : tmp30293;
  assign tmp30297 = l1 ? tmp29620 : tmp28525;
  assign tmp30296 = s0 ? tmp30297 : tmp30093;
  assign tmp30295 = ~(s1 ? tmp30200 : tmp30296);
  assign tmp30289 = s2 ? tmp30290 : tmp30295;
  assign tmp30281 = s3 ? tmp30282 : tmp30289;
  assign tmp30302 = l1 ? tmp29620 : tmp28531;
  assign tmp30301 = s0 ? tmp27858 : tmp30302;
  assign tmp30300 = s1 ? tmp30301 : tmp28896;
  assign tmp30304 = s0 ? tmp27750 : tmp28897;
  assign tmp30306 = l1 ? 1 : tmp28014;
  assign tmp30305 = s0 ? tmp30306 : tmp27750;
  assign tmp30303 = ~(s1 ? tmp30304 : tmp30305);
  assign tmp30299 = s2 ? tmp30300 : tmp30303;
  assign tmp30310 = ~(l1 ? tmp27490 : tmp28531);
  assign tmp30309 = s0 ? tmp30306 : tmp30310;
  assign tmp30312 = ~(l1 ? tmp27490 : tmp27820);
  assign tmp30311 = s0 ? tmp28897 : tmp30312;
  assign tmp30308 = s1 ? tmp30309 : tmp30311;
  assign tmp30307 = ~(s2 ? tmp30308 : tmp30213);
  assign tmp30298 = ~(s3 ? tmp30299 : tmp30307);
  assign tmp30280 = s4 ? tmp30281 : tmp30298;
  assign tmp30317 = s0 ? tmp30093 : tmp29230;
  assign tmp30319 = ~(l1 ? tmp27504 : tmp27971);
  assign tmp30318 = s0 ? tmp29230 : tmp30319;
  assign tmp30316 = s1 ? tmp30317 : tmp30318;
  assign tmp30322 = l1 ? tmp27504 : tmp27971;
  assign tmp30321 = s0 ? tmp30322 : tmp27750;
  assign tmp30320 = ~(s1 ? tmp30321 : tmp27750);
  assign tmp30315 = s2 ? tmp30316 : tmp30320;
  assign tmp30325 = s0 ? tmp27750 : tmp27640;
  assign tmp30324 = s1 ? tmp30325 : tmp30223;
  assign tmp30327 = s0 ? 1 : tmp29958;
  assign tmp30326 = ~(s1 ? tmp30225 : tmp30327);
  assign tmp30323 = ~(s2 ? tmp30324 : tmp30326);
  assign tmp30314 = s3 ? tmp30315 : tmp30323;
  assign tmp30331 = s0 ? tmp27640 : tmp28074;
  assign tmp30330 = s1 ? tmp30331 : tmp30232;
  assign tmp30334 = ~(l1 ? tmp27897 : tmp28014);
  assign tmp30333 = s0 ? tmp29230 : tmp30334;
  assign tmp30332 = ~(s1 ? tmp30333 : tmp27791);
  assign tmp30329 = s2 ? tmp30330 : tmp30332;
  assign tmp30337 = s0 ? tmp30322 : tmp28210;
  assign tmp30338 = ~(s0 ? tmp28196 : tmp28115);
  assign tmp30336 = s1 ? tmp30337 : tmp30338;
  assign tmp30339 = ~(s1 ? tmp30327 : tmp30242);
  assign tmp30335 = s2 ? tmp30336 : tmp30339;
  assign tmp30328 = ~(s3 ? tmp30329 : tmp30335);
  assign tmp30313 = ~(s4 ? tmp30314 : tmp30328);
  assign tmp30279 = ~(s5 ? tmp30280 : tmp30313);
  assign tmp30245 = s6 ? tmp30246 : tmp30279;
  assign tmp30244 = s7 ? tmp30245 : tmp27495;
  assign tmp30243 = s8 ? tmp30160 : tmp30244;
  assign tmp30058 = s9 ? tmp30059 : tmp30243;
  assign tmp30341 = s8 ? tmp30160 : tmp30161;
  assign tmp30340 = s9 ? tmp30341 : tmp27495;
  assign tmp30057 = s10 ? tmp30058 : tmp30340;
  assign tmp30350 = l1 ? tmp28835 : tmp29615;
  assign tmp30351 = s0 ? 1 : tmp29623;
  assign tmp30349 = s1 ? tmp30350 : tmp30351;
  assign tmp30355 = l1 ? tmp28835 : tmp27615;
  assign tmp30354 = s0 ? 1 : tmp30355;
  assign tmp30356 = s0 ? tmp29623 : tmp30355;
  assign tmp30353 = s1 ? tmp30354 : tmp30356;
  assign tmp30357 = s1 ? tmp29625 : tmp30355;
  assign tmp30352 = s2 ? tmp30353 : tmp30357;
  assign tmp30348 = s3 ? tmp30349 : tmp30352;
  assign tmp30360 = s1 ? 1 : tmp30355;
  assign tmp30362 = s0 ? tmp30350 : 1;
  assign tmp30361 = s1 ? tmp30362 : 1;
  assign tmp30359 = s2 ? tmp30360 : tmp30361;
  assign tmp30365 = s0 ? 1 : tmp27838;
  assign tmp30364 = s1 ? 1 : tmp30365;
  assign tmp30368 = l1 ? tmp27760 : tmp27615;
  assign tmp30367 = s0 ? tmp30355 : tmp30368;
  assign tmp30369 = s0 ? tmp27838 : tmp30355;
  assign tmp30366 = s1 ? tmp30367 : tmp30369;
  assign tmp30363 = s2 ? tmp30364 : tmp30366;
  assign tmp30358 = s3 ? tmp30359 : tmp30363;
  assign tmp30347 = s4 ? tmp30348 : tmp30358;
  assign tmp30374 = s1 ? tmp29625 : 1;
  assign tmp30376 = s0 ? tmp30368 : 1;
  assign tmp30375 = s1 ? tmp30351 : tmp30376;
  assign tmp30373 = s2 ? tmp30374 : tmp30375;
  assign tmp30381 = l2 ? tmp27615 : tmp27506;
  assign tmp30380 = l1 ? tmp27760 : tmp30381;
  assign tmp30379 = s0 ? 1 : tmp30380;
  assign tmp30378 = s1 ? tmp29652 : tmp30379;
  assign tmp30383 = s0 ? tmp27838 : tmp27588;
  assign tmp30385 = l1 ? tmp28835 : tmp30381;
  assign tmp30386 = l1 ? tmp27760 : tmp27506;
  assign tmp30384 = s0 ? tmp30385 : tmp30386;
  assign tmp30382 = s1 ? tmp30383 : tmp30384;
  assign tmp30377 = s2 ? tmp30378 : tmp30382;
  assign tmp30372 = s3 ? tmp30373 : tmp30377;
  assign tmp30391 = l1 ? tmp28835 : tmp27897;
  assign tmp30390 = s0 ? tmp27838 : tmp30391;
  assign tmp30389 = s1 ? tmp30390 : 1;
  assign tmp30388 = s2 ? tmp30389 : 1;
  assign tmp30394 = s0 ? 1 : tmp27897;
  assign tmp30395 = s0 ? 1 : tmp30386;
  assign tmp30393 = s1 ? tmp30394 : tmp30395;
  assign tmp30397 = s0 ? tmp27838 : tmp28446;
  assign tmp30396 = s1 ? tmp28446 : tmp30397;
  assign tmp30392 = s2 ? tmp30393 : tmp30396;
  assign tmp30387 = s3 ? tmp30388 : tmp30392;
  assign tmp30371 = s4 ? tmp30372 : tmp30387;
  assign tmp30402 = s0 ? tmp30380 : tmp27588;
  assign tmp30401 = s1 ? tmp30402 : tmp28715;
  assign tmp30403 = s1 ? tmp28236 : 1;
  assign tmp30400 = s2 ? tmp30401 : tmp30403;
  assign tmp30407 = ~(l1 ? tmp27495 : tmp27490);
  assign tmp30406 = s0 ? 1 : tmp30407;
  assign tmp30408 = ~(s0 ? tmp27532 : tmp27495);
  assign tmp30405 = s1 ? tmp30406 : tmp30408;
  assign tmp30411 = ~(l1 ? tmp27504 : tmp27506);
  assign tmp30410 = s0 ? tmp27495 : tmp30411;
  assign tmp30412 = ~(s0 ? tmp27838 : 1);
  assign tmp30409 = ~(s1 ? tmp30410 : tmp30412);
  assign tmp30404 = s2 ? tmp30405 : tmp30409;
  assign tmp30399 = s3 ? tmp30400 : tmp30404;
  assign tmp30416 = s0 ? 1 : tmp27836;
  assign tmp30417 = s0 ? tmp27836 : tmp27838;
  assign tmp30415 = s1 ? tmp30416 : tmp30417;
  assign tmp30420 = l1 ? tmp27760 : 1;
  assign tmp30419 = s0 ? tmp27588 : tmp30420;
  assign tmp30418 = s1 ? tmp30419 : 1;
  assign tmp30414 = s2 ? tmp30415 : tmp30418;
  assign tmp30424 = l1 ? tmp27504 : tmp27898;
  assign tmp30423 = s0 ? tmp27504 : tmp30424;
  assign tmp30426 = ~(l1 ? tmp27760 : tmp27897);
  assign tmp30425 = ~(s0 ? tmp27495 : tmp30426);
  assign tmp30422 = s1 ? tmp30423 : tmp30425;
  assign tmp30428 = s0 ? tmp27838 : 1;
  assign tmp30429 = ~(s0 ? tmp27532 : tmp29728);
  assign tmp30427 = s1 ? tmp30428 : tmp30429;
  assign tmp30421 = s2 ? tmp30422 : tmp30427;
  assign tmp30413 = s3 ? tmp30414 : tmp30421;
  assign tmp30398 = s4 ? tmp30399 : tmp30413;
  assign tmp30370 = s5 ? tmp30371 : tmp30398;
  assign tmp30346 = s6 ? tmp30347 : tmp30370;
  assign tmp30345 = s7 ? tmp30346 : tmp27575;
  assign tmp30434 = s1 ? tmp30355 : tmp30351;
  assign tmp30433 = s3 ? tmp30434 : tmp30352;
  assign tmp30438 = s0 ? tmp30355 : 1;
  assign tmp30437 = s1 ? tmp30438 : 1;
  assign tmp30436 = s2 ? tmp30360 : tmp30437;
  assign tmp30435 = s3 ? tmp30436 : tmp30363;
  assign tmp30432 = s4 ? tmp30433 : tmp30435;
  assign tmp30444 = s0 ? tmp27838 : tmp27697;
  assign tmp30443 = s1 ? tmp30444 : tmp30384;
  assign tmp30442 = s2 ? tmp30378 : tmp30443;
  assign tmp30441 = s3 ? tmp30373 : tmp30442;
  assign tmp30448 = s0 ? 1 : tmp27909;
  assign tmp30447 = s1 ? tmp30448 : tmp30395;
  assign tmp30450 = s0 ? tmp27838 : tmp27640;
  assign tmp30449 = s1 ? tmp27640 : tmp30450;
  assign tmp30446 = s2 ? tmp30447 : tmp30449;
  assign tmp30445 = s3 ? tmp30388 : tmp30446;
  assign tmp30440 = s4 ? tmp30441 : tmp30445;
  assign tmp30455 = s0 ? tmp30380 : tmp27697;
  assign tmp30454 = s1 ? tmp30455 : tmp27868;
  assign tmp30456 = s1 ? tmp27842 : 1;
  assign tmp30453 = s2 ? tmp30454 : tmp30456;
  assign tmp30460 = ~(l1 ? 1 : tmp27490);
  assign tmp30459 = s0 ? 1 : tmp30460;
  assign tmp30461 = ~(s0 ? tmp27642 : 1);
  assign tmp30458 = s1 ? tmp30459 : tmp30461;
  assign tmp30463 = s0 ? 1 : tmp30411;
  assign tmp30462 = ~(s1 ? tmp30463 : tmp30412);
  assign tmp30457 = s2 ? tmp30458 : tmp30462;
  assign tmp30452 = s3 ? tmp30453 : tmp30457;
  assign tmp30467 = s0 ? tmp27697 : tmp30420;
  assign tmp30466 = s1 ? tmp30467 : 1;
  assign tmp30465 = s2 ? tmp30415 : tmp30466;
  assign tmp30471 = l1 ? tmp27504 : tmp28495;
  assign tmp30470 = s0 ? tmp27836 : tmp30471;
  assign tmp30472 = ~(s0 ? 1 : tmp30426);
  assign tmp30469 = s1 ? tmp30470 : tmp30472;
  assign tmp30474 = ~(s0 ? tmp27642 : tmp29728);
  assign tmp30473 = s1 ? tmp30428 : tmp30474;
  assign tmp30468 = s2 ? tmp30469 : tmp30473;
  assign tmp30464 = s3 ? tmp30465 : tmp30468;
  assign tmp30451 = s4 ? tmp30452 : tmp30464;
  assign tmp30439 = s5 ? tmp30440 : tmp30451;
  assign tmp30431 = s6 ? tmp30432 : tmp30439;
  assign tmp30430 = s7 ? tmp30431 : tmp27575;
  assign tmp30344 = s8 ? tmp30345 : tmp30430;
  assign tmp30482 = l2 ? 1 : tmp29979;
  assign tmp30481 = l1 ? tmp28835 : tmp30482;
  assign tmp30483 = s0 ? tmp27750 : tmp29761;
  assign tmp30480 = s1 ? tmp30481 : tmp30483;
  assign tmp30488 = l2 ? tmp27615 : tmp29979;
  assign tmp30487 = l1 ? tmp28835 : tmp30488;
  assign tmp30486 = s0 ? tmp27750 : tmp30487;
  assign tmp30489 = s0 ? tmp29761 : tmp30487;
  assign tmp30485 = s1 ? tmp30486 : tmp30489;
  assign tmp30490 = s1 ? tmp29763 : tmp30487;
  assign tmp30484 = s2 ? tmp30485 : tmp30490;
  assign tmp30479 = s3 ? tmp30480 : tmp30484;
  assign tmp30493 = s1 ? tmp27750 : tmp30487;
  assign tmp30495 = s0 ? tmp30481 : tmp27750;
  assign tmp30494 = s1 ? tmp30495 : tmp27750;
  assign tmp30492 = s2 ? tmp30493 : tmp30494;
  assign tmp30497 = s1 ? tmp27750 : tmp27793;
  assign tmp30500 = l1 ? tmp27760 : tmp30488;
  assign tmp30499 = s0 ? tmp30487 : tmp30500;
  assign tmp30501 = s0 ? tmp27574 : tmp30487;
  assign tmp30498 = s1 ? tmp30499 : tmp30501;
  assign tmp30496 = s2 ? tmp30497 : tmp30498;
  assign tmp30491 = s3 ? tmp30492 : tmp30496;
  assign tmp30478 = s4 ? tmp30479 : tmp30491;
  assign tmp30506 = s1 ? tmp29763 : tmp27750;
  assign tmp30508 = s0 ? tmp30500 : tmp27750;
  assign tmp30507 = s1 ? tmp30483 : tmp30508;
  assign tmp30505 = s2 ? tmp30506 : tmp30507;
  assign tmp30513 = l2 ? tmp27615 : tmp28324;
  assign tmp30512 = l1 ? tmp27760 : tmp30513;
  assign tmp30511 = s0 ? tmp27750 : tmp30512;
  assign tmp30510 = s1 ? tmp29790 : tmp30511;
  assign tmp30515 = s0 ? tmp27574 : tmp27697;
  assign tmp30517 = l1 ? tmp28835 : tmp30513;
  assign tmp30518 = l1 ? tmp27760 : tmp27553;
  assign tmp30516 = s0 ? tmp30517 : tmp30518;
  assign tmp30514 = s1 ? tmp30515 : tmp30516;
  assign tmp30509 = s2 ? tmp30510 : tmp30514;
  assign tmp30504 = s3 ? tmp30505 : tmp30509;
  assign tmp30523 = l1 ? tmp28835 : tmp28323;
  assign tmp30522 = s0 ? tmp27574 : tmp30523;
  assign tmp30521 = s1 ? tmp30522 : tmp27750;
  assign tmp30520 = s2 ? tmp30521 : tmp27750;
  assign tmp30526 = s0 ? tmp27750 : tmp28338;
  assign tmp30527 = s0 ? tmp27750 : tmp30518;
  assign tmp30525 = s1 ? tmp30526 : tmp30527;
  assign tmp30529 = s0 ? tmp27574 : tmp27640;
  assign tmp30528 = s1 ? tmp27640 : tmp30529;
  assign tmp30524 = s2 ? tmp30525 : tmp30528;
  assign tmp30519 = s3 ? tmp30520 : tmp30524;
  assign tmp30503 = s4 ? tmp30504 : tmp30519;
  assign tmp30534 = s0 ? tmp30512 : tmp27697;
  assign tmp30533 = s1 ? tmp30534 : tmp27778;
  assign tmp30532 = s2 ? tmp30533 : tmp27802;
  assign tmp30538 = ~(l1 ? 1 : tmp28080);
  assign tmp30537 = s0 ? tmp27750 : tmp30538;
  assign tmp30536 = s1 ? tmp30537 : tmp29236;
  assign tmp30541 = ~(l1 ? tmp27504 : tmp27553);
  assign tmp30540 = s0 ? 1 : tmp30541;
  assign tmp30542 = ~(s0 ? tmp27574 : tmp27750);
  assign tmp30539 = ~(s1 ? tmp30540 : tmp30542);
  assign tmp30535 = s2 ? tmp30536 : tmp30539;
  assign tmp30531 = s3 ? tmp30532 : tmp30535;
  assign tmp30546 = s0 ? tmp27743 : tmp27574;
  assign tmp30545 = s1 ? tmp27799 : tmp30546;
  assign tmp30549 = l1 ? tmp27760 : tmp27744;
  assign tmp30548 = s0 ? tmp27697 : tmp30549;
  assign tmp30547 = s1 ? tmp30548 : tmp27750;
  assign tmp30544 = s2 ? tmp30545 : tmp30547;
  assign tmp30553 = l1 ? tmp27504 : tmp30049;
  assign tmp30552 = s0 ? tmp27743 : tmp30553;
  assign tmp30555 = ~(l1 ? tmp27760 : tmp27553);
  assign tmp30554 = ~(s0 ? 1 : tmp30555);
  assign tmp30551 = s1 ? tmp30552 : tmp30554;
  assign tmp30557 = s0 ? tmp27574 : tmp27750;
  assign tmp30558 = ~(s0 ? tmp29218 : tmp29816);
  assign tmp30556 = s1 ? tmp30557 : tmp30558;
  assign tmp30550 = s2 ? tmp30551 : tmp30556;
  assign tmp30543 = s3 ? tmp30544 : tmp30550;
  assign tmp30530 = s4 ? tmp30531 : tmp30543;
  assign tmp30502 = s5 ? tmp30503 : tmp30530;
  assign tmp30477 = s6 ? tmp30478 : tmp30502;
  assign tmp30476 = s7 ? tmp30477 : tmp27575;
  assign tmp30475 = s8 ? tmp30430 : tmp30476;
  assign tmp30343 = s9 ? tmp30344 : tmp30475;
  assign tmp30560 = s8 ? tmp30430 : tmp30431;
  assign tmp30559 = s9 ? tmp30560 : tmp27575;
  assign tmp30342 = ~(s10 ? tmp30343 : tmp30559);
  assign tmp30056 = s12 ? tmp30057 : tmp30342;
  assign tmp29602 = s13 ? tmp29603 : tmp30056;
  assign tmp30572 = ~(l1 ? tmp28934 : tmp28490);
  assign tmp30571 = s0 ? tmp28643 : tmp30572;
  assign tmp30570 = s1 ? tmp28643 : tmp30571;
  assign tmp30575 = ~(l1 ? tmp28641 : tmp28643);
  assign tmp30574 = s0 ? tmp29333 : tmp30575;
  assign tmp30577 = s0 ? tmp29333 : 0;
  assign tmp30576 = s1 ? tmp30577 : tmp30575;
  assign tmp30573 = ~(s2 ? tmp30574 : tmp30576);
  assign tmp30569 = s3 ? tmp30570 : tmp30573;
  assign tmp30580 = s1 ? tmp29333 : tmp30575;
  assign tmp30581 = ~(s0 ? tmp28643 : 1);
  assign tmp30579 = s2 ? tmp30580 : tmp30581;
  assign tmp30584 = s0 ? 1 : tmp30067;
  assign tmp30583 = s1 ? tmp28643 : tmp30584;
  assign tmp30587 = l1 ? tmp28641 : tmp28643;
  assign tmp30588 = l1 ? tmp28678 : tmp28643;
  assign tmp30586 = s0 ? tmp30587 : tmp30588;
  assign tmp30590 = l1 ? tmp28661 : tmp28643;
  assign tmp30589 = s0 ? tmp30590 : tmp30587;
  assign tmp30585 = s1 ? tmp30586 : tmp30589;
  assign tmp30582 = ~(s2 ? tmp30583 : tmp30585);
  assign tmp30578 = ~(s3 ? tmp30579 : tmp30582);
  assign tmp30568 = s4 ? tmp30569 : tmp30578;
  assign tmp30597 = l1 ? tmp28934 : tmp28490;
  assign tmp30596 = s0 ? tmp30597 : 0;
  assign tmp30595 = s1 ? tmp30596 : tmp29333;
  assign tmp30600 = ~(l1 ? tmp28934 : tmp28525);
  assign tmp30599 = s0 ? 1 : tmp30600;
  assign tmp30601 = s0 ? tmp30588 : 1;
  assign tmp30598 = ~(s1 ? tmp30599 : tmp30601);
  assign tmp30594 = s2 ? tmp30595 : tmp30598;
  assign tmp30605 = ~(l1 ? tmp28938 : tmp28490);
  assign tmp30604 = s0 ? 1 : tmp30605;
  assign tmp30606 = s0 ? 1 : tmp30588;
  assign tmp30603 = s1 ? tmp30604 : tmp30606;
  assign tmp30607 = s1 ? tmp30590 : tmp30586;
  assign tmp30602 = ~(s2 ? tmp30603 : tmp30607);
  assign tmp30593 = s3 ? tmp30594 : tmp30602;
  assign tmp30611 = s0 ? tmp28643 : tmp30587;
  assign tmp30610 = s1 ? tmp30611 : tmp28693;
  assign tmp30613 = ~(l1 ? tmp28938 : tmp28525);
  assign tmp30612 = s1 ? tmp28693 : tmp30613;
  assign tmp30609 = s2 ? tmp30610 : tmp30612;
  assign tmp30617 = ~(l1 ? tmp28643 : tmp27505);
  assign tmp30616 = s0 ? tmp30119 : tmp30617;
  assign tmp30619 = ~(l1 ? tmp28678 : tmp28643);
  assign tmp30618 = s0 ? tmp27495 : tmp30619;
  assign tmp30615 = s1 ? tmp30616 : tmp30618;
  assign tmp30621 = s0 ? tmp30067 : 1;
  assign tmp30620 = ~(s1 ? 1 : tmp30621);
  assign tmp30614 = ~(s2 ? tmp30615 : tmp30620);
  assign tmp30608 = ~(s3 ? tmp30609 : tmp30614);
  assign tmp30592 = s4 ? tmp30593 : tmp30608;
  assign tmp30627 = ~(l1 ? tmp27517 : tmp27495);
  assign tmp30626 = s0 ? 1 : tmp30627;
  assign tmp30625 = s1 ? tmp30601 : tmp30626;
  assign tmp30629 = s0 ? tmp29880 : tmp28225;
  assign tmp30628 = ~(s1 ? tmp30629 : tmp29392);
  assign tmp30624 = s2 ? tmp30625 : tmp30628;
  assign tmp30633 = ~(l1 ? 1 : tmp28643);
  assign tmp30632 = s0 ? tmp27495 : tmp30633;
  assign tmp30631 = s1 ? tmp30632 : tmp30083;
  assign tmp30636 = l1 ? 1 : tmp27505;
  assign tmp30635 = s0 ? 1 : tmp30636;
  assign tmp30637 = s0 ? tmp30636 : tmp27575;
  assign tmp30634 = ~(s1 ? tmp30635 : tmp30637);
  assign tmp30630 = ~(s2 ? tmp30631 : tmp30634);
  assign tmp30623 = s3 ? tmp30624 : tmp30630;
  assign tmp30641 = s0 ? tmp27495 : tmp29880;
  assign tmp30643 = ~(l1 ? tmp28661 : tmp28643);
  assign tmp30642 = s0 ? tmp29880 : tmp30643;
  assign tmp30640 = s1 ? tmp30641 : tmp30642;
  assign tmp30646 = ~(l1 ? tmp28733 : tmp28525);
  assign tmp30645 = s0 ? 1 : tmp30646;
  assign tmp30644 = ~(s1 ? tmp30645 : tmp29398);
  assign tmp30639 = s2 ? tmp30640 : tmp30644;
  assign tmp30650 = l1 ? tmp27517 : tmp28490;
  assign tmp30649 = s0 ? tmp29880 : tmp30650;
  assign tmp30652 = l1 ? tmp28678 : tmp27505;
  assign tmp30651 = ~(s0 ? 1 : tmp30652);
  assign tmp30648 = s1 ? tmp30649 : tmp30651;
  assign tmp30654 = s0 ? tmp30067 : tmp30627;
  assign tmp30653 = ~(s1 ? tmp30637 : tmp30654);
  assign tmp30647 = s2 ? tmp30648 : tmp30653;
  assign tmp30638 = ~(s3 ? tmp30639 : tmp30647);
  assign tmp30622 = ~(s4 ? tmp30623 : tmp30638);
  assign tmp30591 = ~(s5 ? tmp30592 : tmp30622);
  assign tmp30567 = s6 ? tmp30568 : tmp30591;
  assign tmp30566 = s7 ? tmp30567 : tmp27575;
  assign tmp30660 = l1 ? tmp28643 : tmp27490;
  assign tmp30662 = l1 ? tmp28741 : tmp27490;
  assign tmp30661 = s0 ? tmp27996 : tmp30662;
  assign tmp30659 = s1 ? tmp30660 : tmp30661;
  assign tmp30665 = l1 ? tmp28641 : tmp27490;
  assign tmp30664 = s0 ? tmp27979 : tmp30665;
  assign tmp30667 = s0 ? tmp27979 : tmp27642;
  assign tmp30666 = s1 ? tmp30667 : tmp30665;
  assign tmp30663 = s2 ? tmp30664 : tmp30666;
  assign tmp30658 = s3 ? tmp30659 : tmp30663;
  assign tmp30670 = s1 ? tmp27979 : tmp30665;
  assign tmp30672 = s0 ? tmp30660 : 1;
  assign tmp30671 = s1 ? tmp30672 : tmp27995;
  assign tmp30669 = s2 ? tmp30670 : tmp30671;
  assign tmp30675 = s0 ? 1 : tmp27642;
  assign tmp30674 = s1 ? tmp27996 : tmp30675;
  assign tmp30678 = l1 ? tmp28678 : tmp27490;
  assign tmp30677 = s0 ? tmp30665 : tmp30678;
  assign tmp30680 = l1 ? tmp27891 : tmp27490;
  assign tmp30679 = s0 ? tmp30680 : tmp30665;
  assign tmp30676 = s1 ? tmp30677 : tmp30679;
  assign tmp30673 = s2 ? tmp30674 : tmp30676;
  assign tmp30668 = s3 ? tmp30669 : tmp30673;
  assign tmp30657 = s4 ? tmp30658 : tmp30668;
  assign tmp30686 = s0 ? tmp30662 : 1;
  assign tmp30685 = s1 ? tmp30686 : tmp28009;
  assign tmp30689 = l1 ? tmp28741 : tmp27497;
  assign tmp30688 = s0 ? 1 : tmp30689;
  assign tmp30690 = s0 ? tmp30678 : tmp27642;
  assign tmp30687 = s1 ? tmp30688 : tmp30690;
  assign tmp30684 = s2 ? tmp30685 : tmp30687;
  assign tmp30693 = s0 ? tmp27642 : tmp27979;
  assign tmp30695 = l1 ? tmp29088 : tmp27490;
  assign tmp30694 = s0 ? tmp27642 : tmp30695;
  assign tmp30692 = s1 ? tmp30693 : tmp30694;
  assign tmp30696 = s1 ? tmp30680 : tmp30677;
  assign tmp30691 = s2 ? tmp30692 : tmp30696;
  assign tmp30683 = s3 ? tmp30684 : tmp30691;
  assign tmp30700 = s0 ? tmp27490 : tmp30665;
  assign tmp30699 = s1 ? tmp30700 : tmp28029;
  assign tmp30702 = l1 ? tmp27980 : tmp27497;
  assign tmp30701 = s1 ? tmp28029 : tmp30702;
  assign tmp30698 = s2 ? tmp30699 : tmp30701;
  assign tmp30706 = ~(l1 ? tmp28643 : tmp28226);
  assign tmp30705 = s0 ? tmp27858 : tmp30706;
  assign tmp30707 = ~(s0 ? tmp27697 : tmp30695);
  assign tmp30704 = s1 ? tmp30705 : tmp30707;
  assign tmp30709 = s0 ? tmp27642 : 1;
  assign tmp30708 = ~(s1 ? 1 : tmp30709);
  assign tmp30703 = ~(s2 ? tmp30704 : tmp30708);
  assign tmp30697 = s3 ? tmp30698 : tmp30703;
  assign tmp30682 = s4 ? tmp30683 : tmp30697;
  assign tmp30714 = s0 ? tmp30695 : 1;
  assign tmp30713 = s1 ? tmp30714 : tmp29727;
  assign tmp30716 = s0 ? tmp27836 : tmp27858;
  assign tmp30715 = ~(s1 ? tmp30716 : tmp27964);
  assign tmp30712 = s2 ? tmp30713 : tmp30715;
  assign tmp30720 = l1 ? 1 : tmp28226;
  assign tmp30719 = s0 ? 1 : tmp30720;
  assign tmp30721 = s0 ? tmp30720 : 0;
  assign tmp30718 = ~(s1 ? tmp30719 : tmp30721);
  assign tmp30717 = ~(s2 ? tmp30458 : tmp30718);
  assign tmp30711 = s3 ? tmp30712 : tmp30717;
  assign tmp30726 = ~(l1 ? tmp27891 : tmp27490);
  assign tmp30725 = s0 ? tmp27836 : tmp30726;
  assign tmp30724 = s1 ? tmp30416 : tmp30725;
  assign tmp30729 = ~(l1 ? tmp28835 : tmp27820);
  assign tmp30728 = s0 ? 1 : tmp30729;
  assign tmp30727 = ~(s1 ? tmp30728 : tmp29477);
  assign tmp30723 = s2 ? tmp30724 : tmp30727;
  assign tmp30733 = l1 ? tmp29088 : tmp28226;
  assign tmp30732 = ~(s0 ? 1 : tmp30733);
  assign tmp30731 = s1 ? tmp30417 : tmp30732;
  assign tmp30735 = s0 ? tmp27642 : tmp29728;
  assign tmp30734 = ~(s1 ? tmp30721 : tmp30735);
  assign tmp30730 = s2 ? tmp30731 : tmp30734;
  assign tmp30722 = ~(s3 ? tmp30723 : tmp30730);
  assign tmp30710 = s4 ? tmp30711 : tmp30722;
  assign tmp30681 = s5 ? tmp30682 : tmp30710;
  assign tmp30656 = s6 ? tmp30657 : tmp30681;
  assign tmp30655 = s7 ? tmp30656 : tmp27575;
  assign tmp30565 = s8 ? tmp30566 : tmp30655;
  assign tmp30742 = l1 ? tmp28643 : tmp27980;
  assign tmp30744 = l1 ? tmp28741 : tmp27980;
  assign tmp30743 = s0 ? tmp28740 : tmp30744;
  assign tmp30741 = s1 ? tmp30742 : tmp30743;
  assign tmp30747 = s0 ? tmp29488 : tmp30587;
  assign tmp30749 = l1 ? tmp27980 : tmp28741;
  assign tmp30748 = s0 ? tmp30749 : tmp30587;
  assign tmp30746 = s1 ? tmp30747 : tmp30748;
  assign tmp30751 = s0 ? tmp30749 : tmp27750;
  assign tmp30753 = l1 ? tmp28641 : tmp27980;
  assign tmp30752 = s0 ? tmp30587 : tmp30753;
  assign tmp30750 = s1 ? tmp30751 : tmp30752;
  assign tmp30745 = s2 ? tmp30746 : tmp30750;
  assign tmp30740 = s3 ? tmp30741 : tmp30745;
  assign tmp30757 = s0 ? tmp27980 : tmp27784;
  assign tmp30758 = s0 ? tmp30753 : tmp30587;
  assign tmp30756 = s1 ? tmp30757 : tmp30758;
  assign tmp30760 = s0 ? tmp30742 : tmp27750;
  assign tmp30759 = s1 ? tmp30760 : tmp28853;
  assign tmp30755 = s2 ? tmp30756 : tmp30759;
  assign tmp30763 = s0 ? tmp27750 : tmp27642;
  assign tmp30762 = s1 ? tmp28857 : tmp30763;
  assign tmp30766 = l1 ? tmp27891 : tmp28643;
  assign tmp30765 = s0 ? tmp30766 : tmp30587;
  assign tmp30764 = s1 ? tmp30586 : tmp30765;
  assign tmp30761 = s2 ? tmp30762 : tmp30764;
  assign tmp30754 = s3 ? tmp30755 : tmp30761;
  assign tmp30739 = s4 ? tmp30740 : tmp30754;
  assign tmp30772 = s0 ? tmp30744 : tmp27750;
  assign tmp30771 = s1 ? tmp30772 : tmp29508;
  assign tmp30775 = l1 ? tmp28741 : tmp28014;
  assign tmp30774 = s0 ? tmp27750 : tmp30775;
  assign tmp30776 = s0 ? tmp30588 : tmp27750;
  assign tmp30773 = s1 ? tmp30774 : tmp30776;
  assign tmp30770 = s2 ? tmp30771 : tmp30773;
  assign tmp30779 = s0 ? tmp27750 : tmp30749;
  assign tmp30781 = l1 ? tmp29088 : tmp28643;
  assign tmp30780 = s0 ? tmp27750 : tmp30781;
  assign tmp30778 = s1 ? tmp30779 : tmp30780;
  assign tmp30783 = s0 ? tmp30766 : tmp27750;
  assign tmp30782 = s1 ? tmp30783 : tmp30586;
  assign tmp30777 = s2 ? tmp30778 : tmp30782;
  assign tmp30769 = s3 ? tmp30770 : tmp30777;
  assign tmp30787 = s0 ? tmp27490 : tmp30753;
  assign tmp30786 = s1 ? tmp30787 : tmp28885;
  assign tmp30790 = l1 ? tmp27980 : tmp28014;
  assign tmp30789 = s0 ? tmp30790 : tmp27784;
  assign tmp30788 = s1 ? tmp28885 : tmp30789;
  assign tmp30785 = s2 ? tmp30786 : tmp30788;
  assign tmp30794 = ~(l1 ? tmp28643 : tmp27980);
  assign tmp30793 = s0 ? tmp28546 : tmp30794;
  assign tmp30795 = ~(s0 ? tmp28014 : tmp30695);
  assign tmp30792 = s1 ? tmp30793 : tmp30795;
  assign tmp30797 = s0 ? tmp27642 : tmp27750;
  assign tmp30796 = ~(s1 ? tmp27750 : tmp30797);
  assign tmp30791 = ~(s2 ? tmp30792 : tmp30796);
  assign tmp30784 = s3 ? tmp30785 : tmp30791;
  assign tmp30768 = s4 ? tmp30769 : tmp30784;
  assign tmp30802 = s0 ? tmp30781 : tmp27750;
  assign tmp30804 = ~(l1 ? tmp27504 : tmp28497);
  assign tmp30803 = s0 ? tmp27750 : tmp30804;
  assign tmp30801 = s1 ? tmp30802 : tmp30803;
  assign tmp30807 = l1 ? tmp27504 : tmp28497;
  assign tmp30806 = s0 ? tmp30807 : tmp29230;
  assign tmp30805 = ~(s1 ? tmp30806 : tmp29532);
  assign tmp30800 = s2 ? tmp30801 : tmp30805;
  assign tmp30810 = ~(s0 ? tmp27642 : tmp27750);
  assign tmp30809 = s1 ? tmp30459 : tmp30810;
  assign tmp30812 = s0 ? tmp27750 : tmp30720;
  assign tmp30811 = ~(s1 ? tmp30812 : tmp30721);
  assign tmp30808 = ~(s2 ? tmp30809 : tmp30811);
  assign tmp30799 = s3 ? tmp30800 : tmp30808;
  assign tmp30817 = ~(l1 ? tmp27891 : tmp28643);
  assign tmp30816 = s0 ? tmp27836 : tmp30817;
  assign tmp30815 = s1 ? tmp30416 : tmp30816;
  assign tmp30820 = ~(l1 ? tmp28835 : tmp28531);
  assign tmp30819 = s0 ? tmp27750 : tmp30820;
  assign tmp30818 = ~(s1 ? tmp30819 : tmp29538);
  assign tmp30814 = s2 ? tmp30815 : tmp30818;
  assign tmp30823 = s0 ? tmp30807 : tmp27838;
  assign tmp30824 = ~(s0 ? tmp27750 : tmp30733);
  assign tmp30822 = s1 ? tmp30823 : tmp30824;
  assign tmp30821 = s2 ? tmp30822 : tmp30734;
  assign tmp30813 = ~(s3 ? tmp30814 : tmp30821);
  assign tmp30798 = s4 ? tmp30799 : tmp30813;
  assign tmp30767 = s5 ? tmp30768 : tmp30798;
  assign tmp30738 = s6 ? tmp30739 : tmp30767;
  assign tmp30737 = s7 ? tmp30738 : tmp27575;
  assign tmp30736 = s8 ? tmp30655 : tmp30737;
  assign tmp30564 = s9 ? tmp30565 : tmp30736;
  assign tmp30832 = s0 ? tmp28743 : tmp30744;
  assign tmp30831 = s1 ? tmp30742 : tmp30832;
  assign tmp30835 = s0 ? tmp29549 : tmp30587;
  assign tmp30836 = s0 ? tmp27980 : tmp30587;
  assign tmp30834 = s1 ? tmp30835 : tmp30836;
  assign tmp30838 = s0 ? tmp27980 : 1;
  assign tmp30837 = s1 ? tmp30838 : tmp30752;
  assign tmp30833 = s2 ? tmp30834 : tmp30837;
  assign tmp30830 = s3 ? tmp30831 : tmp30833;
  assign tmp30842 = s0 ? tmp27980 : tmp27991;
  assign tmp30841 = s1 ? tmp30842 : tmp30758;
  assign tmp30844 = s0 ? tmp30742 : 1;
  assign tmp30843 = s1 ? tmp30844 : tmp28760;
  assign tmp30840 = s2 ? tmp30841 : tmp30843;
  assign tmp30846 = s1 ? tmp28764 : tmp30675;
  assign tmp30845 = s2 ? tmp30846 : tmp30764;
  assign tmp30839 = s3 ? tmp30840 : tmp30845;
  assign tmp30829 = s4 ? tmp30830 : tmp30839;
  assign tmp30852 = s0 ? tmp30744 : 1;
  assign tmp30851 = s1 ? tmp30852 : tmp29568;
  assign tmp30854 = s0 ? 1 : tmp30775;
  assign tmp30853 = s1 ? tmp30854 : tmp30601;
  assign tmp30850 = s2 ? tmp30851 : tmp30853;
  assign tmp30857 = s0 ? 1 : tmp27980;
  assign tmp30858 = s0 ? 1 : tmp30781;
  assign tmp30856 = s1 ? tmp30857 : tmp30858;
  assign tmp30860 = s0 ? tmp30766 : 1;
  assign tmp30859 = s1 ? tmp30860 : tmp30586;
  assign tmp30855 = s2 ? tmp30856 : tmp30859;
  assign tmp30849 = s3 ? tmp30850 : tmp30855;
  assign tmp30863 = s1 ? tmp30787 : tmp28792;
  assign tmp30865 = s0 ? tmp30790 : tmp27991;
  assign tmp30864 = s1 ? tmp28792 : tmp30865;
  assign tmp30862 = s2 ? tmp30863 : tmp30864;
  assign tmp30866 = ~(s2 ? tmp30792 : tmp30708);
  assign tmp30861 = s3 ? tmp30862 : tmp30866;
  assign tmp30848 = s4 ? tmp30849 : tmp30861;
  assign tmp30871 = s0 ? tmp30781 : 1;
  assign tmp30873 = ~(l1 ? tmp27504 : tmp27492);
  assign tmp30872 = s0 ? 1 : tmp30873;
  assign tmp30870 = s1 ? tmp30871 : tmp30872;
  assign tmp30875 = s0 ? tmp27703 : tmp28267;
  assign tmp30874 = ~(s1 ? tmp30875 : tmp28818);
  assign tmp30869 = s2 ? tmp30870 : tmp30874;
  assign tmp30868 = s3 ? tmp30869 : tmp30717;
  assign tmp30879 = s0 ? 1 : tmp30820;
  assign tmp30878 = ~(s1 ? tmp30879 : tmp29600);
  assign tmp30877 = s2 ? tmp30815 : tmp30878;
  assign tmp30882 = s0 ? tmp27703 : tmp27838;
  assign tmp30881 = s1 ? tmp30882 : tmp30732;
  assign tmp30880 = s2 ? tmp30881 : tmp30734;
  assign tmp30876 = ~(s3 ? tmp30877 : tmp30880);
  assign tmp30867 = s4 ? tmp30868 : tmp30876;
  assign tmp30847 = s5 ? tmp30848 : tmp30867;
  assign tmp30828 = s6 ? tmp30829 : tmp30847;
  assign tmp30827 = s7 ? tmp30828 : tmp27575;
  assign tmp30826 = s8 ? tmp30827 : tmp30828;
  assign tmp30825 = s9 ? tmp30826 : tmp27575;
  assign tmp30563 = s10 ? tmp30564 : tmp30825;
  assign tmp30891 = l1 ? tmp30069 : tmp28641;
  assign tmp30894 = l2 ? tmp27496 : tmp27487;
  assign tmp30893 = ~(l1 ? tmp30894 : tmp28665);
  assign tmp30892 = s0 ? tmp30067 : tmp30893;
  assign tmp30890 = s1 ? tmp30891 : tmp30892;
  assign tmp30897 = l1 ? tmp29442 : tmp28490;
  assign tmp30899 = l2 ? tmp27554 : tmp27615;
  assign tmp30898 = ~(l1 ? tmp30899 : tmp28641);
  assign tmp30896 = s0 ? tmp30897 : tmp30898;
  assign tmp30901 = s0 ? tmp30897 : 0;
  assign tmp30900 = s1 ? tmp30901 : tmp30898;
  assign tmp30895 = ~(s2 ? tmp30896 : tmp30900);
  assign tmp30889 = s3 ? tmp30890 : tmp30895;
  assign tmp30906 = l1 ? tmp27517 : tmp28665;
  assign tmp30905 = s0 ? tmp30906 : 0;
  assign tmp30904 = s1 ? tmp30905 : tmp30898;
  assign tmp30908 = s0 ? tmp30891 : 1;
  assign tmp30907 = ~(s1 ? tmp30908 : tmp30621);
  assign tmp30903 = s2 ? tmp30904 : tmp30907;
  assign tmp30910 = s1 ? tmp30067 : tmp30105;
  assign tmp30913 = l1 ? tmp30899 : tmp28641;
  assign tmp30915 = l2 ? tmp27554 : tmp27506;
  assign tmp30914 = l1 ? tmp30915 : tmp28641;
  assign tmp30912 = s0 ? tmp30913 : tmp30914;
  assign tmp30917 = l1 ? tmp30915 : tmp28661;
  assign tmp30916 = s0 ? tmp30917 : tmp30913;
  assign tmp30911 = s1 ? tmp30912 : tmp30916;
  assign tmp30909 = ~(s2 ? tmp30910 : tmp30911);
  assign tmp30902 = ~(s3 ? tmp30903 : tmp30909);
  assign tmp30888 = s4 ? tmp30889 : tmp30902;
  assign tmp30924 = l1 ? tmp30894 : tmp28665;
  assign tmp30923 = s0 ? tmp30924 : 0;
  assign tmp30926 = ~(l1 ? tmp27517 : tmp28490);
  assign tmp30925 = ~(s0 ? 1 : tmp30926);
  assign tmp30922 = s1 ? tmp30923 : tmp30925;
  assign tmp30929 = ~(l1 ? tmp30894 : tmp28685);
  assign tmp30928 = s0 ? 1 : tmp30929;
  assign tmp30930 = s0 ? tmp30914 : 1;
  assign tmp30927 = ~(s1 ? tmp30928 : tmp30930);
  assign tmp30921 = s2 ? tmp30922 : tmp30927;
  assign tmp30934 = ~(l1 ? tmp29414 : tmp28490);
  assign tmp30933 = s0 ? 1 : tmp30934;
  assign tmp30936 = l1 ? tmp30915 : tmp28678;
  assign tmp30935 = s0 ? 1 : tmp30936;
  assign tmp30932 = s1 ? tmp30933 : tmp30935;
  assign tmp30938 = s0 ? tmp30917 : tmp28248;
  assign tmp30940 = l1 ? tmp30899 : tmp28678;
  assign tmp30939 = s0 ? tmp30940 : tmp30936;
  assign tmp30937 = s1 ? tmp30938 : tmp30939;
  assign tmp30931 = ~(s2 ? tmp30932 : tmp30937);
  assign tmp30920 = s3 ? tmp30921 : tmp30931;
  assign tmp30945 = l1 ? tmp27504 : tmp28661;
  assign tmp30944 = s0 ? tmp30945 : tmp30940;
  assign tmp30943 = s1 ? tmp30944 : tmp30121;
  assign tmp30948 = l1 ? tmp27517 : tmp28685;
  assign tmp30947 = ~(s0 ? tmp30948 : 0);
  assign tmp30946 = s1 ? tmp30121 : tmp30947;
  assign tmp30942 = s2 ? tmp30943 : tmp30946;
  assign tmp30952 = ~(l1 ? tmp30915 : tmp28702);
  assign tmp30951 = s0 ? tmp30948 : tmp30952;
  assign tmp30953 = ~(s0 ? tmp28446 : tmp30936);
  assign tmp30950 = s1 ? tmp30951 : tmp30953;
  assign tmp30955 = s0 ? tmp30106 : 1;
  assign tmp30954 = ~(s1 ? 1 : tmp30955);
  assign tmp30949 = ~(s2 ? tmp30950 : tmp30954);
  assign tmp30941 = ~(s3 ? tmp30942 : tmp30949);
  assign tmp30919 = s4 ? tmp30920 : tmp30941;
  assign tmp30960 = s0 ? tmp30936 : tmp27504;
  assign tmp30961 = s0 ? tmp27504 : tmp27575;
  assign tmp30959 = s1 ? tmp30960 : tmp30961;
  assign tmp30964 = l1 ? tmp27517 : tmp27833;
  assign tmp30963 = s0 ? tmp27495 : tmp30964;
  assign tmp30965 = s0 ? tmp29880 : tmp30964;
  assign tmp30962 = ~(s1 ? tmp30963 : tmp30965);
  assign tmp30958 = s2 ? tmp30959 : tmp30962;
  assign tmp30967 = s1 ? tmp29902 : tmp29698;
  assign tmp30970 = ~(l1 ? tmp27504 : tmp27960);
  assign tmp30969 = s0 ? tmp28214 : tmp30970;
  assign tmp30972 = l1 ? tmp27504 : tmp27960;
  assign tmp30973 = ~(l1 ? tmp27517 : tmp28733);
  assign tmp30971 = ~(s0 ? tmp30972 : tmp30973);
  assign tmp30968 = s1 ? tmp30969 : tmp30971;
  assign tmp30966 = ~(s2 ? tmp30967 : tmp30968);
  assign tmp30957 = s3 ? tmp30958 : tmp30966;
  assign tmp30978 = l1 ? tmp27517 : tmp28733;
  assign tmp30977 = s0 ? tmp30978 : tmp29414;
  assign tmp30980 = ~(l1 ? tmp30915 : tmp28661);
  assign tmp30979 = s0 ? tmp29414 : tmp30980;
  assign tmp30976 = s1 ? tmp30977 : tmp30979;
  assign tmp30983 = ~(l1 ? tmp29414 : tmp28685);
  assign tmp30982 = s0 ? tmp27504 : tmp30983;
  assign tmp30984 = ~(s0 ? tmp30964 : tmp29880);
  assign tmp30981 = ~(s1 ? tmp30982 : tmp30984);
  assign tmp30975 = s2 ? tmp30976 : tmp30981;
  assign tmp30988 = l1 ? tmp29414 : 0;
  assign tmp30987 = s0 ? tmp27495 : tmp30988;
  assign tmp30989 = s0 ? tmp28214 : tmp30952;
  assign tmp30986 = s1 ? tmp30987 : tmp30989;
  assign tmp30991 = s0 ? tmp30972 : tmp30973;
  assign tmp30992 = s0 ? 1 : tmp27898;
  assign tmp30990 = ~(s1 ? tmp30991 : tmp30992);
  assign tmp30985 = s2 ? tmp30986 : tmp30990;
  assign tmp30974 = ~(s3 ? tmp30975 : tmp30985);
  assign tmp30956 = ~(s4 ? tmp30957 : tmp30974);
  assign tmp30918 = ~(s5 ? tmp30919 : tmp30956);
  assign tmp30887 = s6 ? tmp30888 : tmp30918;
  assign tmp30886 = s7 ? tmp30887 : tmp27575;
  assign tmp30998 = l1 ? tmp30069 : tmp28860;
  assign tmp31000 = l1 ? tmp27614 : tmp28860;
  assign tmp30999 = s0 ? tmp27642 : tmp31000;
  assign tmp30997 = s1 ? tmp30998 : tmp30999;
  assign tmp31003 = l1 ? tmp27488 : tmp27490;
  assign tmp31004 = l1 ? tmp30899 : tmp28860;
  assign tmp31002 = s0 ? tmp31003 : tmp31004;
  assign tmp31006 = s0 ? tmp31003 : tmp27642;
  assign tmp31005 = s1 ? tmp31006 : tmp31004;
  assign tmp31001 = s2 ? tmp31002 : tmp31005;
  assign tmp30996 = s3 ? tmp30997 : tmp31001;
  assign tmp31011 = l1 ? tmp27623 : tmp28860;
  assign tmp31010 = s0 ? tmp31011 : 1;
  assign tmp31009 = s1 ? tmp31010 : tmp31004;
  assign tmp31013 = s0 ? tmp30998 : 1;
  assign tmp31012 = s1 ? tmp31013 : tmp30709;
  assign tmp31008 = s2 ? tmp31009 : tmp31012;
  assign tmp31017 = l1 ? tmp27897 : tmp27891;
  assign tmp31016 = s0 ? 1 : tmp31017;
  assign tmp31015 = s1 ? tmp27642 : tmp31016;
  assign tmp31020 = l1 ? tmp30915 : tmp28860;
  assign tmp31019 = s0 ? tmp31004 : tmp31020;
  assign tmp31022 = l1 ? tmp27624 : tmp27891;
  assign tmp31021 = s0 ? tmp31022 : tmp31004;
  assign tmp31018 = s1 ? tmp31019 : tmp31021;
  assign tmp31014 = s2 ? tmp31015 : tmp31018;
  assign tmp31007 = s3 ? tmp31008 : tmp31014;
  assign tmp30995 = s4 ? tmp30996 : tmp31007;
  assign tmp31028 = s0 ? tmp31000 : 1;
  assign tmp31030 = l1 ? tmp27623 : tmp27490;
  assign tmp31029 = s0 ? 1 : tmp31030;
  assign tmp31027 = s1 ? tmp31028 : tmp31029;
  assign tmp31033 = l1 ? tmp27614 : tmp29088;
  assign tmp31032 = s0 ? 1 : tmp31033;
  assign tmp31034 = s0 ? tmp31020 : tmp27642;
  assign tmp31031 = s1 ? tmp31032 : tmp31034;
  assign tmp31026 = s2 ? tmp31027 : tmp31031;
  assign tmp31038 = ~(l1 ? tmp27496 : tmp27506);
  assign tmp31037 = s0 ? tmp27642 : tmp31038;
  assign tmp31040 = l1 ? tmp27624 : tmp29088;
  assign tmp31039 = s0 ? tmp27642 : tmp31040;
  assign tmp31036 = s1 ? tmp31037 : tmp31039;
  assign tmp31042 = s0 ? tmp31022 : tmp28248;
  assign tmp31044 = l1 ? tmp30899 : tmp29088;
  assign tmp31045 = l1 ? tmp30915 : tmp29088;
  assign tmp31043 = s0 ? tmp31044 : tmp31045;
  assign tmp31041 = s1 ? tmp31042 : tmp31043;
  assign tmp31035 = s2 ? tmp31036 : tmp31041;
  assign tmp31025 = s3 ? tmp31026 : tmp31035;
  assign tmp31050 = l1 ? tmp27504 : tmp27891;
  assign tmp31049 = s0 ? tmp31050 : tmp31044;
  assign tmp31048 = s1 ? tmp31049 : tmp27677;
  assign tmp31053 = l1 ? tmp27623 : tmp29088;
  assign tmp31052 = s0 ? tmp31053 : 1;
  assign tmp31051 = s1 ? tmp27677 : tmp31052;
  assign tmp31047 = s2 ? tmp31048 : tmp31051;
  assign tmp31057 = l1 ? tmp27504 : tmp28802;
  assign tmp31058 = ~(l1 ? tmp30915 : tmp28821);
  assign tmp31056 = s0 ? tmp31057 : tmp31058;
  assign tmp31059 = ~(s0 ? tmp27640 : tmp31040);
  assign tmp31055 = s1 ? tmp31056 : tmp31059;
  assign tmp31061 = s0 ? tmp31017 : 1;
  assign tmp31060 = ~(s1 ? 1 : tmp31061);
  assign tmp31054 = ~(s2 ? tmp31055 : tmp31060);
  assign tmp31046 = s3 ? tmp31047 : tmp31054;
  assign tmp31024 = s4 ? tmp31025 : tmp31046;
  assign tmp31066 = s0 ? tmp31040 : tmp27504;
  assign tmp31067 = s0 ? tmp27504 : 0;
  assign tmp31065 = s1 ? tmp31066 : tmp31067;
  assign tmp31069 = s0 ? 1 : tmp27819;
  assign tmp31070 = s0 ? tmp27836 : tmp27819;
  assign tmp31068 = ~(s1 ? tmp31069 : tmp31070);
  assign tmp31064 = s2 ? tmp31065 : tmp31068;
  assign tmp31072 = s1 ? tmp29954 : tmp29698;
  assign tmp31075 = ~(l1 ? tmp27504 : tmp27833);
  assign tmp31074 = s0 ? tmp28214 : tmp31075;
  assign tmp31077 = ~(l1 ? tmp27504 : tmp28835);
  assign tmp31076 = ~(s0 ? tmp27832 : tmp31077);
  assign tmp31073 = s1 ? tmp31074 : tmp31076;
  assign tmp31071 = ~(s2 ? tmp31072 : tmp31073);
  assign tmp31063 = s3 ? tmp31064 : tmp31071;
  assign tmp31082 = l1 ? tmp27504 : tmp28835;
  assign tmp31081 = s0 ? tmp31082 : tmp27560;
  assign tmp31084 = ~(l1 ? tmp27624 : tmp27891);
  assign tmp31083 = s0 ? tmp27560 : tmp31084;
  assign tmp31080 = s1 ? tmp31081 : tmp31083;
  assign tmp31087 = ~(l1 ? tmp27560 : tmp28802);
  assign tmp31086 = s0 ? tmp27504 : tmp31087;
  assign tmp31088 = ~(s0 ? tmp27819 : tmp27836);
  assign tmp31085 = ~(s1 ? tmp31086 : tmp31088);
  assign tmp31079 = s2 ? tmp31080 : tmp31085;
  assign tmp31091 = s0 ? 1 : tmp28275;
  assign tmp31093 = ~(l1 ? tmp27624 : tmp28821);
  assign tmp31092 = s0 ? tmp28214 : tmp31093;
  assign tmp31090 = s1 ? tmp31091 : tmp31092;
  assign tmp31095 = s0 ? tmp27832 : tmp31077;
  assign tmp31096 = s0 ? 1 : tmp28495;
  assign tmp31094 = ~(s1 ? tmp31095 : tmp31096);
  assign tmp31089 = s2 ? tmp31090 : tmp31094;
  assign tmp31078 = ~(s3 ? tmp31079 : tmp31089);
  assign tmp31062 = s4 ? tmp31063 : tmp31078;
  assign tmp31023 = s5 ? tmp31024 : tmp31062;
  assign tmp30994 = s6 ? tmp30995 : tmp31023;
  assign tmp30993 = s7 ? tmp30994 : tmp27575;
  assign tmp30885 = s8 ? tmp30886 : tmp30993;
  assign tmp31103 = l1 ? tmp30069 : tmp28741;
  assign tmp31105 = l1 ? tmp27614 : tmp28741;
  assign tmp31104 = s0 ? tmp30251 : tmp31105;
  assign tmp31102 = s1 ? tmp31103 : tmp31104;
  assign tmp31108 = l1 ? tmp27488 : tmp28741;
  assign tmp31107 = s0 ? tmp31108 : tmp30913;
  assign tmp31110 = s0 ? tmp31108 : tmp27750;
  assign tmp31112 = l1 ? tmp30899 : tmp28741;
  assign tmp31111 = s0 ? tmp30913 : tmp31112;
  assign tmp31109 = s1 ? tmp31110 : tmp31111;
  assign tmp31106 = s2 ? tmp31107 : tmp31109;
  assign tmp31101 = s3 ? tmp31102 : tmp31106;
  assign tmp31117 = l1 ? tmp27623 : tmp28741;
  assign tmp31116 = s0 ? tmp31117 : tmp27750;
  assign tmp31118 = s0 ? tmp31112 : tmp30913;
  assign tmp31115 = s1 ? tmp31116 : tmp31118;
  assign tmp31120 = s0 ? tmp31103 : tmp27750;
  assign tmp31119 = s1 ? tmp31120 : tmp28916;
  assign tmp31114 = s2 ? tmp31115 : tmp31119;
  assign tmp31124 = l1 ? tmp27897 : tmp28860;
  assign tmp31123 = s0 ? tmp27750 : tmp31124;
  assign tmp31122 = s1 ? tmp30273 : tmp31123;
  assign tmp31127 = l1 ? tmp27624 : tmp28641;
  assign tmp31126 = s0 ? tmp31127 : tmp30913;
  assign tmp31125 = s1 ? tmp30912 : tmp31126;
  assign tmp31121 = s2 ? tmp31122 : tmp31125;
  assign tmp31113 = s3 ? tmp31114 : tmp31121;
  assign tmp31100 = s4 ? tmp31101 : tmp31113;
  assign tmp31133 = s0 ? tmp31105 : tmp27750;
  assign tmp31135 = l1 ? tmp27623 : tmp27744;
  assign tmp31134 = s0 ? tmp27750 : tmp31135;
  assign tmp31132 = s1 ? tmp31133 : tmp31134;
  assign tmp31137 = s0 ? tmp27750 : tmp31105;
  assign tmp31138 = s0 ? tmp30914 : tmp27750;
  assign tmp31136 = s1 ? tmp31137 : tmp31138;
  assign tmp31131 = s2 ? tmp31132 : tmp31136;
  assign tmp31143 = ~(l2 ? tmp27488 : tmp27496);
  assign tmp31142 = ~(l1 ? tmp27496 : tmp31143);
  assign tmp31141 = s0 ? tmp27750 : tmp31142;
  assign tmp31144 = s0 ? tmp27750 : tmp31127;
  assign tmp31140 = s1 ? tmp31141 : tmp31144;
  assign tmp31146 = s0 ? tmp31127 : tmp28378;
  assign tmp31145 = s1 ? tmp31146 : tmp30912;
  assign tmp31139 = s2 ? tmp31140 : tmp31145;
  assign tmp31130 = s3 ? tmp31131 : tmp31139;
  assign tmp31151 = l1 ? tmp27504 : tmp28860;
  assign tmp31150 = s0 ? tmp31151 : tmp31112;
  assign tmp31149 = s1 ? tmp31150 : tmp30304;
  assign tmp31152 = s1 ? tmp30304 : tmp31116;
  assign tmp31148 = s2 ? tmp31149 : tmp31152;
  assign tmp31156 = l1 ? tmp27504 : tmp31143;
  assign tmp31157 = ~(l1 ? tmp30915 : tmp28741);
  assign tmp31155 = s0 ? tmp31156 : tmp31157;
  assign tmp31159 = l1 ? tmp27624 : tmp28860;
  assign tmp31158 = ~(s0 ? tmp28897 : tmp31159);
  assign tmp31154 = s1 ? tmp31155 : tmp31158;
  assign tmp31161 = s0 ? tmp31124 : tmp27750;
  assign tmp31160 = ~(s1 ? tmp27750 : tmp31161);
  assign tmp31153 = ~(s2 ? tmp31154 : tmp31160);
  assign tmp31147 = s3 ? tmp31148 : tmp31153;
  assign tmp31129 = s4 ? tmp31130 : tmp31147;
  assign tmp31166 = s0 ? tmp31127 : tmp27504;
  assign tmp31167 = s0 ? tmp27504 : tmp28515;
  assign tmp31165 = s1 ? tmp31166 : tmp31167;
  assign tmp31169 = s0 ? tmp28496 : tmp29217;
  assign tmp31170 = s0 ? tmp29180 : tmp29217;
  assign tmp31168 = ~(s1 ? tmp31169 : tmp31170);
  assign tmp31164 = s2 ? tmp31165 : tmp31168;
  assign tmp31173 = s0 ? tmp29180 : tmp27791;
  assign tmp31172 = s1 ? tmp31173 : tmp29838;
  assign tmp31176 = ~(l1 ? tmp27504 : tmp27739);
  assign tmp31175 = s0 ? tmp28342 : tmp31176;
  assign tmp31177 = ~(s0 ? tmp27738 : tmp29178);
  assign tmp31174 = s1 ? tmp31175 : tmp31177;
  assign tmp31171 = ~(s2 ? tmp31172 : tmp31174);
  assign tmp31163 = s3 ? tmp31164 : tmp31171;
  assign tmp31183 = l2 ? 1 : tmp27554;
  assign tmp31182 = l1 ? tmp27560 : tmp31183;
  assign tmp31181 = s0 ? tmp29180 : tmp31182;
  assign tmp31185 = ~(l1 ? tmp27624 : tmp28641);
  assign tmp31184 = s0 ? tmp31182 : tmp31185;
  assign tmp31180 = s1 ? tmp31181 : tmp31184;
  assign tmp31188 = ~(l1 ? tmp27560 : tmp31143);
  assign tmp31187 = s0 ? tmp27504 : tmp31188;
  assign tmp31189 = ~(s0 ? tmp29217 : tmp29180);
  assign tmp31186 = ~(s1 ? tmp31187 : tmp31189);
  assign tmp31179 = s2 ? tmp31180 : tmp31186;
  assign tmp31193 = l1 ? tmp27560 : tmp27809;
  assign tmp31192 = s0 ? tmp28496 : tmp31193;
  assign tmp31195 = ~(l1 ? tmp27624 : tmp27739);
  assign tmp31194 = s0 ? tmp28342 : tmp31195;
  assign tmp31191 = s1 ? tmp31192 : tmp31194;
  assign tmp31197 = s0 ? tmp27738 : tmp29178;
  assign tmp31199 = ~(l1 ? tmp27560 : tmp31183);
  assign tmp31198 = s0 ? tmp27750 : tmp31199;
  assign tmp31196 = ~(s1 ? tmp31197 : tmp31198);
  assign tmp31190 = s2 ? tmp31191 : tmp31196;
  assign tmp31178 = ~(s3 ? tmp31179 : tmp31190);
  assign tmp31162 = s4 ? tmp31163 : tmp31178;
  assign tmp31128 = s5 ? tmp31129 : tmp31162;
  assign tmp31099 = s6 ? tmp31100 : tmp31128;
  assign tmp31098 = s7 ? tmp31099 : tmp27575;
  assign tmp31097 = s8 ? tmp30993 : tmp31098;
  assign tmp30884 = s9 ? tmp30885 : tmp31097;
  assign tmp31207 = s0 ? tmp30166 : tmp31105;
  assign tmp31206 = s1 ? tmp31103 : tmp31207;
  assign tmp31210 = l1 ? tmp27488 : tmp27980;
  assign tmp31209 = s0 ? tmp31210 : tmp30913;
  assign tmp31212 = s0 ? tmp31210 : 1;
  assign tmp31211 = s1 ? tmp31212 : tmp31111;
  assign tmp31208 = s2 ? tmp31209 : tmp31211;
  assign tmp31205 = s3 ? tmp31206 : tmp31208;
  assign tmp31216 = s0 ? tmp31117 : 1;
  assign tmp31215 = s1 ? tmp31216 : tmp31118;
  assign tmp31218 = s0 ? tmp31103 : 1;
  assign tmp31217 = s1 ? tmp31218 : tmp28832;
  assign tmp31214 = s2 ? tmp31215 : tmp31217;
  assign tmp31220 = s1 ? tmp30184 : tmp31016;
  assign tmp31223 = l1 ? tmp27624 : tmp28661;
  assign tmp31222 = s0 ? tmp31223 : tmp30913;
  assign tmp31221 = s1 ? tmp30912 : tmp31222;
  assign tmp31219 = s2 ? tmp31220 : tmp31221;
  assign tmp31213 = s3 ? tmp31214 : tmp31219;
  assign tmp31204 = s4 ? tmp31205 : tmp31213;
  assign tmp31229 = s0 ? tmp31105 : 1;
  assign tmp31231 = l1 ? tmp27623 : tmp27560;
  assign tmp31230 = s0 ? 1 : tmp31231;
  assign tmp31228 = s1 ? tmp31229 : tmp31230;
  assign tmp31234 = l1 ? tmp27614 : tmp28779;
  assign tmp31233 = s0 ? 1 : tmp31234;
  assign tmp31232 = s1 ? tmp31233 : tmp30930;
  assign tmp31227 = s2 ? tmp31228 : tmp31232;
  assign tmp31239 = ~(l2 ? tmp27488 : tmp27490);
  assign tmp31238 = ~(l1 ? tmp27496 : tmp31239);
  assign tmp31237 = s0 ? 1 : tmp31238;
  assign tmp31241 = l1 ? tmp27624 : tmp28678;
  assign tmp31240 = s0 ? 1 : tmp31241;
  assign tmp31236 = s1 ? tmp31237 : tmp31240;
  assign tmp31243 = s0 ? tmp31223 : tmp28248;
  assign tmp31242 = s1 ? tmp31243 : tmp30939;
  assign tmp31235 = s2 ? tmp31236 : tmp31242;
  assign tmp31226 = s3 ? tmp31227 : tmp31235;
  assign tmp31248 = l1 ? tmp30899 : tmp28779;
  assign tmp31247 = s0 ? tmp31050 : tmp31248;
  assign tmp31246 = s1 ? tmp31247 : tmp30207;
  assign tmp31251 = l1 ? tmp27623 : tmp28779;
  assign tmp31250 = s0 ? tmp31251 : 1;
  assign tmp31249 = s1 ? tmp30207 : tmp31250;
  assign tmp31245 = s2 ? tmp31246 : tmp31249;
  assign tmp31256 = ~(l2 ? tmp27488 : tmp27492);
  assign tmp31255 = l1 ? tmp27504 : tmp31256;
  assign tmp31257 = ~(l1 ? tmp30915 : tmp28779);
  assign tmp31254 = s0 ? tmp31255 : tmp31257;
  assign tmp31258 = ~(s0 ? tmp28812 : tmp31040);
  assign tmp31253 = s1 ? tmp31254 : tmp31258;
  assign tmp31252 = ~(s2 ? tmp31253 : tmp31060);
  assign tmp31244 = s3 ? tmp31245 : tmp31252;
  assign tmp31225 = s4 ? tmp31226 : tmp31244;
  assign tmp31263 = s0 ? tmp31241 : tmp27504;
  assign tmp31264 = s0 ? tmp27504 : tmp28589;
  assign tmp31262 = s1 ? tmp31263 : tmp31264;
  assign tmp31266 = s0 ? tmp28540 : tmp27832;
  assign tmp31267 = s0 ? tmp27836 : tmp27832;
  assign tmp31265 = ~(s1 ? tmp31266 : tmp31267);
  assign tmp31261 = s2 ? tmp31262 : tmp31265;
  assign tmp31260 = s3 ? tmp31261 : tmp31071;
  assign tmp31272 = ~(l1 ? tmp27624 : tmp28661);
  assign tmp31271 = s0 ? tmp27560 : tmp31272;
  assign tmp31270 = s1 ? tmp31081 : tmp31271;
  assign tmp31275 = ~(l1 ? tmp27560 : tmp31256);
  assign tmp31274 = s0 ? tmp27504 : tmp31275;
  assign tmp31276 = ~(s0 ? tmp27832 : tmp27836);
  assign tmp31273 = ~(s1 ? tmp31274 : tmp31276);
  assign tmp31269 = s2 ? tmp31270 : tmp31273;
  assign tmp31279 = s0 ? tmp28540 : tmp28275;
  assign tmp31278 = s1 ? tmp31279 : tmp31092;
  assign tmp31277 = s2 ? tmp31278 : tmp31094;
  assign tmp31268 = ~(s3 ? tmp31269 : tmp31277);
  assign tmp31259 = s4 ? tmp31260 : tmp31268;
  assign tmp31224 = s5 ? tmp31225 : tmp31259;
  assign tmp31203 = s6 ? tmp31204 : tmp31224;
  assign tmp31202 = s7 ? tmp31203 : tmp27575;
  assign tmp31201 = s8 ? tmp31202 : tmp31203;
  assign tmp31200 = s9 ? tmp31201 : tmp27575;
  assign tmp30883 = s10 ? tmp30884 : tmp31200;
  assign tmp30562 = s12 ? tmp30563 : tmp30883;
  assign tmp31289 = l1 ? 1 : tmp28835;
  assign tmp31291 = l1 ? tmp31183 : tmp28835;
  assign tmp31290 = s0 ? 1 : tmp31291;
  assign tmp31288 = s1 ? tmp31289 : tmp31290;
  assign tmp31293 = s1 ? 1 : tmp31291;
  assign tmp31292 = s2 ? tmp31290 : tmp31293;
  assign tmp31287 = s3 ? tmp31288 : tmp31292;
  assign tmp31297 = s0 ? tmp31289 : 1;
  assign tmp31296 = s1 ? tmp31297 : tmp31291;
  assign tmp31298 = s1 ? tmp31297 : 1;
  assign tmp31295 = s2 ? tmp31296 : tmp31298;
  assign tmp31302 = l1 ? tmp28643 : tmp27504;
  assign tmp31301 = s0 ? 1 : tmp31302;
  assign tmp31300 = s1 ? 1 : tmp31301;
  assign tmp31304 = s0 ? tmp29713 : tmp31291;
  assign tmp31303 = s1 ? tmp31291 : tmp31304;
  assign tmp31299 = s2 ? tmp31300 : tmp31303;
  assign tmp31294 = s3 ? tmp31295 : tmp31299;
  assign tmp31286 = s4 ? tmp31287 : tmp31294;
  assign tmp31310 = s0 ? tmp31291 : 1;
  assign tmp31309 = s1 ? tmp31310 : 1;
  assign tmp31311 = s1 ? tmp31290 : tmp31310;
  assign tmp31308 = s2 ? tmp31309 : tmp31311;
  assign tmp31315 = l1 ? tmp31183 : tmp27760;
  assign tmp31314 = s0 ? 1 : tmp31315;
  assign tmp31313 = s1 ? 1 : tmp31314;
  assign tmp31317 = s0 ? tmp29713 : tmp31302;
  assign tmp31316 = s1 ? tmp31317 : tmp31315;
  assign tmp31312 = s2 ? tmp31313 : tmp31316;
  assign tmp31307 = s3 ? tmp31308 : tmp31312;
  assign tmp31321 = s0 ? tmp27636 : tmp31315;
  assign tmp31320 = s1 ? tmp31321 : 1;
  assign tmp31322 = s1 ? 1 : tmp31297;
  assign tmp31319 = s2 ? tmp31320 : tmp31322;
  assign tmp31325 = s0 ? tmp31289 : tmp27762;
  assign tmp31324 = s1 ? tmp31325 : tmp31314;
  assign tmp31327 = s0 ? tmp31302 : tmp27504;
  assign tmp31326 = s1 ? tmp27504 : tmp31327;
  assign tmp31323 = s2 ? tmp31324 : tmp31326;
  assign tmp31318 = s3 ? tmp31319 : tmp31323;
  assign tmp31306 = s4 ? tmp31307 : tmp31318;
  assign tmp31332 = s0 ? tmp31315 : 1;
  assign tmp31331 = s1 ? tmp31332 : 1;
  assign tmp31330 = s2 ? tmp31331 : 1;
  assign tmp31335 = s0 ? 1 : tmp27575;
  assign tmp31337 = ~(l1 ? tmp28643 : tmp27504);
  assign tmp31336 = ~(s0 ? tmp27495 : tmp31337);
  assign tmp31334 = s1 ? tmp31335 : tmp31336;
  assign tmp31339 = s0 ? tmp31302 : tmp27636;
  assign tmp31340 = s0 ? tmp27636 : tmp28835;
  assign tmp31338 = s1 ? tmp31339 : tmp31340;
  assign tmp31333 = s2 ? tmp31334 : tmp31338;
  assign tmp31329 = s3 ? tmp31330 : tmp31333;
  assign tmp31345 = l1 ? tmp27560 : tmp27575;
  assign tmp31344 = s0 ? tmp28835 : tmp31345;
  assign tmp31346 = s0 ? tmp31345 : tmp29713;
  assign tmp31343 = s1 ? tmp31344 : tmp31346;
  assign tmp31347 = s1 ? tmp31290 : 1;
  assign tmp31342 = s2 ? tmp31343 : tmp31347;
  assign tmp31350 = s0 ? 1 : tmp29713;
  assign tmp31351 = s0 ? tmp31302 : tmp31315;
  assign tmp31349 = s1 ? tmp31350 : tmp31351;
  assign tmp31354 = ~(l1 ? tmp27560 : tmp27575);
  assign tmp31353 = ~(s0 ? tmp27495 : tmp31354);
  assign tmp31352 = s1 ? tmp31340 : tmp31353;
  assign tmp31348 = s2 ? tmp31349 : tmp31352;
  assign tmp31341 = s3 ? tmp31342 : tmp31348;
  assign tmp31328 = s4 ? tmp31329 : tmp31341;
  assign tmp31305 = s5 ? tmp31306 : tmp31328;
  assign tmp31285 = s6 ? tmp31286 : tmp31305;
  assign tmp31284 = s7 ? tmp31285 : tmp27575;
  assign tmp31361 = s0 ? 1 : tmp29736;
  assign tmp31360 = s1 ? 1 : tmp31361;
  assign tmp31359 = s2 ? tmp31360 : tmp31303;
  assign tmp31358 = s3 ? tmp31295 : tmp31359;
  assign tmp31357 = s4 ? tmp31287 : tmp31358;
  assign tmp31367 = s0 ? tmp29713 : tmp29736;
  assign tmp31366 = s1 ? tmp31367 : tmp31315;
  assign tmp31365 = s2 ? tmp31313 : tmp31366;
  assign tmp31364 = s3 ? tmp31308 : tmp31365;
  assign tmp31371 = s0 ? tmp29736 : tmp27504;
  assign tmp31370 = s1 ? tmp27504 : tmp31371;
  assign tmp31369 = s2 ? tmp31324 : tmp31370;
  assign tmp31368 = s3 ? tmp31319 : tmp31369;
  assign tmp31363 = s4 ? tmp31364 : tmp31368;
  assign tmp31376 = ~(s0 ? 1 : tmp29733);
  assign tmp31375 = s1 ? tmp27999 : tmp31376;
  assign tmp31378 = s0 ? tmp29736 : tmp27636;
  assign tmp31377 = s1 ? tmp31378 : tmp31340;
  assign tmp31374 = s2 ? tmp31375 : tmp31377;
  assign tmp31373 = s3 ? tmp31330 : tmp31374;
  assign tmp31382 = s0 ? tmp28835 : tmp28275;
  assign tmp31383 = s0 ? tmp28275 : tmp29713;
  assign tmp31381 = s1 ? tmp31382 : tmp31383;
  assign tmp31380 = s2 ? tmp31381 : tmp31347;
  assign tmp31386 = s0 ? tmp29736 : tmp31315;
  assign tmp31385 = s1 ? tmp31350 : tmp31386;
  assign tmp31389 = ~(l1 ? tmp27560 : 0);
  assign tmp31388 = ~(s0 ? 1 : tmp31389);
  assign tmp31387 = s1 ? tmp31340 : tmp31388;
  assign tmp31384 = s2 ? tmp31385 : tmp31387;
  assign tmp31379 = s3 ? tmp31380 : tmp31384;
  assign tmp31372 = s4 ? tmp31373 : tmp31379;
  assign tmp31362 = s5 ? tmp31363 : tmp31372;
  assign tmp31356 = s6 ? tmp31357 : tmp31362;
  assign tmp31355 = s7 ? tmp31356 : tmp27575;
  assign tmp31283 = s8 ? tmp31284 : tmp31355;
  assign tmp31397 = l2 ? 1 : tmp27509;
  assign tmp31396 = l1 ? 1 : tmp31397;
  assign tmp31399 = l1 ? tmp31183 : tmp27560;
  assign tmp31398 = s0 ? tmp27750 : tmp31399;
  assign tmp31395 = s1 ? tmp31396 : tmp31398;
  assign tmp31402 = l1 ? tmp31183 : tmp31397;
  assign tmp31401 = s0 ? tmp27750 : tmp31402;
  assign tmp31403 = s1 ? tmp27750 : tmp31402;
  assign tmp31400 = s2 ? tmp31401 : tmp31403;
  assign tmp31394 = s3 ? tmp31395 : tmp31400;
  assign tmp31408 = l1 ? 1 : tmp27560;
  assign tmp31407 = s0 ? tmp31408 : tmp27750;
  assign tmp31406 = s1 ? tmp31407 : tmp31402;
  assign tmp31410 = s0 ? tmp31396 : tmp27750;
  assign tmp31409 = s1 ? tmp31410 : tmp27750;
  assign tmp31405 = s2 ? tmp31406 : tmp31409;
  assign tmp31413 = s0 ? tmp27750 : tmp29736;
  assign tmp31412 = s1 ? tmp27750 : tmp31413;
  assign tmp31415 = s0 ? tmp29713 : tmp31402;
  assign tmp31414 = s1 ? tmp31402 : tmp31415;
  assign tmp31411 = s2 ? tmp31412 : tmp31414;
  assign tmp31404 = s3 ? tmp31405 : tmp31411;
  assign tmp31393 = s4 ? tmp31394 : tmp31404;
  assign tmp31421 = s0 ? tmp31399 : tmp27750;
  assign tmp31420 = s1 ? tmp31421 : tmp27750;
  assign tmp31424 = l1 ? tmp31183 : tmp27504;
  assign tmp31423 = s0 ? tmp27750 : tmp31424;
  assign tmp31425 = s0 ? tmp31402 : tmp27750;
  assign tmp31422 = s1 ? tmp31423 : tmp31425;
  assign tmp31419 = s2 ? tmp31420 : tmp31422;
  assign tmp31427 = s1 ? tmp27750 : tmp31423;
  assign tmp31428 = s1 ? tmp31367 : tmp31424;
  assign tmp31426 = s2 ? tmp31427 : tmp31428;
  assign tmp31418 = s3 ? tmp31419 : tmp31426;
  assign tmp31432 = s0 ? tmp27636 : tmp31424;
  assign tmp31431 = s1 ? tmp31432 : tmp27750;
  assign tmp31433 = s1 ? tmp27750 : tmp28365;
  assign tmp31430 = s2 ? tmp31431 : tmp31433;
  assign tmp31435 = s1 ? tmp27636 : tmp31423;
  assign tmp31434 = s2 ? tmp31435 : tmp31370;
  assign tmp31429 = s3 ? tmp31430 : tmp31434;
  assign tmp31417 = s4 ? tmp31418 : tmp31429;
  assign tmp31440 = s0 ? tmp31424 : tmp27750;
  assign tmp31439 = s1 ? tmp31440 : tmp27750;
  assign tmp31438 = s2 ? tmp31439 : tmp27750;
  assign tmp31443 = s0 ? tmp27750 : 0;
  assign tmp31442 = s1 ? tmp31443 : tmp31376;
  assign tmp31444 = s1 ? tmp31378 : tmp27636;
  assign tmp31441 = s2 ? tmp31442 : tmp31444;
  assign tmp31437 = s3 ? tmp31438 : tmp31441;
  assign tmp31448 = s0 ? tmp27636 : tmp28275;
  assign tmp31447 = s1 ? tmp31448 : tmp31383;
  assign tmp31449 = s1 ? tmp31423 : tmp27750;
  assign tmp31446 = s2 ? tmp31447 : tmp31449;
  assign tmp31452 = s0 ? tmp27750 : tmp29713;
  assign tmp31453 = s0 ? tmp29736 : tmp31424;
  assign tmp31451 = s1 ? tmp31452 : tmp31453;
  assign tmp31454 = s1 ? tmp27636 : tmp31388;
  assign tmp31450 = s2 ? tmp31451 : tmp31454;
  assign tmp31445 = s3 ? tmp31446 : tmp31450;
  assign tmp31436 = s4 ? tmp31437 : tmp31445;
  assign tmp31416 = s5 ? tmp31417 : tmp31436;
  assign tmp31392 = s6 ? tmp31393 : tmp31416;
  assign tmp31391 = s7 ? tmp31392 : tmp27575;
  assign tmp31390 = s8 ? tmp31355 : tmp31391;
  assign tmp31282 = s9 ? tmp31283 : tmp31390;
  assign tmp31456 = s8 ? tmp31355 : tmp31356;
  assign tmp31455 = s9 ? tmp31456 : tmp27575;
  assign tmp31281 = s10 ? tmp31282 : tmp31455;
  assign tmp31465 = l1 ? tmp30069 : tmp27560;
  assign tmp31466 = ~(l1 ? tmp29442 : tmp28495);
  assign tmp31464 = s1 ? tmp31465 : tmp31466;
  assign tmp31470 = ~(l1 ? tmp30069 : tmp27560);
  assign tmp31469 = s0 ? tmp30650 : tmp31470;
  assign tmp31472 = l1 ? tmp29442 : tmp28495;
  assign tmp31471 = s0 ? tmp31472 : tmp31470;
  assign tmp31468 = s1 ? tmp31469 : tmp31471;
  assign tmp31474 = s0 ? tmp31472 : 0;
  assign tmp31473 = s1 ? tmp31474 : tmp31470;
  assign tmp31467 = ~(s2 ? tmp31468 : tmp31473);
  assign tmp31463 = s3 ? tmp31464 : tmp31467;
  assign tmp31479 = l1 ? tmp27517 : tmp28495;
  assign tmp31478 = s0 ? tmp31479 : 0;
  assign tmp31477 = s1 ? tmp31478 : tmp31470;
  assign tmp31481 = s0 ? tmp31465 : 1;
  assign tmp31480 = ~(s1 ? tmp31481 : 1);
  assign tmp31476 = s2 ? tmp31477 : tmp31480;
  assign tmp31485 = l1 ? tmp27504 : tmp27560;
  assign tmp31484 = s0 ? 1 : tmp31485;
  assign tmp31483 = s1 ? 1 : tmp31484;
  assign tmp31489 = l2 ? tmp27554 : tmp27491;
  assign tmp31488 = l1 ? tmp31489 : tmp27560;
  assign tmp31487 = s0 ? tmp31465 : tmp31488;
  assign tmp31492 = l2 ? tmp27554 : 0;
  assign tmp31491 = l1 ? tmp31492 : tmp27560;
  assign tmp31490 = s0 ? tmp31491 : tmp31465;
  assign tmp31486 = s1 ? tmp31487 : tmp31490;
  assign tmp31482 = ~(s2 ? tmp31483 : tmp31486);
  assign tmp31475 = ~(s3 ? tmp31476 : tmp31482);
  assign tmp31462 = s4 ? tmp31463 : tmp31475;
  assign tmp31497 = s1 ? tmp31474 : tmp30925;
  assign tmp31500 = ~(l1 ? tmp29442 : tmp27833);
  assign tmp31499 = s0 ? 1 : tmp31500;
  assign tmp31501 = s0 ? tmp31488 : 1;
  assign tmp31498 = ~(s1 ? tmp31499 : tmp31501);
  assign tmp31496 = s2 ? tmp31497 : tmp31498;
  assign tmp31505 = ~(l1 ? tmp29414 : tmp28495);
  assign tmp31504 = s0 ? 1 : tmp31505;
  assign tmp31506 = s0 ? 1 : tmp31488;
  assign tmp31503 = s1 ? tmp31504 : tmp31506;
  assign tmp31508 = s0 ? tmp31491 : tmp27836;
  assign tmp31507 = s1 ? tmp31508 : tmp31487;
  assign tmp31502 = ~(s2 ? tmp31503 : tmp31507);
  assign tmp31495 = s3 ? tmp31496 : tmp31502;
  assign tmp31512 = s0 ? tmp31485 : tmp31465;
  assign tmp31511 = s1 ? tmp31512 : 1;
  assign tmp31514 = ~(s0 ? tmp30964 : 0);
  assign tmp31513 = s1 ? 1 : tmp31514;
  assign tmp31510 = s2 ? tmp31511 : tmp31513;
  assign tmp31518 = ~(l1 ? tmp30915 : tmp27560);
  assign tmp31517 = s0 ? tmp30964 : tmp31518;
  assign tmp31519 = ~(s0 ? 1 : tmp31488);
  assign tmp31516 = s1 ? tmp31517 : tmp31519;
  assign tmp31521 = s0 ? tmp31485 : 1;
  assign tmp31520 = ~(s1 ? 1 : tmp31521);
  assign tmp31515 = ~(s2 ? tmp31516 : tmp31520);
  assign tmp31509 = ~(s3 ? tmp31510 : tmp31515);
  assign tmp31494 = s4 ? tmp31495 : tmp31509;
  assign tmp31526 = s0 ? tmp31488 : tmp27504;
  assign tmp31527 = s0 ? tmp27504 : tmp27530;
  assign tmp31525 = s1 ? tmp31526 : tmp31527;
  assign tmp31529 = s0 ? tmp27533 : tmp30964;
  assign tmp31528 = ~(s1 ? tmp31529 : tmp30965);
  assign tmp31524 = s2 ? tmp31525 : tmp31528;
  assign tmp31533 = l1 ? tmp27495 : tmp28490;
  assign tmp31532 = s0 ? tmp29880 : tmp31533;
  assign tmp31534 = s0 ? tmp31533 : tmp27533;
  assign tmp31531 = s1 ? tmp31532 : tmp31534;
  assign tmp31537 = ~(l1 ? tmp27504 : tmp27560);
  assign tmp31536 = s0 ? tmp27533 : tmp31537;
  assign tmp31539 = ~(l1 ? tmp27517 : tmp27833);
  assign tmp31538 = ~(s0 ? tmp31485 : tmp31539);
  assign tmp31535 = s1 ? tmp31536 : tmp31538;
  assign tmp31530 = ~(s2 ? tmp31531 : tmp31535);
  assign tmp31523 = s3 ? tmp31524 : tmp31530;
  assign tmp31543 = s0 ? tmp30964 : tmp27495;
  assign tmp31545 = ~(l1 ? tmp31492 : tmp27560);
  assign tmp31544 = s0 ? tmp27495 : tmp31545;
  assign tmp31542 = s1 ? tmp31543 : tmp31544;
  assign tmp31548 = ~(l1 ? tmp27496 : tmp27833);
  assign tmp31547 = s0 ? tmp27504 : tmp31548;
  assign tmp31546 = ~(s1 ? tmp31547 : tmp30984);
  assign tmp31541 = s2 ? tmp31542 : tmp31546;
  assign tmp31551 = s0 ? tmp27533 : tmp31533;
  assign tmp31553 = ~(l1 ? tmp31489 : tmp27560);
  assign tmp31552 = s0 ? tmp27533 : tmp31553;
  assign tmp31550 = s1 ? tmp31551 : tmp31552;
  assign tmp31555 = s0 ? tmp31485 : tmp31539;
  assign tmp31556 = ~(s0 ? tmp31533 : tmp27495);
  assign tmp31554 = ~(s1 ? tmp31555 : tmp31556);
  assign tmp31549 = s2 ? tmp31550 : tmp31554;
  assign tmp31540 = ~(s3 ? tmp31541 : tmp31549);
  assign tmp31522 = ~(s4 ? tmp31523 : tmp31540);
  assign tmp31493 = ~(s5 ? tmp31494 : tmp31522);
  assign tmp31461 = s6 ? tmp31462 : tmp31493;
  assign tmp31460 = s7 ? tmp31461 : tmp27575;
  assign tmp31562 = l1 ? tmp30069 : tmp29414;
  assign tmp31563 = l1 ? tmp27488 : tmp29414;
  assign tmp31561 = s1 ? tmp31562 : tmp31563;
  assign tmp31566 = s0 ? tmp31030 : tmp31562;
  assign tmp31567 = s0 ? tmp31563 : tmp31562;
  assign tmp31565 = s1 ? tmp31566 : tmp31567;
  assign tmp31569 = s0 ? tmp31563 : tmp27642;
  assign tmp31568 = s1 ? tmp31569 : tmp31562;
  assign tmp31564 = s2 ? tmp31565 : tmp31568;
  assign tmp31560 = s3 ? tmp31561 : tmp31564;
  assign tmp31574 = l1 ? tmp27623 : tmp29414;
  assign tmp31573 = s0 ? tmp31574 : 1;
  assign tmp31572 = s1 ? tmp31573 : tmp31562;
  assign tmp31576 = s0 ? tmp31562 : 1;
  assign tmp31578 = l1 ? 1 : tmp27496;
  assign tmp31577 = s0 ? tmp31578 : 1;
  assign tmp31575 = s1 ? tmp31576 : tmp31577;
  assign tmp31571 = s2 ? tmp31572 : tmp31575;
  assign tmp31582 = l1 ? 1 : tmp27495;
  assign tmp31581 = s0 ? tmp31578 : tmp31582;
  assign tmp31580 = s1 ? tmp31581 : tmp31484;
  assign tmp31585 = l1 ? tmp31489 : tmp29414;
  assign tmp31584 = s0 ? tmp31562 : tmp31585;
  assign tmp31588 = ~(l2 ? tmp27488 : tmp27506);
  assign tmp31587 = l1 ? tmp27497 : tmp31588;
  assign tmp31586 = s0 ? tmp31587 : tmp31562;
  assign tmp31583 = s1 ? tmp31584 : tmp31586;
  assign tmp31579 = s2 ? tmp31580 : tmp31583;
  assign tmp31570 = s3 ? tmp31571 : tmp31579;
  assign tmp31559 = s4 ? tmp31560 : tmp31570;
  assign tmp31594 = s0 ? tmp31563 : 1;
  assign tmp31593 = s1 ? tmp31594 : tmp31029;
  assign tmp31597 = l1 ? tmp27488 : tmp27517;
  assign tmp31596 = s0 ? 1 : tmp31597;
  assign tmp31598 = s0 ? tmp31585 : tmp27642;
  assign tmp31595 = s1 ? tmp31596 : tmp31598;
  assign tmp31592 = s2 ? tmp31593 : tmp31595;
  assign tmp31602 = ~(l1 ? tmp27496 : tmp27898);
  assign tmp31601 = s0 ? tmp27642 : tmp31602;
  assign tmp31604 = l1 ? tmp27521 : tmp29414;
  assign tmp31603 = s0 ? tmp27642 : tmp31604;
  assign tmp31600 = s1 ? tmp31601 : tmp31603;
  assign tmp31606 = s0 ? tmp31587 : tmp27836;
  assign tmp31608 = l1 ? tmp31489 : tmp31588;
  assign tmp31607 = s0 ? tmp31562 : tmp31608;
  assign tmp31605 = s1 ? tmp31606 : tmp31607;
  assign tmp31599 = s2 ? tmp31600 : tmp31605;
  assign tmp31591 = s3 ? tmp31592 : tmp31599;
  assign tmp31612 = s0 ? tmp31485 : tmp31562;
  assign tmp31613 = s0 ? 1 : tmp28540;
  assign tmp31611 = s1 ? tmp31612 : tmp31613;
  assign tmp31616 = l1 ? tmp27623 : tmp27517;
  assign tmp31615 = s0 ? tmp31616 : 1;
  assign tmp31614 = s1 ? tmp31613 : tmp31615;
  assign tmp31610 = s2 ? tmp31611 : tmp31614;
  assign tmp31620 = ~(l1 ? tmp30915 : tmp31588);
  assign tmp31619 = s0 ? tmp30972 : tmp31620;
  assign tmp31622 = l1 ? tmp27521 : tmp27560;
  assign tmp31621 = ~(s0 ? tmp28540 : tmp31622);
  assign tmp31618 = s1 ? tmp31619 : tmp31621;
  assign tmp31617 = ~(s2 ? tmp31618 : tmp31520);
  assign tmp31609 = s3 ? tmp31610 : tmp31617;
  assign tmp31590 = s4 ? tmp31591 : tmp31609;
  assign tmp31627 = s0 ? tmp31604 : tmp27504;
  assign tmp31628 = s0 ? tmp27504 : tmp29123;
  assign tmp31626 = s1 ? tmp31627 : tmp31628;
  assign tmp31630 = s0 ? tmp28812 : tmp27819;
  assign tmp31629 = ~(s1 ? tmp31630 : tmp31070);
  assign tmp31625 = s2 ? tmp31626 : tmp31629;
  assign tmp31633 = s0 ? tmp27836 : tmp28033;
  assign tmp31634 = s0 ? tmp28033 : tmp27640;
  assign tmp31632 = s1 ? tmp31633 : tmp31634;
  assign tmp31636 = s0 ? tmp27640 : tmp31537;
  assign tmp31637 = ~(s0 ? tmp31485 : tmp31075);
  assign tmp31635 = s1 ? tmp31636 : tmp31637;
  assign tmp31631 = ~(s2 ? tmp31632 : tmp31635);
  assign tmp31624 = s3 ? tmp31625 : tmp31631;
  assign tmp31641 = s0 ? tmp27832 : 1;
  assign tmp31643 = ~(l1 ? tmp27497 : tmp31588);
  assign tmp31642 = s0 ? 1 : tmp31643;
  assign tmp31640 = s1 ? tmp31641 : tmp31642;
  assign tmp31646 = ~(l1 ? tmp27744 : tmp27960);
  assign tmp31645 = s0 ? tmp27504 : tmp31646;
  assign tmp31644 = ~(s1 ? tmp31645 : tmp31088);
  assign tmp31639 = s2 ? tmp31640 : tmp31644;
  assign tmp31649 = s0 ? tmp28812 : tmp28033;
  assign tmp31651 = ~(l1 ? tmp27521 : tmp27560);
  assign tmp31650 = s0 ? tmp27640 : tmp31651;
  assign tmp31648 = s1 ? tmp31649 : tmp31650;
  assign tmp31653 = s0 ? tmp31485 : tmp31075;
  assign tmp31654 = ~(s0 ? tmp28033 : 1);
  assign tmp31652 = ~(s1 ? tmp31653 : tmp31654);
  assign tmp31647 = s2 ? tmp31648 : tmp31652;
  assign tmp31638 = ~(s3 ? tmp31639 : tmp31647);
  assign tmp31623 = s4 ? tmp31624 : tmp31638;
  assign tmp31589 = s5 ? tmp31590 : tmp31623;
  assign tmp31558 = s6 ? tmp31559 : tmp31589;
  assign tmp31557 = s7 ? tmp31558 : tmp27575;
  assign tmp31459 = s8 ? tmp31460 : tmp31557;
  assign tmp31661 = l1 ? tmp27488 : tmp27560;
  assign tmp31660 = s1 ? tmp31465 : tmp31661;
  assign tmp31664 = s0 ? tmp31135 : tmp31465;
  assign tmp31666 = l1 ? tmp27488 : tmp27744;
  assign tmp31665 = s0 ? tmp31666 : tmp31465;
  assign tmp31663 = s1 ? tmp31664 : tmp31665;
  assign tmp31668 = s0 ? tmp31666 : tmp27750;
  assign tmp31667 = s1 ? tmp31668 : tmp31465;
  assign tmp31662 = s2 ? tmp31663 : tmp31667;
  assign tmp31659 = s3 ? tmp31660 : tmp31662;
  assign tmp31672 = s0 ? tmp31231 : tmp27750;
  assign tmp31671 = s1 ? tmp31672 : tmp31465;
  assign tmp31674 = s0 ? tmp31465 : tmp27750;
  assign tmp31673 = s1 ? tmp31674 : tmp27750;
  assign tmp31670 = s2 ? tmp31671 : tmp31673;
  assign tmp31677 = s0 ? tmp27750 : tmp31485;
  assign tmp31676 = s1 ? tmp27750 : tmp31677;
  assign tmp31680 = l1 ? tmp27497 : tmp27560;
  assign tmp31679 = s0 ? tmp31680 : tmp31465;
  assign tmp31678 = s1 ? tmp31487 : tmp31679;
  assign tmp31675 = s2 ? tmp31676 : tmp31678;
  assign tmp31669 = s3 ? tmp31670 : tmp31675;
  assign tmp31658 = s4 ? tmp31659 : tmp31669;
  assign tmp31686 = s0 ? tmp31661 : tmp27750;
  assign tmp31685 = s1 ? tmp31686 : tmp31134;
  assign tmp31689 = l1 ? tmp27488 : tmp27504;
  assign tmp31688 = s0 ? tmp27750 : tmp31689;
  assign tmp31690 = s0 ? tmp31488 : tmp27750;
  assign tmp31687 = s1 ? tmp31688 : tmp31690;
  assign tmp31684 = s2 ? tmp31685 : tmp31687;
  assign tmp31694 = ~(l1 ? tmp27496 : tmp27809);
  assign tmp31693 = s0 ? tmp27750 : tmp31694;
  assign tmp31695 = s0 ? tmp27750 : tmp31622;
  assign tmp31692 = s1 ? tmp31693 : tmp31695;
  assign tmp31697 = s0 ? tmp31680 : tmp27743;
  assign tmp31696 = s1 ? tmp31697 : tmp31487;
  assign tmp31691 = s2 ? tmp31692 : tmp31696;
  assign tmp31683 = s3 ? tmp31684 : tmp31691;
  assign tmp31700 = s1 ? tmp31512 : tmp27750;
  assign tmp31703 = l1 ? tmp27623 : tmp27504;
  assign tmp31702 = s0 ? tmp31703 : tmp27750;
  assign tmp31701 = s1 ? tmp27750 : tmp31702;
  assign tmp31699 = s2 ? tmp31700 : tmp31701;
  assign tmp31706 = s0 ? tmp27832 : tmp31518;
  assign tmp31707 = ~(s0 ? tmp27750 : tmp31622);
  assign tmp31705 = s1 ? tmp31706 : tmp31707;
  assign tmp31709 = s0 ? tmp31485 : tmp27750;
  assign tmp31708 = ~(s1 ? tmp27750 : tmp31709);
  assign tmp31704 = ~(s2 ? tmp31705 : tmp31708);
  assign tmp31698 = s3 ? tmp31699 : tmp31704;
  assign tmp31682 = s4 ? tmp31683 : tmp31698;
  assign tmp31714 = s0 ? tmp31622 : tmp27504;
  assign tmp31715 = s0 ? tmp27504 : tmp29225;
  assign tmp31713 = s1 ? tmp31714 : tmp31715;
  assign tmp31716 = ~(s1 ? tmp29229 : tmp31170);
  assign tmp31712 = s2 ? tmp31713 : tmp31716;
  assign tmp31719 = s0 ? tmp29180 : tmp28033;
  assign tmp31720 = s0 ? tmp28033 : tmp29230;
  assign tmp31718 = s1 ? tmp31719 : tmp31720;
  assign tmp31722 = s0 ? tmp29230 : tmp31537;
  assign tmp31721 = s1 ? tmp31722 : tmp31637;
  assign tmp31717 = ~(s2 ? tmp31718 : tmp31721);
  assign tmp31711 = s3 ? tmp31712 : tmp31717;
  assign tmp31727 = ~(l1 ? tmp27497 : tmp27560);
  assign tmp31726 = s0 ? 1 : tmp31727;
  assign tmp31725 = s1 ? tmp31641 : tmp31726;
  assign tmp31730 = ~(l1 ? tmp27744 : tmp27833);
  assign tmp31729 = s0 ? tmp27504 : tmp31730;
  assign tmp31728 = ~(s1 ? tmp31729 : tmp31189);
  assign tmp31724 = s2 ? tmp31725 : tmp31728;
  assign tmp31733 = s0 ? tmp29230 : tmp28033;
  assign tmp31734 = s0 ? tmp29230 : tmp31651;
  assign tmp31732 = s1 ? tmp31733 : tmp31734;
  assign tmp31731 = s2 ? tmp31732 : tmp31652;
  assign tmp31723 = ~(s3 ? tmp31724 : tmp31731);
  assign tmp31710 = s4 ? tmp31711 : tmp31723;
  assign tmp31681 = s5 ? tmp31682 : tmp31710;
  assign tmp31657 = s6 ? tmp31658 : tmp31681;
  assign tmp31656 = s7 ? tmp31657 : tmp27575;
  assign tmp31655 = s8 ? tmp31557 : tmp31656;
  assign tmp31458 = s9 ? tmp31459 : tmp31655;
  assign tmp31743 = s0 ? tmp31231 : tmp31465;
  assign tmp31744 = s0 ? tmp31661 : tmp31465;
  assign tmp31742 = s1 ? tmp31743 : tmp31744;
  assign tmp31746 = s0 ? tmp31661 : 1;
  assign tmp31745 = s1 ? tmp31746 : tmp31465;
  assign tmp31741 = s2 ? tmp31742 : tmp31745;
  assign tmp31740 = s3 ? tmp31660 : tmp31741;
  assign tmp31750 = s0 ? tmp31231 : 1;
  assign tmp31749 = s1 ? tmp31750 : tmp31465;
  assign tmp31751 = s1 ? tmp31481 : 1;
  assign tmp31748 = s2 ? tmp31749 : tmp31751;
  assign tmp31752 = s2 ? tmp31483 : tmp31678;
  assign tmp31747 = s3 ? tmp31748 : tmp31752;
  assign tmp31739 = s4 ? tmp31740 : tmp31747;
  assign tmp31757 = s1 ? tmp31746 : tmp31230;
  assign tmp31759 = s0 ? 1 : tmp31689;
  assign tmp31758 = s1 ? tmp31759 : tmp31501;
  assign tmp31756 = s2 ? tmp31757 : tmp31758;
  assign tmp31763 = ~(l1 ? tmp27496 : tmp28495);
  assign tmp31762 = s0 ? 1 : tmp31763;
  assign tmp31764 = s0 ? 1 : tmp31622;
  assign tmp31761 = s1 ? tmp31762 : tmp31764;
  assign tmp31766 = s0 ? tmp31680 : tmp27836;
  assign tmp31765 = s1 ? tmp31766 : tmp31487;
  assign tmp31760 = s2 ? tmp31761 : tmp31765;
  assign tmp31755 = s3 ? tmp31756 : tmp31760;
  assign tmp31770 = s0 ? tmp31703 : 1;
  assign tmp31769 = s1 ? 1 : tmp31770;
  assign tmp31768 = s2 ? tmp31511 : tmp31769;
  assign tmp31773 = ~(s0 ? 1 : tmp31622);
  assign tmp31772 = s1 ? tmp31706 : tmp31773;
  assign tmp31771 = ~(s2 ? tmp31772 : tmp31520);
  assign tmp31767 = s3 ? tmp31768 : tmp31771;
  assign tmp31754 = s4 ? tmp31755 : tmp31767;
  assign tmp31778 = s0 ? tmp27504 : tmp29958;
  assign tmp31777 = s1 ? tmp31714 : tmp31778;
  assign tmp31780 = s0 ? tmp27640 : tmp27832;
  assign tmp31779 = ~(s1 ? tmp31780 : tmp31267);
  assign tmp31776 = s2 ? tmp31777 : tmp31779;
  assign tmp31775 = s3 ? tmp31776 : tmp31631;
  assign tmp31783 = ~(s1 ? tmp31729 : tmp31276);
  assign tmp31782 = s2 ? tmp31725 : tmp31783;
  assign tmp31786 = s0 ? tmp27640 : tmp28033;
  assign tmp31785 = s1 ? tmp31786 : tmp31650;
  assign tmp31784 = s2 ? tmp31785 : tmp31652;
  assign tmp31781 = ~(s3 ? tmp31782 : tmp31784);
  assign tmp31774 = s4 ? tmp31775 : tmp31781;
  assign tmp31753 = s5 ? tmp31754 : tmp31774;
  assign tmp31738 = s6 ? tmp31739 : tmp31753;
  assign tmp31737 = s7 ? tmp31738 : tmp27575;
  assign tmp31736 = s8 ? tmp31737 : tmp31738;
  assign tmp31735 = s9 ? tmp31736 : tmp27575;
  assign tmp31457 = s10 ? tmp31458 : tmp31735;
  assign tmp31280 = s12 ? tmp31281 : tmp31457;
  assign tmp30561 = ~(s13 ? tmp30562 : tmp31280);
  assign tmp29601 = ~(s14 ? tmp29602 : tmp30561);
  assign tmp27474 = s15 ? tmp27475 : tmp29601;
  assign tmp31798 = s0 ? tmp29204 : tmp27618;
  assign tmp31797 = s1 ? tmp27613 : tmp31798;
  assign tmp31801 = s0 ? tmp27627 : tmp29204;
  assign tmp31800 = s1 ? tmp31801 : tmp27630;
  assign tmp31799 = s2 ? tmp27620 : tmp31800;
  assign tmp31796 = s3 ? tmp31797 : tmp31799;
  assign tmp31805 = s0 ? tmp27635 : tmp27762;
  assign tmp31804 = s1 ? tmp31805 : tmp27637;
  assign tmp31807 = s0 ? tmp27613 : tmp29230;
  assign tmp31808 = s0 ? tmp29218 : tmp29230;
  assign tmp31806 = s1 ? tmp31807 : tmp31808;
  assign tmp31803 = s2 ? tmp31804 : tmp31806;
  assign tmp31811 = s0 ? tmp29218 : tmp29204;
  assign tmp31810 = s1 ? tmp31811 : tmp29825;
  assign tmp31813 = ~(s0 ? tmp27750 : tmp27649);
  assign tmp31812 = s1 ? tmp27625 : tmp31813;
  assign tmp31809 = s2 ? tmp31810 : tmp31812;
  assign tmp31802 = s3 ? tmp31803 : tmp31809;
  assign tmp31795 = s4 ? tmp31796 : tmp31802;
  assign tmp31819 = s0 ? tmp27618 : tmp27762;
  assign tmp31820 = s0 ? tmp27762 : tmp27622;
  assign tmp31818 = s1 ? tmp31819 : tmp31820;
  assign tmp31822 = s0 ? tmp27762 : tmp27659;
  assign tmp31823 = s0 ? tmp27625 : tmp29204;
  assign tmp31821 = s1 ? tmp31822 : tmp31823;
  assign tmp31817 = s2 ? tmp31818 : tmp31821;
  assign tmp31826 = s0 ? tmp29204 : tmp27664;
  assign tmp31827 = s0 ? tmp29204 : tmp27667;
  assign tmp31825 = s1 ? tmp31826 : tmp31827;
  assign tmp31828 = ~(s1 ? tmp27750 : tmp27669);
  assign tmp31824 = s2 ? tmp31825 : tmp31828;
  assign tmp31816 = s3 ? tmp31817 : tmp31824;
  assign tmp31832 = s0 ? tmp27750 : tmp27674;
  assign tmp31833 = ~(s0 ? 1 : tmp29230);
  assign tmp31831 = s1 ? tmp31832 : tmp31833;
  assign tmp31834 = ~(s1 ? tmp29532 : tmp27678);
  assign tmp31830 = s2 ? tmp31831 : tmp31834;
  assign tmp31837 = ~(s0 ? tmp29230 : tmp27488);
  assign tmp31836 = s1 ? tmp27682 : tmp31837;
  assign tmp31835 = s2 ? tmp31836 : tmp27750;
  assign tmp31829 = ~(s3 ? tmp31830 : tmp31835);
  assign tmp31815 = s4 ? tmp31816 : tmp31829;
  assign tmp31842 = s0 ? tmp27667 : tmp27791;
  assign tmp31841 = s1 ? tmp31842 : tmp27791;
  assign tmp31844 = s0 ? tmp27750 : tmp27694;
  assign tmp31843 = ~(s1 ? tmp31844 : tmp27696);
  assign tmp31840 = s2 ? tmp31841 : tmp31843;
  assign tmp31847 = s0 ? tmp27750 : tmp27703;
  assign tmp31846 = s1 ? tmp27750 : tmp31847;
  assign tmp31845 = ~(s2 ? tmp28901 : tmp31846);
  assign tmp31839 = s3 ? tmp31840 : tmp31845;
  assign tmp31851 = s0 ? tmp27703 : tmp27750;
  assign tmp31850 = s1 ? tmp31851 : tmp27750;
  assign tmp31853 = s0 ? tmp27750 : tmp27710;
  assign tmp31852 = s1 ? tmp31853 : tmp27711;
  assign tmp31849 = s2 ? tmp31850 : tmp31852;
  assign tmp31856 = s0 ? tmp27750 : tmp27715;
  assign tmp31855 = s1 ? tmp27750 : tmp31856;
  assign tmp31857 = s1 ? tmp31847 : tmp27750;
  assign tmp31854 = s2 ? tmp31855 : tmp31857;
  assign tmp31848 = ~(s3 ? tmp31849 : tmp31854);
  assign tmp31838 = s4 ? tmp31839 : tmp31848;
  assign tmp31814 = s5 ? tmp31815 : tmp31838;
  assign tmp31794 = s6 ? tmp31795 : tmp31814;
  assign tmp31793 = s7 ? tmp31794 : tmp27495;
  assign tmp31792 = ~(s8 ? tmp27718 : tmp31793);
  assign tmp31791 = s9 ? tmp27479 : tmp31792;
  assign tmp31859 = s8 ? tmp27718 : tmp27609;
  assign tmp31858 = ~(s9 ? tmp31859 : tmp27495);
  assign tmp31790 = s10 ? tmp31791 : tmp31858;
  assign tmp31869 = l1 ? tmp27971 : tmp27606;
  assign tmp31871 = l1 ? tmp27971 : tmp30018;
  assign tmp31870 = s0 ? tmp28258 : tmp31871;
  assign tmp31868 = s1 ? tmp31869 : tmp31870;
  assign tmp31875 = l1 ? tmp27980 : tmp27833;
  assign tmp31874 = s0 ? tmp31875 : tmp31869;
  assign tmp31877 = l1 ? tmp27971 : tmp27833;
  assign tmp31876 = s0 ? tmp31877 : tmp31869;
  assign tmp31873 = s1 ? tmp31874 : tmp31876;
  assign tmp31879 = s0 ? tmp31877 : tmp28267;
  assign tmp31878 = s1 ? tmp31879 : tmp31869;
  assign tmp31872 = s2 ? tmp31873 : tmp31878;
  assign tmp31867 = s3 ? tmp31868 : tmp31872;
  assign tmp31884 = l1 ? tmp27980 : tmp30018;
  assign tmp31883 = s0 ? tmp31884 : tmp28258;
  assign tmp31882 = s1 ? tmp31883 : tmp31869;
  assign tmp31886 = s0 ? tmp31869 : 1;
  assign tmp31887 = s0 ? tmp31193 : 1;
  assign tmp31885 = s1 ? tmp31886 : tmp31887;
  assign tmp31881 = s2 ? tmp31882 : tmp31885;
  assign tmp31889 = s1 ? tmp28258 : tmp29222;
  assign tmp31892 = ~(l1 ? tmp27971 : tmp27606);
  assign tmp31891 = ~(s0 ? tmp27750 : tmp31892);
  assign tmp31890 = s1 ? tmp31869 : tmp31891;
  assign tmp31888 = s2 ? tmp31889 : tmp31890;
  assign tmp31880 = s3 ? tmp31881 : tmp31888;
  assign tmp31866 = s4 ? tmp31867 : tmp31880;
  assign tmp31898 = s0 ? tmp31871 : tmp28267;
  assign tmp31899 = s0 ? tmp28267 : tmp31875;
  assign tmp31897 = s1 ? tmp31898 : tmp31899;
  assign tmp31902 = l1 ? tmp27971 : tmp27809;
  assign tmp31901 = s0 ? tmp28267 : tmp31902;
  assign tmp31904 = l1 ? tmp28014 : tmp27606;
  assign tmp31903 = s0 ? tmp31904 : tmp28267;
  assign tmp31900 = s1 ? tmp31901 : tmp31903;
  assign tmp31896 = s2 ? tmp31897 : tmp31900;
  assign tmp31908 = l1 ? tmp28014 : tmp27833;
  assign tmp31907 = s0 ? tmp28267 : tmp31908;
  assign tmp31909 = s0 ? tmp28267 : tmp27791;
  assign tmp31906 = s1 ? tmp31907 : tmp31909;
  assign tmp31912 = l1 ? tmp28014 : tmp27809;
  assign tmp31911 = ~(s0 ? tmp31902 : tmp31912);
  assign tmp31910 = ~(s1 ? tmp27750 : tmp31911);
  assign tmp31905 = s2 ? tmp31906 : tmp31910;
  assign tmp31895 = s3 ? tmp31896 : tmp31905;
  assign tmp31917 = ~(l1 ? tmp27971 : tmp27809);
  assign tmp31916 = s0 ? tmp27750 : tmp31917;
  assign tmp31918 = ~(s0 ? tmp31193 : tmp29217);
  assign tmp31915 = s1 ? tmp31916 : tmp31918;
  assign tmp31920 = s0 ? tmp31193 : tmp29217;
  assign tmp31922 = l1 ? tmp27980 : tmp27809;
  assign tmp31921 = s0 ? tmp31922 : tmp31193;
  assign tmp31919 = ~(s1 ? tmp31920 : tmp31921);
  assign tmp31914 = s2 ? tmp31915 : tmp31919;
  assign tmp31926 = ~(l1 ? tmp28014 : tmp27809);
  assign tmp31925 = s0 ? tmp27750 : tmp31926;
  assign tmp31927 = ~(s0 ? tmp29217 : tmp27791);
  assign tmp31924 = s1 ? tmp31925 : tmp31927;
  assign tmp31923 = s2 ? tmp31924 : tmp27750;
  assign tmp31913 = ~(s3 ? tmp31914 : tmp31923);
  assign tmp31894 = s4 ? tmp31895 : tmp31913;
  assign tmp31893 = s5 ? tmp31894 : tmp27791;
  assign tmp31865 = s6 ? tmp31866 : tmp31893;
  assign tmp31864 = s7 ? tmp31865 : tmp27495;
  assign tmp31863 = ~(s8 ? tmp28314 : tmp31864);
  assign tmp31862 = s9 ? tmp28189 : tmp31863;
  assign tmp31929 = s8 ? tmp28314 : tmp28251;
  assign tmp31928 = ~(s9 ? tmp31929 : tmp27495);
  assign tmp31861 = s10 ? tmp31862 : tmp31928;
  assign tmp31860 = s12 ? tmp27877 : tmp31861;
  assign tmp31789 = s13 ? tmp31790 : tmp31860;
  assign tmp31940 = l1 ? tmp27936 : tmp27972;
  assign tmp31942 = l1 ? tmp27517 : tmp27891;
  assign tmp31943 = l1 ? tmp27936 : tmp27490;
  assign tmp31941 = s0 ? tmp31942 : tmp31943;
  assign tmp31939 = s1 ? tmp31940 : tmp31941;
  assign tmp31947 = l1 ? tmp27936 : tmp29414;
  assign tmp31948 = l1 ? tmp27936 : tmp27509;
  assign tmp31946 = s0 ? tmp31947 : tmp31948;
  assign tmp31949 = s0 ? tmp31943 : tmp31948;
  assign tmp31945 = s1 ? tmp31946 : tmp31949;
  assign tmp31951 = s0 ? tmp31943 : tmp29880;
  assign tmp31952 = s0 ? tmp31948 : tmp31940;
  assign tmp31950 = s1 ? tmp31951 : tmp31952;
  assign tmp31944 = s2 ? tmp31945 : tmp31950;
  assign tmp31938 = s3 ? tmp31939 : tmp31944;
  assign tmp31956 = s0 ? tmp31940 : tmp31948;
  assign tmp31955 = s1 ? tmp31951 : tmp31956;
  assign tmp31958 = s0 ? tmp31940 : tmp29880;
  assign tmp31960 = l1 ? tmp27517 : tmp28080;
  assign tmp31959 = s0 ? tmp31960 : tmp29880;
  assign tmp31957 = s1 ? tmp31958 : tmp31959;
  assign tmp31954 = s2 ? tmp31955 : tmp31957;
  assign tmp31962 = s1 ? tmp31942 : tmp29902;
  assign tmp31964 = s0 ? tmp31948 : tmp27509;
  assign tmp31965 = s0 ? tmp27508 : tmp31948;
  assign tmp31963 = s1 ? tmp31964 : tmp31965;
  assign tmp31961 = s2 ? tmp31962 : tmp31963;
  assign tmp31953 = s3 ? tmp31954 : tmp31961;
  assign tmp31937 = s4 ? tmp31938 : tmp31953;
  assign tmp31971 = s0 ? tmp31943 : tmp29907;
  assign tmp31973 = ~(l1 ? tmp27936 : tmp29414);
  assign tmp31972 = ~(s0 ? tmp28446 : tmp31973);
  assign tmp31970 = s1 ? tmp31971 : tmp31972;
  assign tmp31976 = ~(l1 ? tmp27936 : tmp27497);
  assign tmp31975 = s0 ? tmp28446 : tmp31976;
  assign tmp31974 = ~(s1 ? tmp31975 : tmp28468);
  assign tmp31969 = s2 ? tmp31970 : tmp31974;
  assign tmp31979 = s0 ? tmp27495 : tmp31943;
  assign tmp31978 = s1 ? tmp31979 : tmp27935;
  assign tmp31980 = s1 ? tmp27585 : tmp27936;
  assign tmp31977 = s2 ? tmp31978 : tmp31980;
  assign tmp31968 = s3 ? tmp31969 : tmp31977;
  assign tmp31984 = s0 ? 1 : tmp31976;
  assign tmp31986 = l1 ? tmp27517 : tmp27508;
  assign tmp31985 = ~(s0 ? tmp29880 : tmp31986);
  assign tmp31983 = s1 ? tmp31984 : tmp31985;
  assign tmp31988 = s0 ? tmp29880 : tmp31986;
  assign tmp31990 = l1 ? tmp27936 : tmp27497;
  assign tmp31989 = s0 ? tmp31990 : tmp29880;
  assign tmp31987 = ~(s1 ? tmp31988 : tmp31989);
  assign tmp31982 = s2 ? tmp31983 : tmp31987;
  assign tmp31993 = s0 ? tmp27858 : tmp28473;
  assign tmp31994 = ~(s0 ? tmp31986 : 0);
  assign tmp31992 = s1 ? tmp31993 : tmp31994;
  assign tmp31991 = s2 ? tmp31992 : 1;
  assign tmp31981 = ~(s3 ? tmp31982 : tmp31991);
  assign tmp31967 = s4 ? tmp31968 : tmp31981;
  assign tmp31999 = ~(s0 ? 1 : tmp28100);
  assign tmp31998 = s1 ? tmp27956 : tmp31999;
  assign tmp32001 = s0 ? tmp28100 : tmp27959;
  assign tmp32000 = ~(s1 ? tmp32001 : tmp27959);
  assign tmp31997 = s2 ? tmp31998 : tmp32000;
  assign tmp31996 = s3 ? tmp31997 : 0;
  assign tmp32005 = s0 ? 1 : tmp27563;
  assign tmp32004 = s1 ? 1 : tmp32005;
  assign tmp32003 = s2 ? tmp32004 : tmp27963;
  assign tmp32008 = s0 ? tmp28100 : 1;
  assign tmp32007 = s1 ? tmp32008 : 1;
  assign tmp32006 = s2 ? tmp32007 : 1;
  assign tmp32002 = ~(s3 ? tmp32003 : tmp32006);
  assign tmp31995 = s4 ? tmp31996 : tmp32002;
  assign tmp31966 = s5 ? tmp31967 : tmp31995;
  assign tmp31936 = s6 ? tmp31937 : tmp31966;
  assign tmp31935 = s7 ? tmp31936 : tmp27495;
  assign tmp32015 = l2 ? tmp27554 : tmp27509;
  assign tmp32014 = l1 ? tmp28014 : tmp32015;
  assign tmp32017 = l1 ? tmp28014 : tmp28643;
  assign tmp32016 = s0 ? tmp30945 : tmp32017;
  assign tmp32013 = s1 ? tmp32014 : tmp32016;
  assign tmp32021 = l1 ? tmp28014 : tmp27560;
  assign tmp32022 = l1 ? tmp28014 : tmp27971;
  assign tmp32020 = s0 ? tmp32021 : tmp32022;
  assign tmp32023 = s0 ? tmp32017 : tmp32022;
  assign tmp32019 = s1 ? tmp32020 : tmp32023;
  assign tmp32025 = s0 ? tmp32017 : tmp27836;
  assign tmp32026 = s0 ? tmp32022 : tmp32014;
  assign tmp32024 = s1 ? tmp32025 : tmp32026;
  assign tmp32018 = s2 ? tmp32019 : tmp32024;
  assign tmp32012 = s3 ? tmp32013 : tmp32018;
  assign tmp32030 = s0 ? tmp32014 : tmp32022;
  assign tmp32029 = s1 ? tmp32025 : tmp32030;
  assign tmp32032 = s0 ? tmp32014 : tmp27836;
  assign tmp32034 = l1 ? tmp27504 : tmp27554;
  assign tmp32033 = s0 ? tmp32034 : tmp27836;
  assign tmp32031 = s1 ? tmp32032 : tmp32033;
  assign tmp32028 = s2 ? tmp32029 : tmp32031;
  assign tmp32036 = s1 ? tmp30945 : tmp29954;
  assign tmp32038 = s0 ? tmp32022 : tmp27971;
  assign tmp32039 = s0 ? tmp27488 : tmp32022;
  assign tmp32037 = s1 ? tmp32038 : tmp32039;
  assign tmp32035 = s2 ? tmp32036 : tmp32037;
  assign tmp32027 = s3 ? tmp32028 : tmp32035;
  assign tmp32011 = s4 ? tmp32012 : tmp32027;
  assign tmp32045 = s0 ? tmp32017 : tmp29958;
  assign tmp32047 = ~(l1 ? tmp28014 : tmp27560);
  assign tmp32046 = ~(s0 ? tmp27640 : tmp32047);
  assign tmp32044 = s1 ? tmp32045 : tmp32046;
  assign tmp32050 = ~(l1 ? tmp28014 : tmp31492);
  assign tmp32049 = s0 ? tmp27640 : tmp32050;
  assign tmp32051 = ~(s0 ? tmp27971 : 1);
  assign tmp32048 = ~(s1 ? tmp32049 : tmp32051);
  assign tmp32043 = s2 ? tmp32044 : tmp32048;
  assign tmp32054 = s0 ? 1 : tmp32017;
  assign tmp32055 = s0 ? 1 : tmp28014;
  assign tmp32053 = s1 ? tmp32054 : tmp32055;
  assign tmp32056 = s1 ? tmp28533 : tmp28014;
  assign tmp32052 = s2 ? tmp32053 : tmp32056;
  assign tmp32042 = s3 ? tmp32043 : tmp32052;
  assign tmp32060 = s0 ? 1 : tmp32050;
  assign tmp32061 = ~(s0 ? tmp27836 : tmp29118);
  assign tmp32059 = s1 ? tmp32060 : tmp32061;
  assign tmp32063 = s0 ? tmp27836 : tmp29118;
  assign tmp32065 = l1 ? tmp28014 : tmp31492;
  assign tmp32064 = s0 ? tmp32065 : tmp27836;
  assign tmp32062 = ~(s1 ? tmp32063 : tmp32064);
  assign tmp32058 = s2 ? tmp32059 : tmp32062;
  assign tmp32068 = s0 ? tmp28524 : tmp28531;
  assign tmp32069 = ~(s0 ? tmp29118 : 0);
  assign tmp32067 = s1 ? tmp32068 : tmp32069;
  assign tmp32066 = s2 ? tmp32067 : 1;
  assign tmp32057 = ~(s3 ? tmp32058 : tmp32066);
  assign tmp32041 = s4 ? tmp32042 : tmp32057;
  assign tmp32070 = s4 ? tmp28549 : tmp28556;
  assign tmp32040 = s5 ? tmp32041 : tmp32070;
  assign tmp32010 = s6 ? tmp32011 : tmp32040;
  assign tmp32009 = s7 ? tmp32010 : tmp27495;
  assign tmp31934 = s8 ? tmp31935 : tmp32009;
  assign tmp32077 = l1 ? tmp28014 : tmp30069;
  assign tmp32079 = l1 ? tmp28014 : tmp27554;
  assign tmp32078 = s0 ? tmp30945 : tmp32079;
  assign tmp32076 = s1 ? tmp32077 : tmp32078;
  assign tmp32083 = l1 ? tmp28014 : 1;
  assign tmp32084 = l1 ? tmp28014 : tmp27488;
  assign tmp32082 = s0 ? tmp32083 : tmp32084;
  assign tmp32086 = l1 ? tmp28014 : tmp28661;
  assign tmp32085 = s0 ? tmp32086 : tmp32084;
  assign tmp32081 = s1 ? tmp32082 : tmp32085;
  assign tmp32088 = s0 ? tmp32086 : tmp27836;
  assign tmp32089 = s0 ? tmp32084 : tmp32077;
  assign tmp32087 = s1 ? tmp32088 : tmp32089;
  assign tmp32080 = s2 ? tmp32081 : tmp32087;
  assign tmp32075 = s3 ? tmp32076 : tmp32080;
  assign tmp32093 = s0 ? tmp32079 : tmp27836;
  assign tmp32094 = s0 ? tmp32077 : tmp32084;
  assign tmp32092 = s1 ? tmp32093 : tmp32094;
  assign tmp32096 = s0 ? tmp32077 : tmp27836;
  assign tmp32095 = s1 ? tmp32096 : tmp32033;
  assign tmp32091 = s2 ? tmp32092 : tmp32095;
  assign tmp32098 = s1 ? tmp30945 : tmp30032;
  assign tmp32100 = s0 ? tmp27488 : tmp32084;
  assign tmp32099 = s1 ? tmp32084 : tmp32100;
  assign tmp32097 = s2 ? tmp32098 : tmp32099;
  assign tmp32090 = s3 ? tmp32091 : tmp32097;
  assign tmp32074 = s4 ? tmp32075 : tmp32090;
  assign tmp32106 = s0 ? tmp32079 : tmp29958;
  assign tmp32108 = ~(l1 ? tmp28014 : 1);
  assign tmp32107 = ~(s0 ? tmp27640 : tmp32108);
  assign tmp32105 = s1 ? tmp32106 : tmp32107;
  assign tmp32111 = ~(l1 ? tmp28014 : tmp27554);
  assign tmp32110 = s0 ? tmp27640 : tmp32111;
  assign tmp32112 = ~(s0 ? tmp32084 : 1);
  assign tmp32109 = ~(s1 ? tmp32110 : tmp32112);
  assign tmp32104 = s2 ? tmp32105 : tmp32109;
  assign tmp32115 = s0 ? 1 : tmp32086;
  assign tmp32116 = s0 ? 1 : tmp28589;
  assign tmp32114 = s1 ? tmp32115 : tmp32116;
  assign tmp32117 = s1 ? tmp28602 : tmp32084;
  assign tmp32113 = s2 ? tmp32114 : tmp32117;
  assign tmp32103 = s3 ? tmp32104 : tmp32113;
  assign tmp32122 = ~(l1 ? tmp28014 : tmp31489);
  assign tmp32121 = s0 ? tmp27750 : tmp32122;
  assign tmp32120 = s1 ? tmp32121 : tmp32061;
  assign tmp32123 = ~(s1 ? tmp32063 : tmp32093);
  assign tmp32119 = s2 ? tmp32120 : tmp32123;
  assign tmp32128 = l2 ? tmp27488 : tmp27491;
  assign tmp32127 = ~(l1 ? tmp28014 : tmp32128);
  assign tmp32126 = s0 ? tmp28509 : tmp32127;
  assign tmp32129 = ~(s0 ? tmp29118 : tmp27791);
  assign tmp32125 = s1 ? tmp32126 : tmp32129;
  assign tmp32124 = s2 ? tmp32125 : tmp27750;
  assign tmp32118 = ~(s3 ? tmp32119 : tmp32124);
  assign tmp32102 = s4 ? tmp32103 : tmp32118;
  assign tmp32130 = ~(s4 ? tmp28617 : tmp28622);
  assign tmp32101 = s5 ? tmp32102 : tmp32130;
  assign tmp32073 = s6 ? tmp32074 : tmp32101;
  assign tmp32072 = s7 ? tmp32073 : tmp27495;
  assign tmp32071 = s8 ? tmp32009 : tmp32072;
  assign tmp31933 = s9 ? tmp31934 : tmp32071;
  assign tmp32132 = s8 ? tmp32009 : tmp32010;
  assign tmp32131 = s9 ? tmp32132 : tmp27495;
  assign tmp31932 = s10 ? tmp31933 : tmp32131;
  assign tmp32142 = l2 ? tmp27509 : tmp27506;
  assign tmp32141 = l1 ? tmp32142 : tmp28665;
  assign tmp32144 = l1 ? tmp27510 : tmp28665;
  assign tmp32143 = s0 ? tmp29333 : tmp32144;
  assign tmp32140 = s1 ? tmp32141 : tmp32143;
  assign tmp32147 = l1 ? tmp32142 : tmp28490;
  assign tmp32146 = s0 ? tmp32147 : tmp32144;
  assign tmp32149 = s0 ? tmp32147 : tmp30650;
  assign tmp32148 = s1 ? tmp32149 : tmp32144;
  assign tmp32145 = s2 ? tmp32146 : tmp32148;
  assign tmp32139 = s3 ? tmp32140 : tmp32145;
  assign tmp32154 = l1 ? tmp28938 : 0;
  assign tmp32153 = s0 ? tmp32141 : tmp32154;
  assign tmp32152 = s1 ? tmp32153 : tmp32144;
  assign tmp32156 = s0 ? tmp32141 : tmp27517;
  assign tmp32157 = s0 ? tmp29333 : tmp27517;
  assign tmp32155 = s1 ? tmp32156 : tmp32157;
  assign tmp32151 = s2 ? tmp32152 : tmp32155;
  assign tmp32160 = s0 ? tmp27517 : tmp28488;
  assign tmp32159 = s1 ? tmp29333 : tmp32160;
  assign tmp32162 = s0 ? tmp32144 : tmp28680;
  assign tmp32164 = ~(l1 ? tmp27510 : tmp28665);
  assign tmp32163 = ~(s0 ? tmp28667 : tmp32164);
  assign tmp32161 = s1 ? tmp32162 : tmp32163;
  assign tmp32158 = s2 ? tmp32159 : tmp32161;
  assign tmp32150 = s3 ? tmp32151 : tmp32158;
  assign tmp32138 = s4 ? tmp32139 : tmp32150;
  assign tmp32170 = s0 ? tmp32144 : 0;
  assign tmp32172 = ~(l1 ? tmp32142 : tmp28490);
  assign tmp32171 = ~(s0 ? 1 : tmp32172);
  assign tmp32169 = s1 ? tmp32170 : tmp32171;
  assign tmp32175 = ~(l1 ? tmp27510 : tmp28685);
  assign tmp32174 = s0 ? 1 : tmp32175;
  assign tmp32176 = ~(s0 ? tmp28680 : tmp31533);
  assign tmp32173 = ~(s1 ? tmp32174 : tmp32176);
  assign tmp32168 = s2 ? tmp32169 : tmp32173;
  assign tmp32179 = s0 ? tmp31533 : tmp32147;
  assign tmp32180 = s0 ? tmp31533 : tmp28704;
  assign tmp32178 = s1 ? tmp32179 : tmp32180;
  assign tmp32183 = l1 ? tmp27510 : tmp28685;
  assign tmp32182 = ~(s0 ? tmp32183 : tmp28704);
  assign tmp32181 = ~(s1 ? tmp28687 : tmp32182);
  assign tmp32177 = s2 ? tmp32178 : tmp32181;
  assign tmp32167 = s3 ? tmp32168 : tmp32177;
  assign tmp32187 = s0 ? tmp28667 : tmp32175;
  assign tmp32188 = ~(s0 ? tmp32154 : tmp27495);
  assign tmp32186 = s1 ? tmp32187 : tmp32188;
  assign tmp32190 = s0 ? tmp32154 : tmp27495;
  assign tmp32192 = l1 ? tmp32142 : tmp28685;
  assign tmp32191 = s0 ? tmp32192 : tmp32154;
  assign tmp32189 = ~(s1 ? tmp32190 : tmp32191);
  assign tmp32185 = s2 ? tmp32186 : tmp32189;
  assign tmp32196 = ~(l1 ? tmp32142 : tmp28733);
  assign tmp32195 = s0 ? tmp28700 : tmp32196;
  assign tmp32194 = s1 ? tmp32195 : tmp28703;
  assign tmp32193 = s2 ? tmp32194 : tmp28705;
  assign tmp32184 = ~(s3 ? tmp32185 : tmp32193);
  assign tmp32166 = s4 ? tmp32167 : tmp32184;
  assign tmp32202 = l1 ? tmp27504 : tmp31492;
  assign tmp32201 = s0 ? tmp28446 : tmp32202;
  assign tmp32203 = s0 ? tmp27588 : tmp32202;
  assign tmp32200 = ~(s1 ? tmp32201 : tmp32203);
  assign tmp32199 = s2 ? tmp28710 : tmp32200;
  assign tmp32198 = s3 ? tmp32199 : tmp28716;
  assign tmp32207 = s0 ? tmp32202 : tmp27588;
  assign tmp32206 = s1 ? tmp28726 : tmp32207;
  assign tmp32205 = s2 ? tmp28722 : tmp32206;
  assign tmp32204 = ~(s3 ? tmp32205 : tmp28729);
  assign tmp32197 = s4 ? tmp32198 : tmp32204;
  assign tmp32165 = s5 ? tmp32166 : tmp32197;
  assign tmp32137 = s6 ? tmp32138 : tmp32165;
  assign tmp32136 = s7 ? tmp32137 : tmp27495;
  assign tmp32214 = ~(l2 ? tmp27490 : tmp27496);
  assign tmp32213 = l1 ? tmp27665 : tmp32214;
  assign tmp32216 = l1 ? tmp32128 : tmp32214;
  assign tmp32215 = s0 ? tmp27909 : tmp32216;
  assign tmp32212 = s1 ? tmp32213 : tmp32215;
  assign tmp32219 = l1 ? tmp27665 : tmp27506;
  assign tmp32218 = s0 ? tmp32219 : tmp32216;
  assign tmp32221 = s0 ? tmp32219 : tmp27838;
  assign tmp32220 = s1 ? tmp32221 : tmp32216;
  assign tmp32217 = s2 ? tmp32218 : tmp32220;
  assign tmp32211 = s3 ? tmp32212 : tmp32217;
  assign tmp32226 = l1 ? tmp27897 : 0;
  assign tmp32225 = s0 ? tmp32213 : tmp32226;
  assign tmp32224 = s1 ? tmp32225 : tmp32216;
  assign tmp32228 = s0 ? tmp32213 : tmp27504;
  assign tmp32229 = s0 ? tmp27909 : tmp27504;
  assign tmp32227 = s1 ? tmp32228 : tmp32229;
  assign tmp32223 = s2 ? tmp32224 : tmp32227;
  assign tmp32232 = s0 ? tmp27504 : tmp27695;
  assign tmp32231 = s1 ? tmp27909 : tmp32232;
  assign tmp32235 = l1 ? tmp27488 : tmp32214;
  assign tmp32234 = s0 ? tmp32216 : tmp32235;
  assign tmp32237 = ~(l1 ? tmp32128 : tmp32214);
  assign tmp32236 = ~(s0 ? tmp27985 : tmp32237);
  assign tmp32233 = s1 ? tmp32234 : tmp32236;
  assign tmp32230 = s2 ? tmp32231 : tmp32233;
  assign tmp32222 = s3 ? tmp32223 : tmp32230;
  assign tmp32210 = s4 ? tmp32211 : tmp32222;
  assign tmp32243 = s0 ? tmp32216 : 0;
  assign tmp32245 = ~(l1 ? tmp27665 : tmp27506);
  assign tmp32244 = ~(s0 ? 1 : tmp32245);
  assign tmp32242 = s1 ? tmp32243 : tmp32244;
  assign tmp32248 = ~(l1 ? tmp32128 : tmp28802);
  assign tmp32247 = s0 ? 1 : tmp32248;
  assign tmp32249 = ~(s0 ? tmp32235 : tmp28033);
  assign tmp32246 = ~(s1 ? tmp32247 : tmp32249);
  assign tmp32241 = s2 ? tmp32242 : tmp32246;
  assign tmp32252 = s0 ? tmp28033 : tmp32219;
  assign tmp32254 = l1 ? tmp27488 : tmp28802;
  assign tmp32253 = s0 ? tmp28033 : tmp32254;
  assign tmp32251 = s1 ? tmp32252 : tmp32253;
  assign tmp32256 = s0 ? tmp27985 : 1;
  assign tmp32258 = l1 ? tmp32128 : tmp28802;
  assign tmp32257 = ~(s0 ? tmp32258 : tmp32254);
  assign tmp32255 = ~(s1 ? tmp32256 : tmp32257);
  assign tmp32250 = s2 ? tmp32251 : tmp32255;
  assign tmp32240 = s3 ? tmp32241 : tmp32250;
  assign tmp32262 = s0 ? tmp27985 : tmp32248;
  assign tmp32263 = ~(s0 ? tmp32226 : 1);
  assign tmp32261 = s1 ? tmp32262 : tmp32263;
  assign tmp32265 = s0 ? tmp32226 : 1;
  assign tmp32267 = l1 ? tmp27665 : tmp28802;
  assign tmp32266 = s0 ? tmp32267 : tmp32226;
  assign tmp32264 = ~(s1 ? tmp32265 : tmp32266);
  assign tmp32260 = s2 ? tmp32261 : tmp32264;
  assign tmp32271 = l1 ? tmp27504 : tmp29088;
  assign tmp32272 = ~(l1 ? tmp27665 : tmp28835);
  assign tmp32270 = s0 ? tmp32271 : tmp32272;
  assign tmp32273 = ~(s0 ? 1 : tmp32254);
  assign tmp32269 = s1 ? tmp32270 : tmp32273;
  assign tmp32268 = s2 ? tmp32269 : tmp28803;
  assign tmp32259 = ~(s3 ? tmp32260 : tmp32268);
  assign tmp32239 = s4 ? tmp32240 : tmp32259;
  assign tmp32278 = s0 ? tmp32254 : 0;
  assign tmp32277 = s1 ? tmp32278 : tmp27675;
  assign tmp32281 = l1 ? tmp27504 : tmp27497;
  assign tmp32280 = s0 ? tmp27640 : tmp32281;
  assign tmp32282 = s0 ? tmp27697 : tmp32281;
  assign tmp32279 = ~(s1 ? tmp32280 : tmp32282);
  assign tmp32276 = s2 ? tmp32277 : tmp32279;
  assign tmp32275 = s3 ? tmp32276 : tmp28816;
  assign tmp32285 = s1 ? tmp28825 : tmp29307;
  assign tmp32288 = l1 ? tmp27499 : tmp29088;
  assign tmp32287 = s0 ? 1 : tmp32288;
  assign tmp32289 = s0 ? tmp32281 : tmp27697;
  assign tmp32286 = s1 ? tmp32287 : tmp32289;
  assign tmp32284 = s2 ? tmp32285 : tmp32286;
  assign tmp32291 = s1 ? tmp28512 : tmp28833;
  assign tmp32290 = s2 ? tmp32291 : tmp28836;
  assign tmp32283 = ~(s3 ? tmp32284 : tmp32290);
  assign tmp32274 = s4 ? tmp32275 : tmp32283;
  assign tmp32238 = s5 ? tmp32239 : tmp32274;
  assign tmp32209 = s6 ? tmp32210 : tmp32238;
  assign tmp32208 = s7 ? tmp32209 : tmp27495;
  assign tmp32135 = s8 ? tmp32136 : tmp32208;
  assign tmp32300 = l1 ? tmp27897 : tmp27809;
  assign tmp32299 = s0 ? tmp32213 : tmp32300;
  assign tmp32298 = s1 ? tmp32299 : tmp32216;
  assign tmp32302 = s0 ? tmp32213 : tmp29180;
  assign tmp32303 = s0 ? tmp27909 : tmp29180;
  assign tmp32301 = s1 ? tmp32302 : tmp32303;
  assign tmp32297 = s2 ? tmp32298 : tmp32301;
  assign tmp32307 = ~(l1 ? tmp27891 : tmp28860);
  assign tmp32306 = s0 ? tmp29180 : tmp32307;
  assign tmp32305 = s1 ? tmp27909 : tmp32306;
  assign tmp32309 = ~(s0 ? tmp28884 : tmp32237);
  assign tmp32308 = s1 ? tmp32234 : tmp32309;
  assign tmp32304 = s2 ? tmp32305 : tmp32308;
  assign tmp32296 = s3 ? tmp32297 : tmp32304;
  assign tmp32295 = s4 ? tmp32211 : tmp32296;
  assign tmp32315 = s0 ? tmp32216 : tmp27791;
  assign tmp32316 = ~(s0 ? tmp27750 : tmp32245);
  assign tmp32314 = s1 ? tmp32315 : tmp32316;
  assign tmp32318 = s0 ? tmp27750 : tmp32248;
  assign tmp32317 = ~(s1 ? tmp32318 : tmp32249);
  assign tmp32313 = s2 ? tmp32314 : tmp32317;
  assign tmp32321 = s0 ? tmp28884 : tmp27750;
  assign tmp32320 = ~(s1 ? tmp32321 : tmp32257);
  assign tmp32319 = s2 ? tmp32251 : tmp32320;
  assign tmp32312 = s3 ? tmp32313 : tmp32319;
  assign tmp32325 = s0 ? tmp28884 : tmp32248;
  assign tmp32326 = ~(s0 ? tmp32300 : 1);
  assign tmp32324 = s1 ? tmp32325 : tmp32326;
  assign tmp32328 = s0 ? tmp32300 : 1;
  assign tmp32329 = s0 ? tmp32267 : tmp32300;
  assign tmp32327 = ~(s1 ? tmp32328 : tmp32329);
  assign tmp32323 = s2 ? tmp32324 : tmp32327;
  assign tmp32330 = s2 ? tmp32269 : tmp28889;
  assign tmp32322 = ~(s3 ? tmp32323 : tmp32330);
  assign tmp32311 = s4 ? tmp32312 : tmp32322;
  assign tmp32335 = s0 ? tmp32254 : tmp27791;
  assign tmp32336 = ~(s0 ? tmp27750 : tmp27640);
  assign tmp32334 = s1 ? tmp32335 : tmp32336;
  assign tmp32333 = s2 ? tmp32334 : tmp32279;
  assign tmp32332 = s3 ? tmp32333 : tmp28900;
  assign tmp32340 = s0 ? tmp27750 : tmp28884;
  assign tmp32339 = s1 ? tmp28910 : tmp32340;
  assign tmp32342 = s0 ? tmp27750 : tmp32288;
  assign tmp32341 = s1 ? tmp32342 : tmp32289;
  assign tmp32338 = s2 ? tmp32339 : tmp32341;
  assign tmp32344 = s1 ? tmp28586 : tmp28917;
  assign tmp32343 = s2 ? tmp32344 : tmp28918;
  assign tmp32337 = ~(s3 ? tmp32338 : tmp32343);
  assign tmp32331 = s4 ? tmp32332 : tmp32337;
  assign tmp32310 = s5 ? tmp32311 : tmp32331;
  assign tmp32294 = s6 ? tmp32295 : tmp32310;
  assign tmp32293 = s7 ? tmp32294 : tmp27495;
  assign tmp32292 = s8 ? tmp32208 : tmp32293;
  assign tmp32134 = s9 ? tmp32135 : tmp32292;
  assign tmp32346 = s8 ? tmp32208 : tmp32209;
  assign tmp32345 = s9 ? tmp32346 : tmp27495;
  assign tmp32133 = s10 ? tmp32134 : tmp32345;
  assign tmp31931 = s12 ? tmp31932 : tmp32133;
  assign tmp32357 = l1 ? tmp27560 : tmp28608;
  assign tmp32356 = s0 ? tmp32357 : tmp29041;
  assign tmp32355 = s1 ? tmp29038 : tmp32356;
  assign tmp32360 = s0 ? tmp29047 : tmp28905;
  assign tmp32359 = s1 ? tmp32360 : tmp29051;
  assign tmp32358 = s2 ? tmp29043 : tmp32359;
  assign tmp32354 = s3 ? tmp32355 : tmp32358;
  assign tmp32364 = s0 ? tmp29057 : tmp29160;
  assign tmp32363 = s1 ? tmp32364 : tmp29058;
  assign tmp32366 = s0 ? tmp29038 : tmp27750;
  assign tmp32367 = s0 ? tmp29062 : tmp27750;
  assign tmp32365 = s1 ? tmp32366 : tmp32367;
  assign tmp32362 = s2 ? tmp32363 : tmp32365;
  assign tmp32370 = s0 ? tmp29062 : tmp32357;
  assign tmp32369 = s1 ? tmp32370 : tmp27750;
  assign tmp32368 = s2 ? tmp32369 : tmp29066;
  assign tmp32361 = s3 ? tmp32362 : tmp32368;
  assign tmp32353 = s4 ? tmp32354 : tmp32361;
  assign tmp32376 = s0 ? tmp29041 : tmp29178;
  assign tmp32377 = ~(s0 ? tmp29180 : tmp29078);
  assign tmp32375 = s1 ? tmp32376 : tmp32377;
  assign tmp32379 = s0 ? tmp29180 : tmp29081;
  assign tmp32380 = ~(s0 ? tmp29068 : tmp28905);
  assign tmp32378 = ~(s1 ? tmp32379 : tmp32380);
  assign tmp32374 = s2 ? tmp32375 : tmp32378;
  assign tmp32383 = s0 ? tmp28905 : tmp29047;
  assign tmp32384 = s0 ? tmp28905 : tmp29087;
  assign tmp32382 = s1 ? tmp32383 : tmp32384;
  assign tmp32386 = s0 ? tmp29070 : tmp27750;
  assign tmp32385 = s1 ? tmp32386 : tmp29091;
  assign tmp32381 = s2 ? tmp32382 : tmp32385;
  assign tmp32373 = s3 ? tmp32374 : tmp32381;
  assign tmp32390 = s0 ? tmp27750 : tmp29098;
  assign tmp32389 = s1 ? tmp32390 : tmp29099;
  assign tmp32388 = s2 ? tmp32389 : tmp29100;
  assign tmp32391 = ~(s2 ? tmp29104 : tmp27791);
  assign tmp32387 = s3 ? tmp32388 : tmp32391;
  assign tmp32372 = s4 ? tmp32373 : tmp32387;
  assign tmp32396 = s0 ? tmp29087 : tmp27750;
  assign tmp32397 = s0 ? tmp27750 : tmp29115;
  assign tmp32395 = s1 ? tmp32396 : tmp32397;
  assign tmp32394 = s2 ? tmp32395 : tmp29116;
  assign tmp32400 = s0 ? tmp27750 : tmp29123;
  assign tmp32399 = ~(s1 ? tmp27750 : tmp32400);
  assign tmp32398 = ~(s2 ? tmp29221 : tmp32399);
  assign tmp32393 = s3 ? tmp32394 : tmp32398;
  assign tmp32404 = s0 ? tmp28812 : tmp29217;
  assign tmp32405 = s0 ? tmp29217 : tmp29129;
  assign tmp32403 = s1 ? tmp32404 : tmp32405;
  assign tmp32407 = s0 ? tmp27750 : tmp29132;
  assign tmp32406 = ~(s1 ? tmp32407 : 0);
  assign tmp32402 = s2 ? tmp32403 : tmp32406;
  assign tmp32410 = s0 ? tmp29118 : tmp29217;
  assign tmp32411 = ~(s0 ? tmp27750 : tmp29137);
  assign tmp32409 = s1 ? tmp32410 : tmp32411;
  assign tmp32412 = ~(s1 ? tmp32400 : tmp29213);
  assign tmp32408 = s2 ? tmp32409 : tmp32412;
  assign tmp32401 = ~(s3 ? tmp32402 : tmp32408);
  assign tmp32392 = s4 ? tmp32393 : tmp32401;
  assign tmp32371 = s5 ? tmp32372 : tmp32392;
  assign tmp32352 = s6 ? tmp32353 : tmp32371;
  assign tmp32351 = s7 ? tmp32352 : tmp27575;
  assign tmp32350 = s8 ? tmp29033 : tmp32351;
  assign tmp32349 = s9 ? tmp28924 : tmp32350;
  assign tmp32414 = s8 ? tmp29033 : tmp29034;
  assign tmp32413 = s9 ? tmp32414 : tmp27575;
  assign tmp32348 = s10 ? tmp32349 : tmp32413;
  assign tmp32347 = ~(s12 ? tmp32348 : tmp29319);
  assign tmp31930 = ~(s13 ? tmp31931 : tmp32347);
  assign tmp31788 = s14 ? tmp31789 : tmp31930;
  assign tmp32427 = s0 ? tmp31011 : tmp27750;
  assign tmp32426 = s1 ? tmp32427 : tmp31004;
  assign tmp32429 = s0 ? tmp30998 : tmp27750;
  assign tmp32428 = s1 ? tmp32429 : tmp30797;
  assign tmp32425 = s2 ? tmp32426 : tmp32428;
  assign tmp32431 = s1 ? tmp27642 : tmp31123;
  assign tmp32433 = s0 ? tmp31159 : tmp31004;
  assign tmp32432 = s1 ? tmp31019 : tmp32433;
  assign tmp32430 = s2 ? tmp32431 : tmp32432;
  assign tmp32424 = s3 ? tmp32425 : tmp32430;
  assign tmp32423 = s4 ? tmp30996 : tmp32424;
  assign tmp32439 = s0 ? tmp31000 : tmp27750;
  assign tmp32440 = s0 ? tmp27750 : tmp31030;
  assign tmp32438 = s1 ? tmp32439 : tmp32440;
  assign tmp32442 = s0 ? tmp27750 : tmp31033;
  assign tmp32441 = s1 ? tmp32442 : tmp31034;
  assign tmp32437 = s2 ? tmp32438 : tmp32441;
  assign tmp32445 = s0 ? tmp31159 : tmp28378;
  assign tmp32444 = s1 ? tmp32445 : tmp31043;
  assign tmp32443 = s2 ? tmp31036 : tmp32444;
  assign tmp32436 = s3 ? tmp32437 : tmp32443;
  assign tmp32449 = s0 ? tmp31151 : tmp31044;
  assign tmp32448 = s1 ? tmp32449 : tmp30325;
  assign tmp32451 = s0 ? tmp31053 : tmp27750;
  assign tmp32450 = s1 ? tmp30325 : tmp32451;
  assign tmp32447 = s2 ? tmp32448 : tmp32450;
  assign tmp32452 = ~(s2 ? tmp31055 : tmp31160);
  assign tmp32446 = s3 ? tmp32447 : tmp32452;
  assign tmp32435 = s4 ? tmp32436 : tmp32446;
  assign tmp32456 = s1 ? tmp30032 : tmp29838;
  assign tmp32458 = ~(s0 ? tmp27738 : tmp31077);
  assign tmp32457 = s1 ? tmp31175 : tmp32458;
  assign tmp32455 = ~(s2 ? tmp32456 : tmp32457);
  assign tmp32454 = s3 ? tmp31064 : tmp32455;
  assign tmp32462 = s0 ? tmp31082 : tmp31182;
  assign tmp32464 = ~(l1 ? tmp27624 : tmp28860);
  assign tmp32463 = s0 ? tmp31182 : tmp32464;
  assign tmp32461 = s1 ? tmp32462 : tmp32463;
  assign tmp32460 = s2 ? tmp32461 : tmp31085;
  assign tmp32467 = s0 ? 1 : tmp31193;
  assign tmp32468 = s0 ? tmp28342 : tmp31093;
  assign tmp32466 = s1 ? tmp32467 : tmp32468;
  assign tmp32470 = s0 ? tmp27738 : tmp31077;
  assign tmp32469 = ~(s1 ? tmp32470 : tmp31198);
  assign tmp32465 = s2 ? tmp32466 : tmp32469;
  assign tmp32459 = ~(s3 ? tmp32460 : tmp32465);
  assign tmp32453 = s4 ? tmp32454 : tmp32459;
  assign tmp32434 = s5 ? tmp32435 : tmp32453;
  assign tmp32422 = s6 ? tmp32423 : tmp32434;
  assign tmp32421 = s7 ? tmp32422 : tmp27575;
  assign tmp32420 = s8 ? tmp30993 : tmp32421;
  assign tmp32419 = s9 ? tmp30885 : tmp32420;
  assign tmp32472 = s8 ? tmp30993 : tmp30994;
  assign tmp32471 = s9 ? tmp32472 : tmp27575;
  assign tmp32418 = s10 ? tmp32419 : tmp32471;
  assign tmp32417 = s12 ? tmp30563 : tmp32418;
  assign tmp32416 = ~(s13 ? tmp32417 : tmp31280);
  assign tmp32415 = ~(s14 ? tmp29602 : tmp32416);
  assign tmp31787 = s15 ? tmp31788 : tmp32415;
  assign tmp27473 = s16 ? tmp27474 : tmp31787;
  assign tmp32481 = ~(s7 ? tmp28565 : tmp27575);
  assign tmp32480 = s8 ? tmp32009 : tmp32481;
  assign tmp32479 = s9 ? tmp31934 : tmp32480;
  assign tmp32482 = ~(s9 ? tmp28631 : tmp27575);
  assign tmp32478 = s10 ? tmp32479 : tmp32482;
  assign tmp32492 = s0 ? tmp27784 : tmp28644;
  assign tmp32493 = s0 ? tmp28740 : tmp28644;
  assign tmp32491 = s1 ? tmp32492 : tmp32493;
  assign tmp32494 = s1 ? tmp28852 : tmp28752;
  assign tmp32490 = s2 ? tmp32491 : tmp32494;
  assign tmp32489 = s3 ? tmp28842 : tmp32490;
  assign tmp32488 = s4 ? tmp32489 : tmp28847;
  assign tmp32500 = s0 ? tmp27750 : tmp27784;
  assign tmp32499 = s1 ? tmp28869 : tmp32500;
  assign tmp32502 = s0 ? tmp27750 : tmp28744;
  assign tmp32501 = s1 ? tmp32502 : tmp28873;
  assign tmp32498 = s2 ? tmp32499 : tmp32501;
  assign tmp32505 = s0 ? tmp27750 : tmp28740;
  assign tmp32507 = ~(l1 ? tmp27488 : tmp28665);
  assign tmp32506 = s0 ? tmp27750 : tmp32507;
  assign tmp32504 = s1 ? tmp32505 : tmp32506;
  assign tmp32508 = s1 ? tmp28879 : tmp28767;
  assign tmp32503 = s2 ? tmp32504 : tmp32508;
  assign tmp32497 = s3 ? tmp32498 : tmp32503;
  assign tmp32512 = s0 ? tmp28884 : tmp28744;
  assign tmp32511 = s1 ? tmp32512 : tmp28885;
  assign tmp32513 = s1 ? tmp28885 : tmp28850;
  assign tmp32510 = s2 ? tmp32511 : tmp32513;
  assign tmp32517 = l1 ? tmp27504 : tmp28741;
  assign tmp32516 = s0 ? tmp32517 : tmp28740;
  assign tmp32519 = ~(l1 ? tmp27488 : tmp32214);
  assign tmp32518 = s0 ? tmp28014 : tmp32519;
  assign tmp32515 = s1 ? tmp32516 : tmp32518;
  assign tmp32514 = s2 ? tmp32515 : tmp28889;
  assign tmp32509 = s3 ? tmp32510 : tmp32514;
  assign tmp32496 = s4 ? tmp32497 : tmp32509;
  assign tmp32525 = l1 ? tmp27488 : tmp28665;
  assign tmp32524 = s0 ? tmp32525 : tmp27791;
  assign tmp32523 = s1 ? tmp32524 : tmp28896;
  assign tmp32527 = s0 ? tmp28897 : tmp27743;
  assign tmp32528 = s0 ? tmp27504 : tmp27743;
  assign tmp32526 = ~(s1 ? tmp32527 : tmp32528);
  assign tmp32522 = s2 ? tmp32523 : tmp32526;
  assign tmp32531 = s0 ? tmp28905 : tmp27738;
  assign tmp32530 = s1 ? tmp28904 : tmp32531;
  assign tmp32529 = ~(s2 ? tmp27796 : tmp32530);
  assign tmp32521 = s3 ? tmp32522 : tmp32529;
  assign tmp32535 = s0 ? tmp27738 : tmp27750;
  assign tmp32534 = s1 ? tmp32535 : tmp28911;
  assign tmp32538 = l1 ? tmp27499 : tmp28741;
  assign tmp32537 = s0 ? tmp27750 : tmp32538;
  assign tmp32539 = s0 ? tmp27743 : tmp27504;
  assign tmp32536 = s1 ? tmp32537 : tmp32539;
  assign tmp32533 = s2 ? tmp32534 : tmp32536;
  assign tmp32543 = ~(l1 ? tmp27488 : tmp27760);
  assign tmp32542 = s0 ? tmp27750 : tmp32543;
  assign tmp32541 = s1 ? tmp28916 : tmp32542;
  assign tmp32544 = s1 ? tmp32531 : tmp27750;
  assign tmp32540 = s2 ? tmp32541 : tmp32544;
  assign tmp32532 = ~(s3 ? tmp32533 : tmp32540);
  assign tmp32520 = ~(s4 ? tmp32521 : tmp32532);
  assign tmp32495 = s5 ? tmp32496 : tmp32520;
  assign tmp32487 = s6 ? tmp32488 : tmp32495;
  assign tmp32486 = ~(s7 ? tmp32487 : tmp27575);
  assign tmp32485 = s8 ? tmp32208 : tmp32486;
  assign tmp32484 = s9 ? tmp32135 : tmp32485;
  assign tmp32545 = ~(s9 ? tmp28920 : tmp27575);
  assign tmp32483 = s10 ? tmp32484 : tmp32545;
  assign tmp32477 = s12 ? tmp32478 : tmp32483;
  assign tmp32546 = ~(s12 ? tmp28922 : tmp29319);
  assign tmp32476 = ~(s13 ? tmp32477 : tmp32546);
  assign tmp32475 = s14 ? tmp27476 : tmp32476;
  assign tmp32474 = s15 ? tmp32475 : tmp29601;
  assign tmp32473 = s16 ? tmp32474 : tmp31787;
  assign tmp27472 = s17 ? tmp27473 : tmp32473;
  assign s7n = tmp27472;

  assign tmp32561 = l4 ? 1 : 0;
  assign tmp32560 = l3 ? tmp32561 : 0;
  assign tmp32562 = ~(l3 ? 1 : tmp32561);
  assign tmp32559 = l2 ? tmp32560 : tmp32562;
  assign tmp32564 = l3 ? 1 : 0;
  assign tmp32563 = l2 ? tmp32564 : tmp32560;
  assign tmp32558 = l1 ? tmp32559 : tmp32563;
  assign tmp32569 = ~(l4 ? 1 : 0);
  assign tmp32568 = l3 ? 1 : tmp32569;
  assign tmp32567 = l2 ? tmp32568 : tmp32569;
  assign tmp32570 = l2 ? tmp32564 : 1;
  assign tmp32566 = l1 ? tmp32567 : tmp32570;
  assign tmp32572 = l2 ? tmp32564 : 0;
  assign tmp32571 = l1 ? tmp32572 : tmp32564;
  assign tmp32565 = s0 ? tmp32566 : tmp32571;
  assign tmp32557 = s1 ? tmp32558 : tmp32565;
  assign tmp32577 = l2 ? tmp32564 : tmp32569;
  assign tmp32579 = ~(l3 ? 1 : tmp32569);
  assign tmp32578 = ~(l2 ? tmp32561 : tmp32579);
  assign tmp32576 = l1 ? tmp32577 : tmp32578;
  assign tmp32581 = l2 ? tmp32560 : 0;
  assign tmp32583 = ~(l3 ? tmp32561 : 0);
  assign tmp32582 = ~(l2 ? 1 : tmp32583);
  assign tmp32580 = l1 ? tmp32581 : tmp32582;
  assign tmp32575 = s0 ? tmp32576 : tmp32580;
  assign tmp32586 = l2 ? tmp32564 : tmp32562;
  assign tmp32587 = l2 ? tmp32564 : tmp32568;
  assign tmp32585 = l1 ? tmp32586 : tmp32587;
  assign tmp32584 = s0 ? tmp32585 : tmp32580;
  assign tmp32574 = s1 ? tmp32575 : tmp32584;
  assign tmp32591 = l2 ? tmp32568 : tmp32583;
  assign tmp32592 = ~(l2 ? tmp32561 : 0);
  assign tmp32590 = l1 ? tmp32591 : tmp32592;
  assign tmp32589 = s0 ? tmp32585 : tmp32590;
  assign tmp32594 = l1 ? tmp32581 : tmp32563;
  assign tmp32593 = s0 ? tmp32580 : tmp32594;
  assign tmp32588 = s1 ? tmp32589 : tmp32593;
  assign tmp32573 = s2 ? tmp32574 : tmp32588;
  assign tmp32556 = s3 ? tmp32557 : tmp32573;
  assign tmp32599 = l1 ? tmp32577 : tmp32564;
  assign tmp32601 = ~(l2 ? tmp32560 : 0);
  assign tmp32600 = l1 ? tmp32567 : tmp32601;
  assign tmp32598 = s0 ? tmp32599 : tmp32600;
  assign tmp32602 = s0 ? tmp32594 : tmp32580;
  assign tmp32597 = s1 ? tmp32598 : tmp32602;
  assign tmp32605 = l1 ? tmp32591 : 1;
  assign tmp32604 = s0 ? tmp32558 : tmp32605;
  assign tmp32609 = l3 ? tmp32561 : 1;
  assign tmp32608 = ~(l2 ? tmp32609 : 0);
  assign tmp32607 = l1 ? tmp32567 : tmp32608;
  assign tmp32606 = s0 ? tmp32607 : tmp32605;
  assign tmp32603 = s1 ? tmp32604 : tmp32606;
  assign tmp32596 = s2 ? tmp32597 : tmp32603;
  assign tmp32612 = s0 ? tmp32605 : 0;
  assign tmp32611 = s1 ? tmp32607 : tmp32612;
  assign tmp32615 = l1 ? tmp32560 : tmp32582;
  assign tmp32614 = s0 ? tmp32580 : tmp32615;
  assign tmp32617 = ~(l1 ? tmp32581 : tmp32582);
  assign tmp32616 = ~(s0 ? 1 : tmp32617);
  assign tmp32613 = s1 ? tmp32614 : tmp32616;
  assign tmp32610 = s2 ? tmp32611 : tmp32613;
  assign tmp32595 = s3 ? tmp32596 : tmp32610;
  assign tmp32555 = s4 ? tmp32556 : tmp32595;
  assign tmp32625 = l2 ? 1 : tmp32583;
  assign tmp32624 = l1 ? tmp32625 : tmp32601;
  assign tmp32623 = s0 ? tmp32571 : tmp32624;
  assign tmp32626 = s0 ? tmp32624 : tmp32576;
  assign tmp32622 = s1 ? tmp32623 : tmp32626;
  assign tmp32631 = ~(l3 ? 1 : 0);
  assign tmp32630 = ~(l2 ? tmp32609 : tmp32631);
  assign tmp32629 = l1 ? tmp32572 : tmp32630;
  assign tmp32628 = s0 ? tmp32624 : tmp32629;
  assign tmp32634 = l2 ? tmp32568 : 1;
  assign tmp32633 = l1 ? tmp32634 : tmp32592;
  assign tmp32632 = s0 ? tmp32615 : tmp32633;
  assign tmp32627 = s1 ? tmp32628 : tmp32632;
  assign tmp32621 = s2 ? tmp32622 : tmp32627;
  assign tmp32640 = l3 ? tmp32561 : tmp32569;
  assign tmp32639 = l2 ? tmp32564 : tmp32640;
  assign tmp32638 = l1 ? tmp32639 : tmp32587;
  assign tmp32637 = s0 ? tmp32633 : tmp32638;
  assign tmp32641 = s0 ? tmp32633 : 0;
  assign tmp32636 = s1 ? tmp32637 : tmp32641;
  assign tmp32645 = l2 ? tmp32609 : tmp32561;
  assign tmp32644 = ~(l1 ? tmp32645 : tmp32609);
  assign tmp32643 = s0 ? 1 : tmp32644;
  assign tmp32646 = ~(s0 ? tmp32580 : tmp32560);
  assign tmp32642 = ~(s1 ? tmp32643 : tmp32646);
  assign tmp32635 = s2 ? tmp32636 : tmp32642;
  assign tmp32620 = s3 ? tmp32621 : tmp32635;
  assign tmp32651 = l1 ? tmp32609 : tmp32561;
  assign tmp32653 = ~(l2 ? tmp32609 : tmp32583);
  assign tmp32652 = l1 ? tmp32581 : tmp32653;
  assign tmp32650 = s0 ? tmp32651 : tmp32652;
  assign tmp32649 = s1 ? tmp32650 : 0;
  assign tmp32648 = s2 ? tmp32649 : 0;
  assign tmp32647 = s3 ? tmp32648 : 0;
  assign tmp32619 = s4 ? tmp32620 : tmp32647;
  assign tmp32618 = s5 ? tmp32619 : 0;
  assign tmp32554 = s6 ? tmp32555 : tmp32618;
  assign tmp32658 = s1 ? tmp32604 : tmp32607;
  assign tmp32657 = s2 ? tmp32597 : tmp32658;
  assign tmp32660 = s1 ? tmp32566 : 0;
  assign tmp32659 = s2 ? tmp32660 : tmp32613;
  assign tmp32656 = s3 ? tmp32657 : tmp32659;
  assign tmp32655 = s4 ? tmp32556 : tmp32656;
  assign tmp32665 = s1 ? tmp32623 : tmp32576;
  assign tmp32666 = s1 ? tmp32629 : tmp32632;
  assign tmp32664 = s2 ? tmp32665 : tmp32666;
  assign tmp32668 = s1 ? tmp32638 : 0;
  assign tmp32667 = s2 ? tmp32668 : tmp32642;
  assign tmp32663 = s3 ? tmp32664 : tmp32667;
  assign tmp32662 = s4 ? tmp32663 : tmp32647;
  assign tmp32661 = s5 ? tmp32662 : 0;
  assign tmp32654 = s6 ? tmp32655 : tmp32661;
  assign tmp32553 = s7 ? tmp32554 : tmp32654;
  assign tmp32670 = s8 ? tmp32553 : tmp32554;
  assign tmp32669 = s9 ? tmp32670 : tmp32654;
  assign tmp32552 = s10 ? tmp32553 : tmp32669;
  assign tmp32681 = s1 ? tmp32566 : tmp32612;
  assign tmp32680 = s2 ? tmp32681 : tmp32613;
  assign tmp32679 = s3 ? tmp32596 : tmp32680;
  assign tmp32678 = s4 ? tmp32556 : tmp32679;
  assign tmp32677 = s6 ? tmp32678 : tmp32618;
  assign tmp32676 = s7 ? tmp32554 : tmp32677;
  assign tmp32686 = s3 ? tmp32621 : tmp32667;
  assign tmp32685 = s4 ? tmp32686 : tmp32647;
  assign tmp32684 = s5 ? tmp32685 : 0;
  assign tmp32683 = s6 ? tmp32655 : tmp32684;
  assign tmp32682 = s7 ? tmp32554 : tmp32683;
  assign tmp32675 = s8 ? tmp32676 : tmp32682;
  assign tmp32674 = s9 ? tmp32675 : tmp32682;
  assign tmp32688 = s8 ? tmp32682 : tmp32554;
  assign tmp32693 = s3 ? tmp32596 : tmp32659;
  assign tmp32692 = s4 ? tmp32556 : tmp32693;
  assign tmp32697 = s2 ? tmp32622 : tmp32666;
  assign tmp32699 = s1 ? tmp32637 : 0;
  assign tmp32698 = s2 ? tmp32699 : tmp32642;
  assign tmp32696 = s3 ? tmp32697 : tmp32698;
  assign tmp32695 = s4 ? tmp32696 : tmp32647;
  assign tmp32694 = s5 ? tmp32695 : 0;
  assign tmp32691 = s6 ? tmp32692 : tmp32694;
  assign tmp32703 = s3 ? tmp32697 : tmp32667;
  assign tmp32702 = s4 ? tmp32703 : tmp32647;
  assign tmp32701 = s5 ? tmp32702 : 0;
  assign tmp32700 = s6 ? tmp32655 : tmp32701;
  assign tmp32690 = s7 ? tmp32691 : tmp32700;
  assign tmp32689 = s8 ? tmp32690 : tmp32700;
  assign tmp32687 = s9 ? tmp32688 : tmp32689;
  assign tmp32673 = s10 ? tmp32674 : tmp32687;
  assign tmp32707 = s7 ? tmp32677 : tmp32683;
  assign tmp32706 = s8 ? tmp32707 : tmp32683;
  assign tmp32705 = s9 ? tmp32688 : tmp32706;
  assign tmp32704 = s10 ? tmp32674 : tmp32705;
  assign tmp32672 = s11 ? tmp32673 : tmp32704;
  assign tmp32713 = s6 ? tmp32678 : tmp32661;
  assign tmp32712 = s7 ? tmp32554 : tmp32713;
  assign tmp32711 = s8 ? tmp32712 : tmp32553;
  assign tmp32710 = s9 ? tmp32711 : tmp32553;
  assign tmp32717 = s6 ? tmp32692 : tmp32661;
  assign tmp32716 = s7 ? tmp32717 : tmp32654;
  assign tmp32715 = s8 ? tmp32716 : tmp32654;
  assign tmp32714 = s9 ? tmp32670 : tmp32715;
  assign tmp32709 = s10 ? tmp32710 : tmp32714;
  assign tmp32721 = s7 ? tmp32713 : tmp32654;
  assign tmp32720 = s8 ? tmp32721 : tmp32654;
  assign tmp32719 = s9 ? tmp32670 : tmp32720;
  assign tmp32718 = s10 ? tmp32710 : tmp32719;
  assign tmp32708 = s11 ? tmp32709 : tmp32718;
  assign tmp32671 = s12 ? tmp32672 : tmp32708;
  assign tmp32551 = s13 ? tmp32552 : tmp32671;
  assign tmp32732 = s3 ? tmp32664 : tmp32635;
  assign tmp32731 = s4 ? tmp32732 : tmp32647;
  assign tmp32730 = s5 ? tmp32731 : 0;
  assign tmp32729 = s6 ? tmp32655 : tmp32730;
  assign tmp32728 = s7 ? tmp32554 : tmp32729;
  assign tmp32727 = s8 ? tmp32728 : tmp32553;
  assign tmp32726 = s9 ? tmp32727 : tmp32553;
  assign tmp32739 = s3 ? tmp32664 : tmp32698;
  assign tmp32738 = s4 ? tmp32739 : tmp32647;
  assign tmp32737 = s5 ? tmp32738 : 0;
  assign tmp32736 = s6 ? tmp32655 : tmp32737;
  assign tmp32735 = s7 ? tmp32736 : tmp32654;
  assign tmp32734 = s8 ? tmp32735 : tmp32654;
  assign tmp32733 = s9 ? tmp32670 : tmp32734;
  assign tmp32725 = s10 ? tmp32726 : tmp32733;
  assign tmp32743 = s7 ? tmp32729 : tmp32654;
  assign tmp32742 = s8 ? tmp32743 : tmp32654;
  assign tmp32741 = s9 ? tmp32670 : tmp32742;
  assign tmp32740 = s10 ? tmp32726 : tmp32741;
  assign tmp32724 = s11 ? tmp32725 : tmp32740;
  assign tmp32723 = s12 ? tmp32724 : tmp32552;
  assign tmp32722 = s13 ? tmp32723 : tmp32552;
  assign tmp32550 = s14 ? tmp32551 : tmp32722;
  assign tmp32549 = s15 ? tmp32550 : tmp32552;
  assign tmp32751 = s8 ? tmp32712 : tmp32554;
  assign tmp32750 = s9 ? tmp32751 : tmp32717;
  assign tmp32749 = s10 ? tmp32712 : tmp32750;
  assign tmp32753 = s9 ? tmp32751 : tmp32713;
  assign tmp32752 = s10 ? tmp32712 : tmp32753;
  assign tmp32748 = s11 ? tmp32749 : tmp32752;
  assign tmp32747 = s12 ? tmp32672 : tmp32748;
  assign tmp32746 = s13 ? tmp32552 : tmp32747;
  assign tmp32759 = s8 ? tmp32728 : tmp32554;
  assign tmp32758 = s9 ? tmp32759 : tmp32736;
  assign tmp32757 = s10 ? tmp32728 : tmp32758;
  assign tmp32761 = s9 ? tmp32759 : tmp32729;
  assign tmp32760 = s10 ? tmp32728 : tmp32761;
  assign tmp32756 = s11 ? tmp32757 : tmp32760;
  assign tmp32755 = s12 ? tmp32756 : tmp32552;
  assign tmp32754 = s13 ? tmp32755 : tmp32552;
  assign tmp32745 = s14 ? tmp32746 : tmp32754;
  assign tmp32744 = s15 ? tmp32745 : tmp32552;
  assign tmp32548 = s16 ? tmp32549 : tmp32744;
  assign tmp32769 = s9 ? tmp32712 : tmp32711;
  assign tmp32770 = s9 ? tmp32670 : tmp32716;
  assign tmp32768 = s10 ? tmp32769 : tmp32770;
  assign tmp32772 = s9 ? tmp32670 : tmp32721;
  assign tmp32771 = s10 ? tmp32769 : tmp32772;
  assign tmp32767 = s11 ? tmp32768 : tmp32771;
  assign tmp32766 = s12 ? tmp32672 : tmp32767;
  assign tmp32765 = s13 ? tmp32552 : tmp32766;
  assign tmp32777 = s9 ? tmp32728 : tmp32727;
  assign tmp32778 = s9 ? tmp32670 : tmp32735;
  assign tmp32776 = s10 ? tmp32777 : tmp32778;
  assign tmp32780 = s9 ? tmp32670 : tmp32743;
  assign tmp32779 = s10 ? tmp32777 : tmp32780;
  assign tmp32775 = s11 ? tmp32776 : tmp32779;
  assign tmp32774 = s12 ? tmp32775 : tmp32552;
  assign tmp32773 = s13 ? tmp32774 : tmp32552;
  assign tmp32764 = s14 ? tmp32765 : tmp32773;
  assign tmp32763 = s15 ? tmp32764 : tmp32552;
  assign tmp32762 = s16 ? tmp32763 : tmp32744;
  assign tmp32547 = s17 ? tmp32548 : tmp32762;
  assign s6n = tmp32547;

  assign tmp32797 = ~(l4 ? 1 : 0);
  assign tmp32796 = l3 ? 1 : tmp32797;
  assign tmp32799 = l4 ? 1 : 0;
  assign tmp32798 = ~(l3 ? tmp32799 : 0);
  assign tmp32795 = l2 ? tmp32796 : tmp32798;
  assign tmp32800 = l2 ? tmp32796 : 1;
  assign tmp32794 = l1 ? tmp32795 : tmp32800;
  assign tmp32805 = ~(l2 ? tmp32799 : 0);
  assign tmp32804 = l1 ? tmp32795 : tmp32805;
  assign tmp32808 = l3 ? 1 : tmp32799;
  assign tmp32807 = ~(l2 ? tmp32808 : 0);
  assign tmp32806 = l1 ? tmp32795 : tmp32807;
  assign tmp32803 = s0 ? tmp32804 : tmp32806;
  assign tmp32809 = s0 ? tmp32794 : tmp32806;
  assign tmp32802 = s1 ? tmp32803 : tmp32809;
  assign tmp32811 = s0 ? tmp32794 : tmp32804;
  assign tmp32812 = s0 ? tmp32806 : tmp32794;
  assign tmp32810 = s1 ? tmp32811 : tmp32812;
  assign tmp32801 = s2 ? tmp32802 : tmp32810;
  assign tmp32793 = s3 ? tmp32794 : tmp32801;
  assign tmp32819 = l3 ? tmp32799 : 0;
  assign tmp32818 = ~(l2 ? tmp32819 : 0);
  assign tmp32817 = l1 ? tmp32795 : tmp32818;
  assign tmp32816 = s0 ? tmp32794 : tmp32817;
  assign tmp32815 = s1 ? tmp32816 : tmp32809;
  assign tmp32822 = l1 ? tmp32795 : 1;
  assign tmp32821 = s0 ? tmp32794 : tmp32822;
  assign tmp32823 = s0 ? tmp32804 : tmp32822;
  assign tmp32820 = s1 ? tmp32821 : tmp32823;
  assign tmp32814 = s2 ? tmp32815 : tmp32820;
  assign tmp32829 = l3 ? tmp32799 : 1;
  assign tmp32828 = l2 ? tmp32829 : tmp32799;
  assign tmp32830 = l2 ? tmp32808 : tmp32799;
  assign tmp32827 = ~(l1 ? tmp32828 : tmp32830);
  assign tmp32826 = s0 ? tmp32822 : tmp32827;
  assign tmp32825 = s1 ? tmp32804 : tmp32826;
  assign tmp32833 = l1 ? tmp32800 : tmp32807;
  assign tmp32832 = s0 ? tmp32806 : tmp32833;
  assign tmp32835 = l1 ? tmp32799 : tmp32830;
  assign tmp32836 = ~(l1 ? tmp32795 : tmp32807);
  assign tmp32834 = ~(s0 ? tmp32835 : tmp32836);
  assign tmp32831 = s1 ? tmp32832 : tmp32834;
  assign tmp32824 = s2 ? tmp32825 : tmp32831;
  assign tmp32813 = s3 ? tmp32814 : tmp32824;
  assign tmp32792 = s4 ? tmp32793 : tmp32813;
  assign tmp32844 = l2 ? 1 : tmp32798;
  assign tmp32843 = l1 ? tmp32844 : tmp32818;
  assign tmp32842 = s0 ? tmp32794 : tmp32843;
  assign tmp32845 = s0 ? tmp32843 : tmp32804;
  assign tmp32841 = s1 ? tmp32842 : tmp32845;
  assign tmp32848 = l1 ? tmp32800 : tmp32805;
  assign tmp32847 = s0 ? tmp32833 : tmp32848;
  assign tmp32846 = s1 ? tmp32845 : tmp32847;
  assign tmp32840 = s2 ? tmp32841 : tmp32846;
  assign tmp32851 = s0 ? tmp32848 : tmp32800;
  assign tmp32854 = l2 ? tmp32799 : tmp32819;
  assign tmp32855 = l2 ? tmp32808 : tmp32819;
  assign tmp32853 = ~(l1 ? tmp32854 : tmp32855);
  assign tmp32852 = s0 ? tmp32848 : tmp32853;
  assign tmp32850 = s1 ? tmp32851 : tmp32852;
  assign tmp32859 = l2 ? tmp32829 : 1;
  assign tmp32858 = ~(l1 ? 1 : tmp32859);
  assign tmp32857 = s0 ? tmp32835 : tmp32858;
  assign tmp32863 = l3 ? tmp32799 : tmp32797;
  assign tmp32862 = l2 ? tmp32863 : 1;
  assign tmp32861 = l1 ? tmp32800 : tmp32862;
  assign tmp32860 = ~(s0 ? tmp32806 : tmp32861);
  assign tmp32856 = ~(s1 ? tmp32857 : tmp32860);
  assign tmp32849 = s2 ? tmp32850 : tmp32856;
  assign tmp32839 = s3 ? tmp32840 : tmp32849;
  assign tmp32868 = l1 ? 1 : tmp32859;
  assign tmp32867 = s0 ? tmp32868 : tmp32804;
  assign tmp32871 = l2 ? 1 : tmp32796;
  assign tmp32870 = l1 ? tmp32871 : 1;
  assign tmp32873 = l2 ? tmp32808 : 1;
  assign tmp32872 = l1 ? tmp32871 : tmp32873;
  assign tmp32869 = ~(s0 ? tmp32870 : tmp32872);
  assign tmp32866 = s1 ? tmp32867 : tmp32869;
  assign tmp32875 = s0 ? tmp32870 : tmp32872;
  assign tmp32878 = l2 ? tmp32808 : tmp32796;
  assign tmp32880 = l3 ? 1 : 0;
  assign tmp32879 = l2 ? tmp32808 : tmp32880;
  assign tmp32877 = l1 ? tmp32878 : tmp32879;
  assign tmp32876 = s0 ? tmp32877 : tmp32870;
  assign tmp32874 = ~(s1 ? tmp32875 : tmp32876);
  assign tmp32865 = s2 ? tmp32866 : tmp32874;
  assign tmp32885 = l2 ? tmp32799 : tmp32863;
  assign tmp32884 = l1 ? tmp32885 : tmp32855;
  assign tmp32883 = s0 ? tmp32877 : tmp32884;
  assign tmp32887 = l1 ? tmp32854 : tmp32855;
  assign tmp32886 = s0 ? tmp32872 : tmp32887;
  assign tmp32882 = s1 ? tmp32883 : tmp32886;
  assign tmp32890 = l2 ? 1 : tmp32829;
  assign tmp32889 = l1 ? tmp32859 : tmp32890;
  assign tmp32892 = l1 ? tmp32828 : tmp32830;
  assign tmp32891 = s0 ? tmp32892 : tmp32889;
  assign tmp32888 = s1 ? tmp32889 : tmp32891;
  assign tmp32881 = ~(s2 ? tmp32882 : tmp32888);
  assign tmp32864 = s3 ? tmp32865 : tmp32881;
  assign tmp32838 = s4 ? tmp32839 : tmp32864;
  assign tmp32898 = l1 ? tmp32829 : 1;
  assign tmp32897 = s0 ? tmp32887 : tmp32898;
  assign tmp32901 = l2 ? tmp32808 : tmp32829;
  assign tmp32900 = l1 ? tmp32901 : tmp32873;
  assign tmp32899 = s0 ? tmp32898 : tmp32900;
  assign tmp32896 = s1 ? tmp32897 : tmp32899;
  assign tmp32904 = l1 ? tmp32878 : tmp32871;
  assign tmp32903 = s0 ? tmp32900 : tmp32904;
  assign tmp32902 = s1 ? tmp32903 : tmp32904;
  assign tmp32895 = s2 ? tmp32896 : tmp32902;
  assign tmp32907 = s0 ? tmp32904 : 0;
  assign tmp32910 = l2 ? 1 : tmp32799;
  assign tmp32909 = ~(l1 ? tmp32910 : tmp32890);
  assign tmp32908 = ~(s0 ? 1 : tmp32909);
  assign tmp32906 = s1 ? tmp32907 : tmp32908;
  assign tmp32913 = l1 ? tmp32910 : tmp32890;
  assign tmp32912 = s0 ? tmp32913 : 0;
  assign tmp32911 = s1 ? tmp32912 : 0;
  assign tmp32905 = s2 ? tmp32906 : tmp32911;
  assign tmp32894 = s3 ? tmp32895 : tmp32905;
  assign tmp32918 = ~(l1 ? tmp32799 : tmp32830);
  assign tmp32917 = s0 ? 1 : tmp32918;
  assign tmp32916 = s1 ? 1 : tmp32917;
  assign tmp32921 = l1 ? tmp32855 : tmp32879;
  assign tmp32920 = s0 ? tmp32898 : tmp32921;
  assign tmp32919 = ~(s1 ? tmp32920 : tmp32904);
  assign tmp32915 = s2 ? tmp32916 : tmp32919;
  assign tmp32925 = l1 ? tmp32830 : tmp32910;
  assign tmp32924 = s0 ? tmp32900 : tmp32925;
  assign tmp32923 = s1 ? tmp32924 : tmp32912;
  assign tmp32922 = ~(s2 ? tmp32923 : 0);
  assign tmp32914 = ~(s3 ? tmp32915 : tmp32922);
  assign tmp32893 = ~(s4 ? tmp32894 : tmp32914);
  assign tmp32837 = s5 ? tmp32838 : tmp32893;
  assign tmp32791 = s6 ? tmp32792 : tmp32837;
  assign tmp32930 = s1 ? tmp32821 : tmp32804;
  assign tmp32929 = s2 ? tmp32815 : tmp32930;
  assign tmp32932 = s1 ? tmp32794 : tmp32827;
  assign tmp32931 = s2 ? tmp32932 : tmp32831;
  assign tmp32928 = s3 ? tmp32929 : tmp32931;
  assign tmp32927 = s4 ? tmp32793 : tmp32928;
  assign tmp32937 = s1 ? tmp32842 : tmp32804;
  assign tmp32938 = s1 ? tmp32804 : tmp32847;
  assign tmp32936 = s2 ? tmp32937 : tmp32938;
  assign tmp32940 = s1 ? tmp32800 : tmp32853;
  assign tmp32939 = s2 ? tmp32940 : tmp32856;
  assign tmp32935 = s3 ? tmp32936 : tmp32939;
  assign tmp32943 = ~(s1 ? tmp32870 : tmp32876);
  assign tmp32942 = s2 ? tmp32866 : tmp32943;
  assign tmp32945 = s1 ? tmp32883 : tmp32887;
  assign tmp32946 = s1 ? tmp32889 : tmp32892;
  assign tmp32944 = ~(s2 ? tmp32945 : tmp32946);
  assign tmp32941 = s3 ? tmp32942 : tmp32944;
  assign tmp32934 = s4 ? tmp32935 : tmp32941;
  assign tmp32950 = s1 ? tmp32897 : tmp32900;
  assign tmp32949 = s2 ? tmp32950 : tmp32904;
  assign tmp32952 = s1 ? 1 : tmp32909;
  assign tmp32951 = ~(s2 ? tmp32952 : 1);
  assign tmp32948 = s3 ? tmp32949 : tmp32951;
  assign tmp32955 = s1 ? 1 : tmp32918;
  assign tmp32956 = ~(l1 ? tmp32855 : tmp32879);
  assign tmp32954 = s2 ? tmp32955 : tmp32956;
  assign tmp32957 = ~(s1 ? tmp32925 : 0);
  assign tmp32953 = ~(s3 ? tmp32954 : tmp32957);
  assign tmp32947 = ~(s4 ? tmp32948 : tmp32953);
  assign tmp32933 = s5 ? tmp32934 : tmp32947;
  assign tmp32926 = s6 ? tmp32927 : tmp32933;
  assign tmp32790 = s7 ? tmp32791 : tmp32926;
  assign tmp32964 = ~(l1 ? tmp32878 : tmp32879);
  assign tmp32963 = s2 ? tmp32866 : tmp32964;
  assign tmp32962 = s3 ? tmp32963 : tmp32944;
  assign tmp32961 = s4 ? tmp32935 : tmp32962;
  assign tmp32960 = s5 ? tmp32961 : tmp32947;
  assign tmp32959 = s6 ? tmp32927 : tmp32960;
  assign tmp32958 = s7 ? tmp32791 : tmp32959;
  assign tmp32789 = s8 ? tmp32790 : tmp32958;
  assign tmp32788 = s9 ? tmp32789 : tmp32958;
  assign tmp32966 = s8 ? tmp32958 : tmp32791;
  assign tmp32974 = ~(s1 ? tmp32870 : tmp32877);
  assign tmp32973 = s2 ? tmp32866 : tmp32974;
  assign tmp32972 = s3 ? tmp32973 : tmp32944;
  assign tmp32971 = s4 ? tmp32935 : tmp32972;
  assign tmp32970 = s5 ? tmp32971 : tmp32947;
  assign tmp32969 = s6 ? tmp32927 : tmp32970;
  assign tmp32968 = s7 ? tmp32969 : tmp32959;
  assign tmp32967 = s8 ? tmp32968 : tmp32959;
  assign tmp32965 = s9 ? tmp32966 : tmp32967;
  assign tmp32787 = s10 ? tmp32788 : tmp32965;
  assign tmp32978 = s7 ? tmp32926 : tmp32959;
  assign tmp32977 = s8 ? tmp32978 : tmp32959;
  assign tmp32976 = s9 ? tmp32966 : tmp32977;
  assign tmp32975 = s10 ? tmp32788 : tmp32976;
  assign tmp32786 = s11 ? tmp32787 : tmp32975;
  assign tmp32989 = s1 ? tmp32794 : tmp32826;
  assign tmp32988 = s2 ? tmp32989 : tmp32831;
  assign tmp32987 = s3 ? tmp32814 : tmp32988;
  assign tmp32986 = s4 ? tmp32793 : tmp32987;
  assign tmp32991 = s4 ? tmp32839 : tmp32962;
  assign tmp32990 = s5 ? tmp32991 : tmp32947;
  assign tmp32985 = s6 ? tmp32986 : tmp32990;
  assign tmp32984 = s7 ? tmp32791 : tmp32985;
  assign tmp32996 = s3 ? tmp32840 : tmp32939;
  assign tmp32995 = s4 ? tmp32996 : tmp32962;
  assign tmp32994 = s5 ? tmp32995 : tmp32947;
  assign tmp32993 = s6 ? tmp32927 : tmp32994;
  assign tmp32992 = s7 ? tmp32791 : tmp32993;
  assign tmp32983 = s8 ? tmp32984 : tmp32992;
  assign tmp32982 = s9 ? tmp32983 : tmp32992;
  assign tmp32998 = s8 ? tmp32992 : tmp32791;
  assign tmp33003 = s3 ? tmp32814 : tmp32931;
  assign tmp33002 = s4 ? tmp32793 : tmp33003;
  assign tmp33007 = s2 ? tmp32841 : tmp32938;
  assign tmp33009 = s1 ? tmp32851 : tmp32853;
  assign tmp33008 = s2 ? tmp33009 : tmp32856;
  assign tmp33006 = s3 ? tmp33007 : tmp33008;
  assign tmp33005 = s4 ? tmp33006 : tmp32962;
  assign tmp33004 = s5 ? tmp33005 : tmp32947;
  assign tmp33001 = s6 ? tmp33002 : tmp33004;
  assign tmp33013 = s3 ? tmp33007 : tmp32939;
  assign tmp33012 = s4 ? tmp33013 : tmp32962;
  assign tmp33011 = s5 ? tmp33012 : tmp32947;
  assign tmp33010 = s6 ? tmp32927 : tmp33011;
  assign tmp33000 = s7 ? tmp33001 : tmp33010;
  assign tmp32999 = s8 ? tmp33000 : tmp33010;
  assign tmp32997 = s9 ? tmp32998 : tmp32999;
  assign tmp32981 = s10 ? tmp32982 : tmp32997;
  assign tmp33017 = s7 ? tmp32985 : tmp32993;
  assign tmp33016 = s8 ? tmp33017 : tmp32993;
  assign tmp33015 = s9 ? tmp32998 : tmp33016;
  assign tmp33014 = s10 ? tmp32982 : tmp33015;
  assign tmp32980 = s11 ? tmp32981 : tmp33014;
  assign tmp33023 = s6 ? tmp32986 : tmp32960;
  assign tmp33022 = s7 ? tmp32791 : tmp33023;
  assign tmp33021 = s8 ? tmp33022 : tmp32958;
  assign tmp33020 = s9 ? tmp33021 : tmp32958;
  assign tmp33027 = s6 ? tmp33002 : tmp32960;
  assign tmp33026 = s7 ? tmp33027 : tmp32959;
  assign tmp33025 = s8 ? tmp33026 : tmp32959;
  assign tmp33024 = s9 ? tmp32966 : tmp33025;
  assign tmp33019 = s10 ? tmp33020 : tmp33024;
  assign tmp33031 = s7 ? tmp33023 : tmp32959;
  assign tmp33030 = s8 ? tmp33031 : tmp32959;
  assign tmp33029 = s9 ? tmp32966 : tmp33030;
  assign tmp33028 = s10 ? tmp33020 : tmp33029;
  assign tmp33018 = s11 ? tmp33019 : tmp33028;
  assign tmp32979 = s12 ? tmp32980 : tmp33018;
  assign tmp32785 = s13 ? tmp32786 : tmp32979;
  assign tmp33042 = s3 ? tmp32936 : tmp32849;
  assign tmp33041 = s4 ? tmp33042 : tmp32962;
  assign tmp33040 = s5 ? tmp33041 : tmp32947;
  assign tmp33039 = s6 ? tmp32927 : tmp33040;
  assign tmp33038 = s7 ? tmp32791 : tmp33039;
  assign tmp33037 = s8 ? tmp33038 : tmp32958;
  assign tmp33036 = s9 ? tmp33037 : tmp32958;
  assign tmp33049 = s3 ? tmp32936 : tmp33008;
  assign tmp33048 = s4 ? tmp33049 : tmp32962;
  assign tmp33047 = s5 ? tmp33048 : tmp32947;
  assign tmp33046 = s6 ? tmp32927 : tmp33047;
  assign tmp33045 = s7 ? tmp33046 : tmp32959;
  assign tmp33044 = s8 ? tmp33045 : tmp32959;
  assign tmp33043 = s9 ? tmp32966 : tmp33044;
  assign tmp33035 = s10 ? tmp33036 : tmp33043;
  assign tmp33053 = s7 ? tmp33039 : tmp32959;
  assign tmp33052 = s8 ? tmp33053 : tmp32959;
  assign tmp33051 = s9 ? tmp32966 : tmp33052;
  assign tmp33050 = s10 ? tmp33036 : tmp33051;
  assign tmp33034 = s11 ? tmp33035 : tmp33050;
  assign tmp33064 = ~(s1 ? tmp32872 : tmp32877);
  assign tmp33063 = s2 ? tmp32866 : tmp33064;
  assign tmp33065 = ~(s2 ? tmp32882 : tmp32946);
  assign tmp33062 = s3 ? tmp33063 : tmp33065;
  assign tmp33061 = s4 ? tmp32935 : tmp33062;
  assign tmp33060 = s5 ? tmp33061 : tmp32947;
  assign tmp33059 = s6 ? tmp32927 : tmp33060;
  assign tmp33058 = s7 ? tmp32791 : tmp33059;
  assign tmp33057 = s8 ? tmp33058 : tmp32958;
  assign tmp33056 = s9 ? tmp33057 : tmp32958;
  assign tmp33072 = s3 ? tmp33063 : tmp32944;
  assign tmp33071 = s4 ? tmp32935 : tmp33072;
  assign tmp33070 = s5 ? tmp33071 : tmp32947;
  assign tmp33069 = s6 ? tmp32927 : tmp33070;
  assign tmp33068 = s7 ? tmp33069 : tmp32959;
  assign tmp33067 = s8 ? tmp33068 : tmp32959;
  assign tmp33066 = s9 ? tmp32966 : tmp33067;
  assign tmp33055 = s10 ? tmp33056 : tmp33066;
  assign tmp33076 = s7 ? tmp33059 : tmp32959;
  assign tmp33075 = s8 ? tmp33076 : tmp32959;
  assign tmp33074 = s9 ? tmp32966 : tmp33075;
  assign tmp33073 = s10 ? tmp33056 : tmp33074;
  assign tmp33054 = s11 ? tmp33055 : tmp33073;
  assign tmp33033 = s12 ? tmp33034 : tmp33054;
  assign tmp33085 = s1 ? tmp32907 : tmp32913;
  assign tmp33084 = s2 ? tmp33085 : 0;
  assign tmp33083 = s3 ? tmp32949 : tmp33084;
  assign tmp33088 = ~(s1 ? tmp32921 : tmp32904);
  assign tmp33087 = s2 ? tmp32955 : tmp33088;
  assign tmp33086 = ~(s3 ? tmp33087 : tmp32957);
  assign tmp33082 = ~(s4 ? tmp33083 : tmp33086);
  assign tmp33081 = s5 ? tmp32961 : tmp33082;
  assign tmp33080 = s6 ? tmp32927 : tmp33081;
  assign tmp33079 = s7 ? tmp32791 : tmp33080;
  assign tmp33090 = s8 ? tmp33079 : tmp32791;
  assign tmp33093 = ~(s4 ? tmp33083 : tmp32953);
  assign tmp33092 = s5 ? tmp32961 : tmp33093;
  assign tmp33091 = s6 ? tmp32927 : tmp33092;
  assign tmp33089 = s9 ? tmp33090 : tmp33091;
  assign tmp33078 = s10 ? tmp33079 : tmp33089;
  assign tmp33095 = s9 ? tmp33090 : tmp33080;
  assign tmp33094 = s10 ? tmp33079 : tmp33095;
  assign tmp33077 = s11 ? tmp33078 : tmp33094;
  assign tmp33032 = s13 ? tmp33033 : tmp33077;
  assign tmp32784 = s14 ? tmp32785 : tmp33032;
  assign tmp33106 = s2 ? tmp32896 : tmp32904;
  assign tmp33105 = s3 ? tmp33106 : tmp32951;
  assign tmp33109 = ~(s0 ? tmp32898 : tmp32921);
  assign tmp33108 = s2 ? tmp32955 : tmp33109;
  assign tmp33107 = ~(s3 ? tmp33108 : tmp32957);
  assign tmp33104 = ~(s4 ? tmp33105 : tmp33107);
  assign tmp33103 = s5 ? tmp32961 : tmp33104;
  assign tmp33102 = s6 ? tmp32927 : tmp33103;
  assign tmp33101 = s7 ? tmp32791 : tmp33102;
  assign tmp33111 = s8 ? tmp33101 : tmp32791;
  assign tmp33114 = ~(s4 ? tmp33105 : tmp32953);
  assign tmp33113 = s5 ? tmp32961 : tmp33114;
  assign tmp33112 = s6 ? tmp32927 : tmp33113;
  assign tmp33110 = s9 ? tmp33111 : tmp33112;
  assign tmp33100 = s10 ? tmp33101 : tmp33110;
  assign tmp33116 = s9 ? tmp33111 : tmp33102;
  assign tmp33115 = s10 ? tmp33101 : tmp33116;
  assign tmp33099 = s11 ? tmp33100 : tmp33115;
  assign tmp33124 = ~(s2 ? tmp32945 : tmp32888);
  assign tmp33123 = s3 ? tmp32963 : tmp33124;
  assign tmp33122 = s4 ? tmp32935 : tmp33123;
  assign tmp33121 = s5 ? tmp33122 : tmp32947;
  assign tmp33120 = s6 ? tmp32927 : tmp33121;
  assign tmp33119 = s7 ? tmp32791 : tmp33120;
  assign tmp33126 = s8 ? tmp33119 : tmp32791;
  assign tmp33125 = s9 ? tmp33126 : tmp32959;
  assign tmp33118 = s10 ? tmp33119 : tmp33125;
  assign tmp33128 = s9 ? tmp33126 : tmp33120;
  assign tmp33127 = s10 ? tmp33119 : tmp33128;
  assign tmp33117 = s11 ? tmp33118 : tmp33127;
  assign tmp33098 = s12 ? tmp33099 : tmp33117;
  assign tmp33137 = s1 ? tmp32925 : 0;
  assign tmp33136 = ~(s2 ? tmp33137 : 0);
  assign tmp33135 = ~(s3 ? tmp32954 : tmp33136);
  assign tmp33134 = ~(s4 ? tmp32948 : tmp33135);
  assign tmp33133 = s5 ? tmp32961 : tmp33134;
  assign tmp33132 = s6 ? tmp32927 : tmp33133;
  assign tmp33131 = s7 ? tmp32791 : tmp33132;
  assign tmp33139 = s8 ? tmp33131 : tmp32791;
  assign tmp33138 = s9 ? tmp33139 : tmp33132;
  assign tmp33130 = s10 ? tmp33131 : tmp33138;
  assign tmp33148 = ~(s1 ? tmp32912 : 0);
  assign tmp33147 = ~(s2 ? tmp32952 : tmp33148);
  assign tmp33146 = s3 ? tmp32949 : tmp33147;
  assign tmp33150 = ~(s1 ? tmp32925 : tmp32912);
  assign tmp33149 = ~(s3 ? tmp32954 : tmp33150);
  assign tmp33145 = ~(s4 ? tmp33146 : tmp33149);
  assign tmp33144 = s5 ? tmp32961 : tmp33145;
  assign tmp33143 = s6 ? tmp32927 : tmp33144;
  assign tmp33142 = s7 ? tmp32791 : tmp33143;
  assign tmp33152 = s8 ? tmp33142 : tmp32791;
  assign tmp33155 = ~(s4 ? tmp33146 : tmp32953);
  assign tmp33154 = s5 ? tmp32961 : tmp33155;
  assign tmp33153 = s6 ? tmp32927 : tmp33154;
  assign tmp33151 = s9 ? tmp33152 : tmp33153;
  assign tmp33141 = s10 ? tmp33142 : tmp33151;
  assign tmp33157 = s9 ? tmp33152 : tmp33143;
  assign tmp33156 = s10 ? tmp33142 : tmp33157;
  assign tmp33140 = s11 ? tmp33141 : tmp33156;
  assign tmp33129 = s12 ? tmp33130 : tmp33140;
  assign tmp33097 = s13 ? tmp33098 : tmp33129;
  assign tmp33168 = ~(s3 ? tmp33087 : tmp33136);
  assign tmp33167 = ~(s4 ? tmp33083 : tmp33168);
  assign tmp33166 = s5 ? tmp33061 : tmp33167;
  assign tmp33165 = s6 ? tmp32927 : tmp33166;
  assign tmp33164 = s7 ? tmp32791 : tmp33165;
  assign tmp33171 = s5 ? tmp32961 : tmp33167;
  assign tmp33170 = s6 ? tmp32927 : tmp33171;
  assign tmp33169 = s7 ? tmp32791 : tmp33170;
  assign tmp33163 = s8 ? tmp33164 : tmp33169;
  assign tmp33162 = s9 ? tmp33163 : tmp33169;
  assign tmp33173 = s8 ? tmp33169 : tmp32791;
  assign tmp33177 = s5 ? tmp33071 : tmp33093;
  assign tmp33176 = s6 ? tmp32927 : tmp33177;
  assign tmp33175 = s7 ? tmp33176 : tmp33091;
  assign tmp33174 = s8 ? tmp33175 : tmp33091;
  assign tmp33172 = s9 ? tmp33173 : tmp33174;
  assign tmp33161 = s10 ? tmp33162 : tmp33172;
  assign tmp33181 = s7 ? tmp33165 : tmp33170;
  assign tmp33180 = s8 ? tmp33181 : tmp33170;
  assign tmp33179 = s9 ? tmp33173 : tmp33180;
  assign tmp33178 = s10 ? tmp33162 : tmp33179;
  assign tmp33160 = s11 ? tmp33161 : tmp33178;
  assign tmp33191 = s2 ? tmp32950 : tmp32902;
  assign tmp33190 = s3 ? tmp33191 : tmp32951;
  assign tmp33193 = ~(s1 ? tmp32924 : 0);
  assign tmp33192 = ~(s3 ? tmp32954 : tmp33193);
  assign tmp33189 = ~(s4 ? tmp33190 : tmp33192);
  assign tmp33188 = s5 ? tmp32961 : tmp33189;
  assign tmp33187 = s6 ? tmp32927 : tmp33188;
  assign tmp33186 = s7 ? tmp32791 : tmp33187;
  assign tmp33185 = s8 ? tmp33186 : tmp32958;
  assign tmp33184 = s9 ? tmp33185 : tmp32958;
  assign tmp33199 = ~(s4 ? tmp33190 : tmp32953);
  assign tmp33198 = s5 ? tmp32961 : tmp33199;
  assign tmp33197 = s6 ? tmp32927 : tmp33198;
  assign tmp33196 = s7 ? tmp33197 : tmp32959;
  assign tmp33195 = s8 ? tmp33196 : tmp32959;
  assign tmp33194 = s9 ? tmp32966 : tmp33195;
  assign tmp33183 = s10 ? tmp33184 : tmp33194;
  assign tmp33203 = s7 ? tmp33187 : tmp32959;
  assign tmp33202 = s8 ? tmp33203 : tmp32959;
  assign tmp33201 = s9 ? tmp32966 : tmp33202;
  assign tmp33200 = s10 ? tmp33184 : tmp33201;
  assign tmp33182 = s11 ? tmp33183 : tmp33200;
  assign tmp33159 = s12 ? tmp33160 : tmp33182;
  assign tmp33212 = s0 ? 1 : tmp32909;
  assign tmp33211 = s1 ? 1 : tmp33212;
  assign tmp33210 = ~(s2 ? tmp33211 : 1);
  assign tmp33209 = s3 ? tmp32949 : tmp33210;
  assign tmp33214 = s2 ? tmp32916 : tmp32956;
  assign tmp33213 = ~(s3 ? tmp33214 : tmp33136);
  assign tmp33208 = ~(s4 ? tmp33209 : tmp33213);
  assign tmp33207 = s5 ? tmp32961 : tmp33208;
  assign tmp33206 = s6 ? tmp32927 : tmp33207;
  assign tmp33205 = s7 ? tmp32791 : tmp33206;
  assign tmp33216 = s8 ? tmp33205 : tmp32791;
  assign tmp33215 = s9 ? tmp33216 : tmp33206;
  assign tmp33204 = s10 ? tmp33205 : tmp33215;
  assign tmp33158 = s13 ? tmp33159 : tmp33204;
  assign tmp33096 = s14 ? tmp33097 : tmp33158;
  assign tmp32783 = s15 ? tmp32784 : tmp33096;
  assign tmp33223 = s8 ? tmp32790 : tmp32791;
  assign tmp33222 = s9 ? tmp33223 : tmp32969;
  assign tmp33221 = s10 ? tmp32790 : tmp33222;
  assign tmp33225 = s9 ? tmp33223 : tmp32926;
  assign tmp33224 = s10 ? tmp32790 : tmp33225;
  assign tmp33220 = s11 ? tmp33221 : tmp33224;
  assign tmp33230 = s8 ? tmp33022 : tmp32791;
  assign tmp33229 = s9 ? tmp33230 : tmp33027;
  assign tmp33228 = s10 ? tmp33022 : tmp33229;
  assign tmp33232 = s9 ? tmp33230 : tmp33023;
  assign tmp33231 = s10 ? tmp33022 : tmp33232;
  assign tmp33227 = s11 ? tmp33228 : tmp33231;
  assign tmp33226 = s12 ? tmp32980 : tmp33227;
  assign tmp33219 = s13 ? tmp33220 : tmp33226;
  assign tmp33238 = s8 ? tmp33038 : tmp32791;
  assign tmp33237 = s9 ? tmp33238 : tmp33046;
  assign tmp33236 = s10 ? tmp33038 : tmp33237;
  assign tmp33240 = s9 ? tmp33238 : tmp33039;
  assign tmp33239 = s10 ? tmp33038 : tmp33240;
  assign tmp33235 = s11 ? tmp33236 : tmp33239;
  assign tmp33244 = s8 ? tmp33058 : tmp32791;
  assign tmp33243 = s9 ? tmp33244 : tmp33069;
  assign tmp33242 = s10 ? tmp33058 : tmp33243;
  assign tmp33246 = s9 ? tmp33244 : tmp33059;
  assign tmp33245 = s10 ? tmp33058 : tmp33246;
  assign tmp33241 = s11 ? tmp33242 : tmp33245;
  assign tmp33234 = s12 ? tmp33235 : tmp33241;
  assign tmp33250 = s8 ? tmp32958 : tmp33079;
  assign tmp33249 = s9 ? tmp32958 : tmp33250;
  assign tmp33253 = s7 ? tmp32959 : tmp33091;
  assign tmp33252 = s8 ? tmp33253 : tmp32959;
  assign tmp33251 = s9 ? tmp32966 : tmp33252;
  assign tmp33248 = s10 ? tmp33249 : tmp33251;
  assign tmp33257 = s7 ? tmp32959 : tmp33080;
  assign tmp33256 = s8 ? tmp33257 : tmp32959;
  assign tmp33255 = s9 ? tmp32966 : tmp33256;
  assign tmp33254 = s10 ? tmp33249 : tmp33255;
  assign tmp33247 = s11 ? tmp33248 : tmp33254;
  assign tmp33233 = s13 ? tmp33234 : tmp33247;
  assign tmp33218 = s14 ? tmp33219 : tmp33233;
  assign tmp33264 = s8 ? tmp32958 : tmp33169;
  assign tmp33263 = s9 ? tmp33057 : tmp33264;
  assign tmp33267 = s7 ? tmp33069 : tmp33091;
  assign tmp33266 = s8 ? tmp33267 : tmp32959;
  assign tmp33265 = s9 ? tmp32966 : tmp33266;
  assign tmp33262 = s10 ? tmp33263 : tmp33265;
  assign tmp33271 = s7 ? tmp33059 : tmp33170;
  assign tmp33270 = s8 ? tmp33271 : tmp32959;
  assign tmp33269 = s9 ? tmp32966 : tmp33270;
  assign tmp33268 = s10 ? tmp33263 : tmp33269;
  assign tmp33261 = s11 ? tmp33262 : tmp33268;
  assign tmp33275 = s8 ? tmp33186 : tmp32791;
  assign tmp33274 = s9 ? tmp33275 : tmp33197;
  assign tmp33273 = s10 ? tmp33186 : tmp33274;
  assign tmp33277 = s9 ? tmp33275 : tmp33187;
  assign tmp33276 = s10 ? tmp33186 : tmp33277;
  assign tmp33272 = s11 ? tmp33273 : tmp33276;
  assign tmp33260 = s12 ? tmp33261 : tmp33272;
  assign tmp33259 = s13 ? tmp33260 : tmp33204;
  assign tmp33258 = s14 ? tmp33097 : tmp33259;
  assign tmp33217 = s15 ? tmp33218 : tmp33258;
  assign tmp32782 = s16 ? tmp32783 : tmp33217;
  assign tmp33284 = s9 ? tmp32790 : tmp32789;
  assign tmp33285 = s9 ? tmp32966 : tmp32968;
  assign tmp33283 = s10 ? tmp33284 : tmp33285;
  assign tmp33287 = s9 ? tmp32966 : tmp32978;
  assign tmp33286 = s10 ? tmp33284 : tmp33287;
  assign tmp33282 = s11 ? tmp33283 : tmp33286;
  assign tmp33291 = s9 ? tmp33022 : tmp33021;
  assign tmp33292 = s9 ? tmp32966 : tmp33026;
  assign tmp33290 = s10 ? tmp33291 : tmp33292;
  assign tmp33294 = s9 ? tmp32966 : tmp33031;
  assign tmp33293 = s10 ? tmp33291 : tmp33294;
  assign tmp33289 = s11 ? tmp33290 : tmp33293;
  assign tmp33288 = s12 ? tmp32980 : tmp33289;
  assign tmp33281 = s13 ? tmp33282 : tmp33288;
  assign tmp33299 = s9 ? tmp33038 : tmp33037;
  assign tmp33300 = s9 ? tmp32966 : tmp33045;
  assign tmp33298 = s10 ? tmp33299 : tmp33300;
  assign tmp33302 = s9 ? tmp32966 : tmp33053;
  assign tmp33301 = s10 ? tmp33299 : tmp33302;
  assign tmp33297 = s11 ? tmp33298 : tmp33301;
  assign tmp33305 = s9 ? tmp33058 : tmp33057;
  assign tmp33306 = s9 ? tmp32966 : tmp33068;
  assign tmp33304 = s10 ? tmp33305 : tmp33306;
  assign tmp33308 = s9 ? tmp32966 : tmp33076;
  assign tmp33307 = s10 ? tmp33305 : tmp33308;
  assign tmp33303 = s11 ? tmp33304 : tmp33307;
  assign tmp33296 = s12 ? tmp33297 : tmp33303;
  assign tmp33295 = s13 ? tmp33296 : tmp33077;
  assign tmp33280 = s14 ? tmp33281 : tmp33295;
  assign tmp33314 = s9 ? tmp33186 : tmp33185;
  assign tmp33315 = s9 ? tmp32966 : tmp33196;
  assign tmp33313 = s10 ? tmp33314 : tmp33315;
  assign tmp33317 = s9 ? tmp32966 : tmp33203;
  assign tmp33316 = s10 ? tmp33314 : tmp33317;
  assign tmp33312 = s11 ? tmp33313 : tmp33316;
  assign tmp33311 = s12 ? tmp33160 : tmp33312;
  assign tmp33310 = s13 ? tmp33311 : tmp33204;
  assign tmp33309 = s14 ? tmp33097 : tmp33310;
  assign tmp33279 = s15 ? tmp33280 : tmp33309;
  assign tmp33320 = s13 ? tmp33234 : tmp33077;
  assign tmp33319 = s14 ? tmp33219 : tmp33320;
  assign tmp33323 = s12 ? tmp33160 : tmp33272;
  assign tmp33322 = s13 ? tmp33323 : tmp33204;
  assign tmp33321 = s14 ? tmp33097 : tmp33322;
  assign tmp33318 = s15 ? tmp33319 : tmp33321;
  assign tmp33278 = s16 ? tmp33279 : tmp33318;
  assign tmp32781 = ~(s17 ? tmp32782 : tmp33278);
  assign s5n = tmp32781;

  assign tmp33346 = l4 ? 1 : 0;
  assign tmp33345 = l3 ? 1 : tmp33346;
  assign tmp33344 = l2 ? tmp33345 : 1;
  assign tmp33349 = ~(l4 ? 1 : 0);
  assign tmp33348 = l3 ? tmp33346 : tmp33349;
  assign tmp33347 = ~(l2 ? tmp33346 : tmp33348);
  assign tmp33343 = ~(l1 ? tmp33344 : tmp33347);
  assign tmp33342 = s0 ? 1 : tmp33343;
  assign tmp33353 = l3 ? tmp33346 : 0;
  assign tmp33352 = ~(l2 ? tmp33346 : tmp33353);
  assign tmp33351 = l1 ? 1 : tmp33352;
  assign tmp33354 = l1 ? tmp33344 : tmp33347;
  assign tmp33350 = ~(s0 ? tmp33351 : tmp33354);
  assign tmp33341 = s1 ? tmp33342 : tmp33350;
  assign tmp33340 = s2 ? 1 : tmp33341;
  assign tmp33360 = l3 ? 1 : tmp33349;
  assign tmp33359 = l2 ? tmp33360 : tmp33349;
  assign tmp33361 = l2 ? 1 : tmp33360;
  assign tmp33358 = l1 ? tmp33359 : tmp33361;
  assign tmp33363 = ~(l2 ? tmp33345 : tmp33348);
  assign tmp33362 = ~(l1 ? tmp33344 : tmp33363);
  assign tmp33357 = s0 ? tmp33358 : tmp33362;
  assign tmp33365 = l1 ? tmp33344 : tmp33352;
  assign tmp33366 = l1 ? tmp33344 : tmp33363;
  assign tmp33364 = ~(s0 ? tmp33365 : tmp33366);
  assign tmp33356 = s1 ? tmp33357 : tmp33364;
  assign tmp33368 = s0 ? tmp33365 : tmp33351;
  assign tmp33369 = s0 ? tmp33366 : tmp33354;
  assign tmp33367 = ~(s1 ? tmp33368 : tmp33369);
  assign tmp33355 = s2 ? tmp33356 : tmp33367;
  assign tmp33339 = s3 ? tmp33340 : tmp33355;
  assign tmp33375 = ~(l3 ? tmp33346 : 0);
  assign tmp33374 = l1 ? 1 : tmp33375;
  assign tmp33373 = s0 ? tmp33354 : tmp33374;
  assign tmp33376 = s0 ? tmp33354 : tmp33366;
  assign tmp33372 = s1 ? tmp33373 : tmp33376;
  assign tmp33380 = l2 ? 1 : tmp33375;
  assign tmp33379 = l1 ? 1 : tmp33380;
  assign tmp33378 = s0 ? tmp33354 : tmp33379;
  assign tmp33383 = ~(l2 ? tmp33346 : 0);
  assign tmp33382 = l1 ? 1 : tmp33383;
  assign tmp33381 = s0 ? tmp33382 : tmp33379;
  assign tmp33377 = s1 ? tmp33378 : tmp33381;
  assign tmp33371 = s2 ? tmp33372 : tmp33377;
  assign tmp33389 = l3 ? tmp33346 : 1;
  assign tmp33388 = ~(l2 ? tmp33389 : 0);
  assign tmp33387 = l1 ? tmp33361 : tmp33388;
  assign tmp33386 = s0 ? tmp33387 : tmp33351;
  assign tmp33392 = l2 ? tmp33389 : tmp33345;
  assign tmp33391 = l1 ? 1 : tmp33392;
  assign tmp33390 = s0 ? tmp33379 : tmp33391;
  assign tmp33385 = s1 ? tmp33386 : tmp33390;
  assign tmp33396 = l2 ? tmp33348 : tmp33353;
  assign tmp33397 = l2 ? tmp33345 : tmp33348;
  assign tmp33395 = ~(l1 ? tmp33396 : tmp33397);
  assign tmp33394 = s0 ? tmp33366 : tmp33395;
  assign tmp33400 = l2 ? tmp33348 : tmp33345;
  assign tmp33399 = l1 ? tmp33344 : tmp33400;
  assign tmp33398 = s0 ? tmp33399 : tmp33366;
  assign tmp33393 = s1 ? tmp33394 : tmp33398;
  assign tmp33384 = s2 ? tmp33385 : tmp33393;
  assign tmp33370 = ~(s3 ? tmp33371 : tmp33384);
  assign tmp33338 = s4 ? tmp33339 : tmp33370;
  assign tmp33337 = s5 ? 1 : tmp33338;
  assign tmp33407 = ~(l1 ? tmp33380 : 1);
  assign tmp33406 = s0 ? tmp33354 : tmp33407;
  assign tmp33409 = l1 ? tmp33380 : 1;
  assign tmp33408 = ~(s0 ? tmp33409 : tmp33358);
  assign tmp33405 = s1 ? tmp33406 : tmp33408;
  assign tmp33413 = l2 ? tmp33360 : 0;
  assign tmp33414 = l2 ? tmp33345 : tmp33360;
  assign tmp33412 = l1 ? tmp33413 : tmp33414;
  assign tmp33411 = s0 ? tmp33409 : tmp33412;
  assign tmp33416 = l1 ? tmp33396 : tmp33397;
  assign tmp33418 = l2 ? tmp33360 : 1;
  assign tmp33417 = l1 ? tmp33418 : 1;
  assign tmp33415 = s0 ? tmp33416 : tmp33417;
  assign tmp33410 = ~(s1 ? tmp33411 : tmp33415);
  assign tmp33404 = s2 ? tmp33405 : tmp33410;
  assign tmp33423 = l2 ? tmp33360 : tmp33348;
  assign tmp33422 = l1 ? tmp33423 : tmp33414;
  assign tmp33421 = s0 ? tmp33417 : tmp33422;
  assign tmp33427 = ~(l3 ? 1 : tmp33346);
  assign tmp33426 = ~(l2 ? tmp33345 : tmp33427);
  assign tmp33425 = ~(l1 ? tmp33344 : tmp33426);
  assign tmp33424 = s0 ? tmp33417 : tmp33425;
  assign tmp33420 = s1 ? tmp33421 : tmp33424;
  assign tmp33431 = l2 ? tmp33389 : tmp33346;
  assign tmp33432 = l2 ? 1 : tmp33389;
  assign tmp33430 = ~(l1 ? tmp33431 : tmp33432);
  assign tmp33429 = s0 ? tmp33399 : tmp33430;
  assign tmp33435 = l2 ? tmp33348 : 0;
  assign tmp33434 = l1 ? tmp33435 : tmp33397;
  assign tmp33433 = ~(s0 ? tmp33434 : tmp33416);
  assign tmp33428 = ~(s1 ? tmp33429 : tmp33433);
  assign tmp33419 = ~(s2 ? tmp33420 : tmp33428);
  assign tmp33403 = s3 ? tmp33404 : tmp33419;
  assign tmp33441 = l2 ? tmp33345 : tmp33389;
  assign tmp33440 = l1 ? tmp33389 : tmp33441;
  assign tmp33439 = s0 ? tmp33440 : tmp33434;
  assign tmp33444 = ~(l2 ? tmp33353 : 0);
  assign tmp33443 = l1 ? 1 : tmp33444;
  assign tmp33445 = l1 ? 1 : tmp33418;
  assign tmp33442 = ~(s0 ? tmp33443 : tmp33445);
  assign tmp33438 = s1 ? tmp33439 : tmp33442;
  assign tmp33448 = l1 ? tmp33361 : tmp33444;
  assign tmp33451 = l3 ? 1 : 0;
  assign tmp33450 = l2 ? tmp33451 : 1;
  assign tmp33449 = l1 ? tmp33361 : tmp33450;
  assign tmp33447 = s0 ? tmp33448 : tmp33449;
  assign tmp33454 = ~(l2 ? tmp33346 : tmp33427);
  assign tmp33453 = l1 ? tmp33344 : tmp33454;
  assign tmp33452 = s0 ? tmp33453 : tmp33448;
  assign tmp33446 = ~(s1 ? tmp33447 : tmp33452);
  assign tmp33437 = s2 ? tmp33438 : tmp33446;
  assign tmp33459 = l2 ? tmp33360 : tmp33345;
  assign tmp33458 = l1 ? tmp33344 : tmp33459;
  assign tmp33457 = s0 ? tmp33453 : tmp33458;
  assign tmp33461 = l1 ? tmp33344 : tmp33392;
  assign tmp33460 = s0 ? tmp33449 : tmp33461;
  assign tmp33456 = s1 ? tmp33457 : tmp33460;
  assign tmp33465 = l2 ? tmp33389 : 1;
  assign tmp33464 = l1 ? 1 : tmp33465;
  assign tmp33466 = l1 ? tmp33465 : tmp33389;
  assign tmp33463 = s0 ? tmp33464 : tmp33466;
  assign tmp33467 = s0 ? tmp33391 : tmp33466;
  assign tmp33462 = s1 ? tmp33463 : tmp33467;
  assign tmp33455 = ~(s2 ? tmp33456 : tmp33462);
  assign tmp33436 = ~(s3 ? tmp33437 : tmp33455);
  assign tmp33402 = s4 ? tmp33403 : tmp33436;
  assign tmp33473 = l1 ? tmp33344 : tmp33426;
  assign tmp33474 = ~(l1 ? tmp33389 : 1);
  assign tmp33472 = s0 ? tmp33473 : tmp33474;
  assign tmp33476 = l1 ? tmp33432 : tmp33344;
  assign tmp33475 = ~(s0 ? 1 : tmp33476);
  assign tmp33471 = s1 ? tmp33472 : tmp33475;
  assign tmp33478 = s0 ? 1 : tmp33361;
  assign tmp33479 = s0 ? tmp33361 : 1;
  assign tmp33477 = ~(s1 ? tmp33478 : tmp33479);
  assign tmp33470 = s2 ? tmp33471 : tmp33477;
  assign tmp33484 = l2 ? 1 : tmp33345;
  assign tmp33483 = l1 ? tmp33484 : tmp33432;
  assign tmp33482 = s0 ? 1 : tmp33483;
  assign tmp33487 = l2 ? 1 : tmp33346;
  assign tmp33486 = l1 ? tmp33487 : tmp33432;
  assign tmp33485 = s0 ? 1 : tmp33486;
  assign tmp33481 = s1 ? tmp33482 : tmp33485;
  assign tmp33489 = s0 ? 1 : tmp33440;
  assign tmp33491 = l1 ? tmp33361 : tmp33414;
  assign tmp33490 = s0 ? 1 : tmp33491;
  assign tmp33488 = s1 ? tmp33489 : tmp33490;
  assign tmp33480 = ~(s2 ? tmp33481 : tmp33488);
  assign tmp33469 = s3 ? tmp33470 : tmp33480;
  assign tmp33496 = l1 ? tmp33487 : 1;
  assign tmp33495 = s0 ? 1 : tmp33496;
  assign tmp33498 = ~(l1 ? tmp33344 : tmp33400);
  assign tmp33497 = s0 ? 1 : tmp33498;
  assign tmp33494 = s1 ? tmp33495 : tmp33497;
  assign tmp33502 = l2 ? 1 : tmp33353;
  assign tmp33501 = l1 ? tmp33502 : tmp33414;
  assign tmp33500 = s0 ? 1 : tmp33501;
  assign tmp33499 = s1 ? tmp33500 : 1;
  assign tmp33493 = s2 ? tmp33494 : tmp33499;
  assign tmp33506 = ~(l1 ? tmp33344 : tmp33484);
  assign tmp33505 = s0 ? 1 : tmp33506;
  assign tmp33504 = s1 ? tmp33485 : tmp33505;
  assign tmp33503 = s2 ? tmp33504 : 1;
  assign tmp33492 = ~(s3 ? tmp33493 : tmp33503);
  assign tmp33468 = s4 ? tmp33469 : tmp33492;
  assign tmp33401 = ~(s5 ? tmp33402 : tmp33468);
  assign tmp33336 = s6 ? tmp33337 : tmp33401;
  assign tmp33514 = ~(l1 ? 1 : tmp33347);
  assign tmp33513 = s0 ? 1 : tmp33514;
  assign tmp33516 = l1 ? 1 : tmp33347;
  assign tmp33515 = ~(s0 ? tmp33351 : tmp33516);
  assign tmp33512 = s1 ? tmp33513 : tmp33515;
  assign tmp33511 = s2 ? 1 : tmp33512;
  assign tmp33521 = l2 ? tmp33451 : tmp33349;
  assign tmp33520 = l1 ? tmp33521 : tmp33361;
  assign tmp33522 = ~(l1 ? 1 : tmp33363);
  assign tmp33519 = s0 ? tmp33520 : tmp33522;
  assign tmp33524 = l1 ? 1 : tmp33363;
  assign tmp33523 = ~(s0 ? tmp33351 : tmp33524);
  assign tmp33518 = s1 ? tmp33519 : tmp33523;
  assign tmp33526 = s0 ? tmp33524 : tmp33516;
  assign tmp33525 = ~(s1 ? tmp33351 : tmp33526);
  assign tmp33517 = s2 ? tmp33518 : tmp33525;
  assign tmp33510 = s3 ? tmp33511 : tmp33517;
  assign tmp33530 = s0 ? tmp33516 : tmp33374;
  assign tmp33531 = s0 ? tmp33516 : tmp33524;
  assign tmp33529 = s1 ? tmp33530 : tmp33531;
  assign tmp33533 = s0 ? tmp33516 : tmp33379;
  assign tmp33534 = s0 ? tmp33382 : 0;
  assign tmp33532 = s1 ? tmp33533 : tmp33534;
  assign tmp33528 = s2 ? tmp33529 : tmp33532;
  assign tmp33538 = ~(l1 ? 1 : tmp33352);
  assign tmp33537 = s0 ? 1 : tmp33538;
  assign tmp33540 = ~(l1 ? 1 : tmp33392);
  assign tmp33539 = s0 ? 1 : tmp33540;
  assign tmp33536 = s1 ? tmp33537 : tmp33539;
  assign tmp33543 = ~(l1 ? tmp33353 : tmp33397);
  assign tmp33542 = s0 ? tmp33524 : tmp33543;
  assign tmp33545 = l1 ? 1 : tmp33400;
  assign tmp33544 = s0 ? tmp33545 : tmp33524;
  assign tmp33541 = ~(s1 ? tmp33542 : tmp33544);
  assign tmp33535 = ~(s2 ? tmp33536 : tmp33541);
  assign tmp33527 = ~(s3 ? tmp33528 : tmp33535);
  assign tmp33509 = s4 ? tmp33510 : tmp33527;
  assign tmp33508 = s5 ? 1 : tmp33509;
  assign tmp33551 = s0 ? tmp33516 : tmp33407;
  assign tmp33552 = ~(s0 ? 1 : tmp33520);
  assign tmp33550 = s1 ? tmp33551 : tmp33552;
  assign tmp33556 = l2 ? tmp33451 : 0;
  assign tmp33555 = l1 ? tmp33556 : tmp33414;
  assign tmp33554 = s0 ? 1 : tmp33555;
  assign tmp33558 = l1 ? tmp33353 : tmp33397;
  assign tmp33557 = s0 ? tmp33558 : tmp33417;
  assign tmp33553 = ~(s1 ? tmp33554 : tmp33557);
  assign tmp33549 = s2 ? tmp33550 : tmp33553;
  assign tmp33563 = l2 ? tmp33451 : tmp33348;
  assign tmp33562 = l1 ? tmp33563 : tmp33414;
  assign tmp33561 = s0 ? 1 : tmp33562;
  assign tmp33565 = ~(l1 ? 1 : tmp33426);
  assign tmp33564 = s0 ? 1 : tmp33565;
  assign tmp33560 = s1 ? tmp33561 : tmp33564;
  assign tmp33567 = s0 ? tmp33545 : tmp33430;
  assign tmp33570 = l2 ? tmp33353 : 0;
  assign tmp33569 = l1 ? tmp33570 : tmp33397;
  assign tmp33568 = ~(s0 ? tmp33569 : tmp33558);
  assign tmp33566 = ~(s1 ? tmp33567 : tmp33568);
  assign tmp33559 = ~(s2 ? tmp33560 : tmp33566);
  assign tmp33548 = s3 ? tmp33549 : tmp33559;
  assign tmp33574 = s0 ? tmp33440 : tmp33569;
  assign tmp33573 = s1 ? tmp33574 : tmp33442;
  assign tmp33576 = s0 ? tmp33448 : 0;
  assign tmp33578 = l1 ? 1 : tmp33454;
  assign tmp33577 = s0 ? tmp33578 : tmp33448;
  assign tmp33575 = ~(s1 ? tmp33576 : tmp33577);
  assign tmp33572 = s2 ? tmp33573 : tmp33575;
  assign tmp33582 = l1 ? 1 : tmp33459;
  assign tmp33581 = s0 ? tmp33578 : tmp33582;
  assign tmp33583 = ~(s0 ? 1 : tmp33540);
  assign tmp33580 = s1 ? tmp33581 : tmp33583;
  assign tmp33585 = s0 ? tmp33464 : 0;
  assign tmp33586 = s0 ? tmp33391 : 0;
  assign tmp33584 = s1 ? tmp33585 : tmp33586;
  assign tmp33579 = ~(s2 ? tmp33580 : tmp33584);
  assign tmp33571 = ~(s3 ? tmp33572 : tmp33579);
  assign tmp33547 = s4 ? tmp33548 : tmp33571;
  assign tmp33592 = l1 ? 1 : tmp33426;
  assign tmp33591 = s0 ? tmp33592 : tmp33474;
  assign tmp33594 = l1 ? tmp33441 : tmp33344;
  assign tmp33593 = ~(s0 ? 1 : tmp33594);
  assign tmp33590 = s1 ? tmp33591 : tmp33593;
  assign tmp33597 = l1 ? tmp33414 : tmp33361;
  assign tmp33596 = s0 ? 1 : tmp33597;
  assign tmp33598 = s0 ? tmp33597 : 1;
  assign tmp33595 = ~(s1 ? tmp33596 : tmp33598);
  assign tmp33589 = s2 ? tmp33590 : tmp33595;
  assign tmp33601 = s0 ? 1 : tmp33414;
  assign tmp33600 = s1 ? tmp33489 : tmp33601;
  assign tmp33599 = ~(s2 ? tmp33481 : tmp33600);
  assign tmp33588 = s3 ? tmp33589 : tmp33599;
  assign tmp33607 = l2 ? tmp33345 : tmp33346;
  assign tmp33606 = l1 ? tmp33607 : 1;
  assign tmp33605 = s0 ? 1 : tmp33606;
  assign tmp33609 = ~(l1 ? 1 : tmp33400);
  assign tmp33608 = s0 ? 1 : tmp33609;
  assign tmp33604 = s1 ? tmp33605 : tmp33608;
  assign tmp33613 = l2 ? tmp33345 : tmp33353;
  assign tmp33612 = l1 ? tmp33613 : tmp33414;
  assign tmp33611 = s0 ? 1 : tmp33612;
  assign tmp33610 = s1 ? tmp33611 : 1;
  assign tmp33603 = s2 ? tmp33604 : tmp33610;
  assign tmp33617 = l1 ? tmp33607 : tmp33432;
  assign tmp33616 = s0 ? 1 : tmp33617;
  assign tmp33619 = ~(l1 ? 1 : tmp33484);
  assign tmp33618 = s0 ? 1 : tmp33619;
  assign tmp33615 = s1 ? tmp33616 : tmp33618;
  assign tmp33614 = s2 ? tmp33615 : 1;
  assign tmp33602 = ~(s3 ? tmp33603 : tmp33614);
  assign tmp33587 = s4 ? tmp33588 : tmp33602;
  assign tmp33546 = ~(s5 ? tmp33547 : tmp33587);
  assign tmp33507 = s6 ? tmp33508 : tmp33546;
  assign tmp33335 = s7 ? tmp33336 : tmp33507;
  assign tmp33627 = ~(s0 ? tmp33578 : 0);
  assign tmp33626 = s1 ? 1 : tmp33627;
  assign tmp33625 = s2 ? tmp33573 : tmp33626;
  assign tmp33624 = ~(s3 ? tmp33625 : tmp33579);
  assign tmp33623 = s4 ? tmp33548 : tmp33624;
  assign tmp33622 = ~(s5 ? tmp33623 : tmp33587);
  assign tmp33621 = s6 ? tmp33508 : tmp33622;
  assign tmp33620 = s7 ? tmp33336 : tmp33621;
  assign tmp33334 = s8 ? tmp33335 : tmp33620;
  assign tmp33333 = s9 ? tmp33334 : tmp33620;
  assign tmp33629 = s8 ? tmp33620 : tmp33336;
  assign tmp33638 = s0 ? tmp33578 : 0;
  assign tmp33637 = ~(s1 ? tmp33576 : tmp33638);
  assign tmp33636 = s2 ? tmp33573 : tmp33637;
  assign tmp33635 = ~(s3 ? tmp33636 : tmp33579);
  assign tmp33634 = s4 ? tmp33548 : tmp33635;
  assign tmp33633 = ~(s5 ? tmp33634 : tmp33587);
  assign tmp33632 = s6 ? tmp33508 : tmp33633;
  assign tmp33631 = s7 ? tmp33632 : tmp33621;
  assign tmp33630 = s8 ? tmp33631 : tmp33621;
  assign tmp33628 = s9 ? tmp33629 : tmp33630;
  assign tmp33332 = s10 ? tmp33333 : tmp33628;
  assign tmp33642 = s7 ? tmp33507 : tmp33621;
  assign tmp33641 = s8 ? tmp33642 : tmp33621;
  assign tmp33640 = s9 ? tmp33629 : tmp33641;
  assign tmp33639 = s10 ? tmp33333 : tmp33640;
  assign tmp33331 = s11 ? tmp33332 : tmp33639;
  assign tmp33330 = s12 ? 1 : tmp33331;
  assign tmp33654 = s1 ? tmp33533 : tmp33381;
  assign tmp33653 = s2 ? tmp33529 : tmp33654;
  assign tmp33657 = ~(s0 ? tmp33379 : tmp33391);
  assign tmp33656 = s1 ? tmp33537 : tmp33657;
  assign tmp33655 = ~(s2 ? tmp33656 : tmp33541);
  assign tmp33652 = ~(s3 ? tmp33653 : tmp33655);
  assign tmp33651 = s4 ? tmp33510 : tmp33652;
  assign tmp33650 = s5 ? 1 : tmp33651;
  assign tmp33663 = ~(s0 ? tmp33409 : tmp33520);
  assign tmp33662 = s1 ? tmp33551 : tmp33663;
  assign tmp33665 = s0 ? tmp33409 : tmp33555;
  assign tmp33664 = ~(s1 ? tmp33665 : tmp33557);
  assign tmp33661 = s2 ? tmp33662 : tmp33664;
  assign tmp33668 = s0 ? tmp33417 : tmp33562;
  assign tmp33669 = s0 ? tmp33417 : tmp33565;
  assign tmp33667 = s1 ? tmp33668 : tmp33669;
  assign tmp33666 = ~(s2 ? tmp33667 : tmp33566);
  assign tmp33660 = s3 ? tmp33661 : tmp33666;
  assign tmp33659 = s4 ? tmp33660 : tmp33624;
  assign tmp33658 = ~(s5 ? tmp33659 : tmp33587);
  assign tmp33649 = s6 ? tmp33650 : tmp33658;
  assign tmp33648 = s7 ? tmp33336 : tmp33649;
  assign tmp33674 = s3 ? tmp33661 : tmp33559;
  assign tmp33673 = s4 ? tmp33674 : tmp33624;
  assign tmp33672 = ~(s5 ? tmp33673 : tmp33587);
  assign tmp33671 = s6 ? tmp33508 : tmp33672;
  assign tmp33670 = s7 ? tmp33336 : tmp33671;
  assign tmp33647 = s8 ? tmp33648 : tmp33670;
  assign tmp33646 = s9 ? tmp33647 : tmp33670;
  assign tmp33676 = s8 ? tmp33670 : tmp33336;
  assign tmp33682 = ~(s3 ? tmp33653 : tmp33535);
  assign tmp33681 = s4 ? tmp33510 : tmp33682;
  assign tmp33680 = s5 ? 1 : tmp33681;
  assign tmp33686 = s2 ? tmp33662 : tmp33553;
  assign tmp33688 = s1 ? tmp33668 : tmp33564;
  assign tmp33687 = ~(s2 ? tmp33688 : tmp33566);
  assign tmp33685 = s3 ? tmp33686 : tmp33687;
  assign tmp33684 = s4 ? tmp33685 : tmp33624;
  assign tmp33683 = ~(s5 ? tmp33684 : tmp33587);
  assign tmp33679 = s6 ? tmp33680 : tmp33683;
  assign tmp33692 = s3 ? tmp33686 : tmp33559;
  assign tmp33691 = s4 ? tmp33692 : tmp33624;
  assign tmp33690 = ~(s5 ? tmp33691 : tmp33587);
  assign tmp33689 = s6 ? tmp33508 : tmp33690;
  assign tmp33678 = s7 ? tmp33679 : tmp33689;
  assign tmp33677 = s8 ? tmp33678 : tmp33689;
  assign tmp33675 = s9 ? tmp33676 : tmp33677;
  assign tmp33645 = s10 ? tmp33646 : tmp33675;
  assign tmp33696 = s7 ? tmp33649 : tmp33671;
  assign tmp33695 = s8 ? tmp33696 : tmp33671;
  assign tmp33694 = s9 ? tmp33676 : tmp33695;
  assign tmp33693 = s10 ? tmp33646 : tmp33694;
  assign tmp33644 = s11 ? tmp33645 : tmp33693;
  assign tmp33702 = s6 ? tmp33650 : tmp33622;
  assign tmp33701 = s7 ? tmp33336 : tmp33702;
  assign tmp33700 = s8 ? tmp33701 : tmp33620;
  assign tmp33699 = s9 ? tmp33700 : tmp33620;
  assign tmp33706 = s6 ? tmp33680 : tmp33622;
  assign tmp33705 = s7 ? tmp33706 : tmp33621;
  assign tmp33704 = s8 ? tmp33705 : tmp33621;
  assign tmp33703 = s9 ? tmp33629 : tmp33704;
  assign tmp33698 = s10 ? tmp33699 : tmp33703;
  assign tmp33710 = s7 ? tmp33702 : tmp33621;
  assign tmp33709 = s8 ? tmp33710 : tmp33621;
  assign tmp33708 = s9 ? tmp33629 : tmp33709;
  assign tmp33707 = s10 ? tmp33699 : tmp33708;
  assign tmp33697 = s11 ? tmp33698 : tmp33707;
  assign tmp33643 = s12 ? tmp33644 : tmp33697;
  assign tmp33329 = s13 ? tmp33330 : tmp33643;
  assign tmp33721 = s3 ? tmp33549 : tmp33666;
  assign tmp33720 = s4 ? tmp33721 : tmp33624;
  assign tmp33719 = ~(s5 ? tmp33720 : tmp33587);
  assign tmp33718 = s6 ? tmp33508 : tmp33719;
  assign tmp33717 = s7 ? tmp33336 : tmp33718;
  assign tmp33716 = s8 ? tmp33717 : tmp33620;
  assign tmp33715 = s9 ? tmp33716 : tmp33620;
  assign tmp33728 = s3 ? tmp33549 : tmp33687;
  assign tmp33727 = s4 ? tmp33728 : tmp33624;
  assign tmp33726 = ~(s5 ? tmp33727 : tmp33587);
  assign tmp33725 = s6 ? tmp33508 : tmp33726;
  assign tmp33724 = s7 ? tmp33725 : tmp33621;
  assign tmp33723 = s8 ? tmp33724 : tmp33621;
  assign tmp33722 = s9 ? tmp33629 : tmp33723;
  assign tmp33714 = s10 ? tmp33715 : tmp33722;
  assign tmp33732 = s7 ? tmp33718 : tmp33621;
  assign tmp33731 = s8 ? tmp33732 : tmp33621;
  assign tmp33730 = s9 ? tmp33629 : tmp33731;
  assign tmp33729 = s10 ? tmp33715 : tmp33730;
  assign tmp33713 = s11 ? tmp33714 : tmp33729;
  assign tmp33745 = ~(l1 ? tmp33361 : tmp33450);
  assign tmp33744 = s0 ? 1 : tmp33745;
  assign tmp33743 = s1 ? tmp33744 : tmp33627;
  assign tmp33742 = s2 ? tmp33573 : tmp33743;
  assign tmp33748 = s0 ? tmp33449 : tmp33391;
  assign tmp33747 = s1 ? tmp33581 : tmp33748;
  assign tmp33746 = ~(s2 ? tmp33747 : tmp33584);
  assign tmp33741 = ~(s3 ? tmp33742 : tmp33746);
  assign tmp33740 = s4 ? tmp33548 : tmp33741;
  assign tmp33739 = ~(s5 ? tmp33740 : tmp33587);
  assign tmp33738 = s6 ? tmp33508 : tmp33739;
  assign tmp33737 = s7 ? tmp33336 : tmp33738;
  assign tmp33736 = s8 ? tmp33737 : tmp33620;
  assign tmp33735 = s9 ? tmp33736 : tmp33620;
  assign tmp33755 = ~(s3 ? tmp33742 : tmp33579);
  assign tmp33754 = s4 ? tmp33548 : tmp33755;
  assign tmp33753 = ~(s5 ? tmp33754 : tmp33587);
  assign tmp33752 = s6 ? tmp33508 : tmp33753;
  assign tmp33751 = s7 ? tmp33752 : tmp33621;
  assign tmp33750 = s8 ? tmp33751 : tmp33621;
  assign tmp33749 = s9 ? tmp33629 : tmp33750;
  assign tmp33734 = s10 ? tmp33735 : tmp33749;
  assign tmp33759 = s7 ? tmp33738 : tmp33621;
  assign tmp33758 = s8 ? tmp33759 : tmp33621;
  assign tmp33757 = s9 ? tmp33629 : tmp33758;
  assign tmp33756 = s10 ? tmp33735 : tmp33757;
  assign tmp33733 = s11 ? tmp33734 : tmp33756;
  assign tmp33712 = s12 ? tmp33713 : tmp33733;
  assign tmp33767 = s1 ? tmp33378 : tmp33534;
  assign tmp33766 = s2 ? tmp33372 : tmp33767;
  assign tmp33769 = ~(s1 ? tmp33394 : tmp33398);
  assign tmp33768 = ~(s2 ? tmp33536 : tmp33769);
  assign tmp33765 = ~(s3 ? tmp33766 : tmp33768);
  assign tmp33764 = s4 ? tmp33339 : tmp33765;
  assign tmp33763 = s5 ? 1 : tmp33764;
  assign tmp33775 = ~(s0 ? 1 : tmp33358);
  assign tmp33774 = s1 ? tmp33406 : tmp33775;
  assign tmp33777 = s0 ? 1 : tmp33412;
  assign tmp33776 = ~(s1 ? tmp33777 : tmp33415);
  assign tmp33773 = s2 ? tmp33774 : tmp33776;
  assign tmp33780 = s0 ? 1 : tmp33422;
  assign tmp33781 = s0 ? 1 : tmp33425;
  assign tmp33779 = s1 ? tmp33780 : tmp33781;
  assign tmp33778 = ~(s2 ? tmp33779 : tmp33428);
  assign tmp33772 = s3 ? tmp33773 : tmp33778;
  assign tmp33785 = ~(s0 ? tmp33453 : 0);
  assign tmp33784 = s1 ? 1 : tmp33785;
  assign tmp33783 = s2 ? tmp33438 : tmp33784;
  assign tmp33789 = ~(l1 ? tmp33344 : tmp33392);
  assign tmp33788 = ~(s0 ? 1 : tmp33789);
  assign tmp33787 = s1 ? tmp33457 : tmp33788;
  assign tmp33786 = ~(s2 ? tmp33787 : tmp33584);
  assign tmp33782 = ~(s3 ? tmp33783 : tmp33786);
  assign tmp33771 = s4 ? tmp33772 : tmp33782;
  assign tmp33770 = ~(s5 ? tmp33771 : tmp33468);
  assign tmp33762 = s6 ? tmp33763 : tmp33770;
  assign tmp33761 = s7 ? tmp33336 : tmp33762;
  assign tmp33791 = s8 ? tmp33761 : tmp33336;
  assign tmp33790 = s9 ? tmp33791 : tmp33762;
  assign tmp33760 = s10 ? tmp33761 : tmp33790;
  assign tmp33711 = s13 ? tmp33712 : tmp33760;
  assign tmp33328 = s14 ? tmp33329 : tmp33711;
  assign tmp33796 = s9 ? tmp33629 : tmp33621;
  assign tmp33795 = s10 ? tmp33620 : tmp33796;
  assign tmp33804 = ~(s2 ? tmp33580 : tmp33462);
  assign tmp33803 = ~(s3 ? tmp33625 : tmp33804);
  assign tmp33802 = s4 ? tmp33548 : tmp33803;
  assign tmp33801 = ~(s5 ? tmp33802 : tmp33587);
  assign tmp33800 = s6 ? tmp33508 : tmp33801;
  assign tmp33799 = s7 ? tmp33336 : tmp33800;
  assign tmp33806 = s8 ? tmp33799 : tmp33336;
  assign tmp33812 = s1 ? tmp33463 : tmp33586;
  assign tmp33811 = ~(s2 ? tmp33580 : tmp33812);
  assign tmp33810 = ~(s3 ? tmp33625 : tmp33811);
  assign tmp33809 = s4 ? tmp33548 : tmp33810;
  assign tmp33808 = ~(s5 ? tmp33809 : tmp33587);
  assign tmp33807 = s6 ? tmp33508 : tmp33808;
  assign tmp33805 = s9 ? tmp33806 : tmp33807;
  assign tmp33798 = s10 ? tmp33799 : tmp33805;
  assign tmp33814 = s9 ? tmp33806 : tmp33800;
  assign tmp33813 = s10 ? tmp33799 : tmp33814;
  assign tmp33797 = s11 ? tmp33798 : tmp33813;
  assign tmp33794 = s12 ? tmp33795 : tmp33797;
  assign tmp33793 = s13 ? tmp33794 : tmp33795;
  assign tmp33827 = s1 ? tmp33744 : tmp33785;
  assign tmp33826 = s2 ? tmp33438 : tmp33827;
  assign tmp33828 = ~(s2 ? tmp33456 : tmp33584);
  assign tmp33825 = ~(s3 ? tmp33826 : tmp33828);
  assign tmp33824 = s4 ? tmp33772 : tmp33825;
  assign tmp33823 = ~(s5 ? tmp33824 : tmp33468);
  assign tmp33822 = s6 ? tmp33763 : tmp33823;
  assign tmp33821 = s7 ? tmp33336 : tmp33822;
  assign tmp33820 = s8 ? tmp33821 : tmp33761;
  assign tmp33819 = s9 ? tmp33820 : tmp33761;
  assign tmp33835 = ~(s3 ? tmp33826 : tmp33786);
  assign tmp33834 = s4 ? tmp33772 : tmp33835;
  assign tmp33833 = ~(s5 ? tmp33834 : tmp33468);
  assign tmp33832 = s6 ? tmp33763 : tmp33833;
  assign tmp33831 = s7 ? tmp33832 : tmp33762;
  assign tmp33830 = s8 ? tmp33831 : tmp33762;
  assign tmp33829 = s9 ? tmp33791 : tmp33830;
  assign tmp33818 = s10 ? tmp33819 : tmp33829;
  assign tmp33839 = s7 ? tmp33822 : tmp33762;
  assign tmp33838 = s8 ? tmp33839 : tmp33762;
  assign tmp33837 = s9 ? tmp33791 : tmp33838;
  assign tmp33836 = s10 ? tmp33819 : tmp33837;
  assign tmp33817 = s11 ? tmp33818 : tmp33836;
  assign tmp33816 = s12 ? tmp33817 : tmp33760;
  assign tmp33840 = s12 ? tmp33795 : tmp33760;
  assign tmp33815 = s13 ? tmp33816 : tmp33840;
  assign tmp33792 = s14 ? tmp33793 : tmp33815;
  assign tmp33327 = s15 ? tmp33328 : tmp33792;
  assign tmp33848 = s8 ? tmp33335 : tmp33336;
  assign tmp33847 = s9 ? tmp33848 : tmp33632;
  assign tmp33846 = s10 ? tmp33335 : tmp33847;
  assign tmp33850 = s9 ? tmp33848 : tmp33507;
  assign tmp33849 = s10 ? tmp33335 : tmp33850;
  assign tmp33845 = s11 ? tmp33846 : tmp33849;
  assign tmp33844 = s12 ? 1 : tmp33845;
  assign tmp33855 = s8 ? tmp33701 : tmp33336;
  assign tmp33854 = s9 ? tmp33855 : tmp33706;
  assign tmp33853 = s10 ? tmp33701 : tmp33854;
  assign tmp33857 = s9 ? tmp33855 : tmp33702;
  assign tmp33856 = s10 ? tmp33701 : tmp33857;
  assign tmp33852 = s11 ? tmp33853 : tmp33856;
  assign tmp33851 = s12 ? tmp33644 : tmp33852;
  assign tmp33843 = s13 ? tmp33844 : tmp33851;
  assign tmp33863 = s8 ? tmp33717 : tmp33336;
  assign tmp33862 = s9 ? tmp33863 : tmp33725;
  assign tmp33861 = s10 ? tmp33717 : tmp33862;
  assign tmp33865 = s9 ? tmp33863 : tmp33718;
  assign tmp33864 = s10 ? tmp33717 : tmp33865;
  assign tmp33860 = s11 ? tmp33861 : tmp33864;
  assign tmp33869 = s8 ? tmp33737 : tmp33336;
  assign tmp33868 = s9 ? tmp33869 : tmp33752;
  assign tmp33867 = s10 ? tmp33737 : tmp33868;
  assign tmp33871 = s9 ? tmp33869 : tmp33738;
  assign tmp33870 = s10 ? tmp33737 : tmp33871;
  assign tmp33866 = s11 ? tmp33867 : tmp33870;
  assign tmp33859 = s12 ? tmp33860 : tmp33866;
  assign tmp33858 = s13 ? tmp33859 : tmp33760;
  assign tmp33842 = s14 ? tmp33843 : tmp33858;
  assign tmp33841 = s15 ? tmp33842 : tmp33792;
  assign tmp33326 = s16 ? tmp33327 : tmp33841;
  assign tmp33879 = s9 ? tmp33335 : tmp33334;
  assign tmp33880 = s9 ? tmp33629 : tmp33631;
  assign tmp33878 = s10 ? tmp33879 : tmp33880;
  assign tmp33882 = s9 ? tmp33629 : tmp33642;
  assign tmp33881 = s10 ? tmp33879 : tmp33882;
  assign tmp33877 = s11 ? tmp33878 : tmp33881;
  assign tmp33876 = s12 ? 1 : tmp33877;
  assign tmp33886 = s9 ? tmp33701 : tmp33700;
  assign tmp33887 = s9 ? tmp33629 : tmp33705;
  assign tmp33885 = s10 ? tmp33886 : tmp33887;
  assign tmp33889 = s9 ? tmp33629 : tmp33710;
  assign tmp33888 = s10 ? tmp33886 : tmp33889;
  assign tmp33884 = s11 ? tmp33885 : tmp33888;
  assign tmp33883 = s12 ? tmp33644 : tmp33884;
  assign tmp33875 = s13 ? tmp33876 : tmp33883;
  assign tmp33894 = s9 ? tmp33717 : tmp33716;
  assign tmp33895 = s9 ? tmp33629 : tmp33724;
  assign tmp33893 = s10 ? tmp33894 : tmp33895;
  assign tmp33897 = s9 ? tmp33629 : tmp33732;
  assign tmp33896 = s10 ? tmp33894 : tmp33897;
  assign tmp33892 = s11 ? tmp33893 : tmp33896;
  assign tmp33900 = s9 ? tmp33737 : tmp33736;
  assign tmp33901 = s9 ? tmp33629 : tmp33751;
  assign tmp33899 = s10 ? tmp33900 : tmp33901;
  assign tmp33903 = s9 ? tmp33629 : tmp33759;
  assign tmp33902 = s10 ? tmp33900 : tmp33903;
  assign tmp33898 = s11 ? tmp33899 : tmp33902;
  assign tmp33891 = s12 ? tmp33892 : tmp33898;
  assign tmp33890 = s13 ? tmp33891 : tmp33760;
  assign tmp33874 = s14 ? tmp33875 : tmp33890;
  assign tmp33873 = s15 ? tmp33874 : tmp33792;
  assign tmp33872 = s16 ? tmp33873 : tmp33841;
  assign tmp33325 = s17 ? tmp33326 : tmp33872;
  assign tmp33324 = ~(s18 ? 1 : tmp33325);
  assign s4n = tmp33324;

  assign tmp33920 = l4 ? 1 : 0;
  assign tmp33921 = ~(l4 ? 1 : 0);
  assign tmp33919 = l2 ? tmp33920 : tmp33921;
  assign tmp33923 = l3 ? 1 : 0;
  assign tmp33924 = ~(l3 ? tmp33920 : tmp33921);
  assign tmp33922 = l2 ? tmp33923 : tmp33924;
  assign tmp33918 = l1 ? tmp33919 : tmp33922;
  assign tmp33927 = l2 ? 1 : tmp33921;
  assign tmp33929 = ~(l3 ? tmp33920 : 0);
  assign tmp33928 = l2 ? tmp33923 : tmp33929;
  assign tmp33926 = l1 ? tmp33927 : tmp33928;
  assign tmp33932 = l3 ? 1 : tmp33920;
  assign tmp33931 = l2 ? tmp33932 : tmp33921;
  assign tmp33930 = l1 ? tmp33931 : tmp33922;
  assign tmp33925 = s0 ? tmp33926 : tmp33930;
  assign tmp33917 = s1 ? tmp33918 : tmp33925;
  assign tmp33938 = l3 ? 1 : tmp33921;
  assign tmp33937 = l2 ? tmp33938 : 1;
  assign tmp33939 = l2 ? 1 : tmp33938;
  assign tmp33936 = l1 ? tmp33937 : tmp33939;
  assign tmp33942 = l3 ? tmp33920 : 1;
  assign tmp33943 = l3 ? tmp33920 : tmp33921;
  assign tmp33941 = ~(l2 ? tmp33942 : tmp33943);
  assign tmp33940 = ~(l1 ? tmp33919 : tmp33941);
  assign tmp33935 = s0 ? tmp33936 : tmp33940;
  assign tmp33946 = l2 ? tmp33938 : tmp33942;
  assign tmp33948 = l3 ? tmp33920 : 0;
  assign tmp33949 = ~(l3 ? 1 : tmp33921);
  assign tmp33947 = ~(l2 ? tmp33948 : tmp33949);
  assign tmp33945 = l1 ? tmp33946 : tmp33947;
  assign tmp33944 = s0 ? tmp33945 : tmp33940;
  assign tmp33934 = s1 ? tmp33935 : tmp33944;
  assign tmp33952 = l1 ? tmp33937 : 1;
  assign tmp33951 = s0 ? tmp33945 : tmp33952;
  assign tmp33954 = l1 ? tmp33919 : tmp33941;
  assign tmp33953 = ~(s0 ? tmp33954 : tmp33918);
  assign tmp33950 = s1 ? tmp33951 : tmp33953;
  assign tmp33933 = ~(s2 ? tmp33934 : tmp33950);
  assign tmp33916 = s3 ? tmp33917 : tmp33933;
  assign tmp33959 = l1 ? tmp33937 : tmp33947;
  assign tmp33960 = ~(l1 ? tmp33927 : tmp33929);
  assign tmp33958 = s0 ? tmp33959 : tmp33960;
  assign tmp33961 = ~(s0 ? tmp33918 : tmp33954);
  assign tmp33957 = s1 ? tmp33958 : tmp33961;
  assign tmp33964 = l2 ? 1 : tmp33929;
  assign tmp33963 = s0 ? tmp33918 : tmp33964;
  assign tmp33967 = ~(l2 ? tmp33942 : 0);
  assign tmp33966 = l1 ? tmp33927 : tmp33967;
  assign tmp33968 = l1 ? tmp33964 : 1;
  assign tmp33965 = s0 ? tmp33966 : tmp33968;
  assign tmp33962 = ~(s1 ? tmp33963 : tmp33965);
  assign tmp33956 = s2 ? tmp33957 : tmp33962;
  assign tmp33973 = ~(l2 ? tmp33948 : 0);
  assign tmp33972 = l1 ? tmp33927 : tmp33973;
  assign tmp33975 = ~(l2 ? tmp33942 : tmp33948);
  assign tmp33974 = l1 ? tmp33927 : tmp33975;
  assign tmp33971 = s0 ? tmp33972 : tmp33974;
  assign tmp33978 = l2 ? tmp33942 : 1;
  assign tmp33977 = l1 ? tmp33978 : tmp33932;
  assign tmp33976 = s0 ? tmp33968 : tmp33977;
  assign tmp33970 = s1 ? tmp33971 : tmp33976;
  assign tmp33982 = l2 ? tmp33938 : tmp33920;
  assign tmp33983 = l2 ? tmp33942 : tmp33943;
  assign tmp33981 = ~(l1 ? tmp33982 : tmp33983);
  assign tmp33980 = s0 ? tmp33954 : tmp33981;
  assign tmp33986 = l2 ? tmp33920 : 1;
  assign tmp33987 = l2 ? tmp33923 : tmp33932;
  assign tmp33985 = l1 ? tmp33986 : tmp33987;
  assign tmp33984 = s0 ? tmp33985 : tmp33954;
  assign tmp33979 = s1 ? tmp33980 : tmp33984;
  assign tmp33969 = ~(s2 ? tmp33970 : tmp33979);
  assign tmp33955 = ~(s3 ? tmp33956 : tmp33969);
  assign tmp33915 = s4 ? tmp33916 : tmp33955;
  assign tmp33993 = s0 ? tmp33930 : 0;
  assign tmp33995 = l1 ? 1 : tmp33964;
  assign tmp33994 = ~(s0 ? tmp33995 : tmp33936);
  assign tmp33992 = s1 ? tmp33993 : tmp33994;
  assign tmp33998 = l1 ? tmp33982 : tmp33939;
  assign tmp33997 = s0 ? tmp33995 : tmp33998;
  assign tmp34000 = l1 ? tmp33982 : tmp33983;
  assign tmp34002 = ~(l2 ? tmp33920 : tmp33948);
  assign tmp34001 = ~(l1 ? 1 : tmp34002);
  assign tmp33999 = s0 ? tmp34000 : tmp34001;
  assign tmp33996 = ~(s1 ? tmp33997 : tmp33999);
  assign tmp33991 = s2 ? tmp33992 : tmp33996;
  assign tmp34006 = ~(l1 ? tmp33946 : tmp33947);
  assign tmp34005 = s0 ? 1 : tmp34006;
  assign tmp34009 = l2 ? tmp33920 : tmp33938;
  assign tmp34011 = ~(l3 ? 1 : tmp33920);
  assign tmp34010 = ~(l2 ? tmp33942 : tmp34011);
  assign tmp34008 = l1 ? tmp34009 : tmp34010;
  assign tmp34007 = s0 ? 1 : tmp34008;
  assign tmp34004 = s1 ? tmp34005 : tmp34007;
  assign tmp34014 = l1 ? tmp33978 : 1;
  assign tmp34013 = s0 ? tmp33985 : tmp34014;
  assign tmp34016 = l1 ? tmp33919 : tmp34010;
  assign tmp34017 = l1 ? tmp34009 : tmp33987;
  assign tmp34015 = s0 ? tmp34016 : tmp34017;
  assign tmp34012 = s1 ? tmp34013 : tmp34015;
  assign tmp34003 = s2 ? tmp34004 : tmp34012;
  assign tmp33990 = s3 ? tmp33991 : tmp34003;
  assign tmp34021 = s0 ? tmp33977 : tmp34016;
  assign tmp34024 = l2 ? tmp33923 : 1;
  assign tmp34023 = ~(l1 ? tmp33939 : tmp34024);
  assign tmp34022 = ~(s0 ? tmp33952 : tmp34023);
  assign tmp34020 = s1 ? tmp34021 : tmp34022;
  assign tmp34027 = ~(l1 ? tmp33939 : 1);
  assign tmp34026 = s0 ? tmp33952 : tmp34027;
  assign tmp34028 = s0 ? tmp33936 : tmp33952;
  assign tmp34025 = ~(s1 ? tmp34026 : tmp34028);
  assign tmp34019 = s2 ? tmp34020 : tmp34025;
  assign tmp34032 = l1 ? 1 : tmp33939;
  assign tmp34034 = l2 ? 1 : tmp33943;
  assign tmp34033 = l1 ? tmp33946 : tmp34034;
  assign tmp34031 = s0 ? tmp34032 : tmp34033;
  assign tmp34036 = l1 ? tmp33939 : 1;
  assign tmp34037 = l1 ? tmp34009 : tmp33932;
  assign tmp34035 = ~(s0 ? tmp34036 : tmp34037);
  assign tmp34030 = s1 ? tmp34031 : tmp34035;
  assign tmp34039 = s0 ? tmp33977 : tmp34014;
  assign tmp34038 = ~(s1 ? tmp34014 : tmp34039);
  assign tmp34029 = ~(s2 ? tmp34030 : tmp34038);
  assign tmp34018 = s3 ? tmp34019 : tmp34029;
  assign tmp33989 = s4 ? tmp33990 : tmp34018;
  assign tmp34046 = l2 ? 1 : tmp33942;
  assign tmp34045 = ~(l1 ? tmp34046 : tmp33978);
  assign tmp34044 = s0 ? tmp34008 : tmp34045;
  assign tmp34048 = l1 ? tmp34046 : tmp33978;
  assign tmp34050 = l2 ? tmp33932 : 1;
  assign tmp34049 = ~(l1 ? tmp34050 : tmp34024);
  assign tmp34047 = ~(s0 ? tmp34048 : tmp34049);
  assign tmp34043 = s1 ? tmp34044 : tmp34047;
  assign tmp34053 = ~(l1 ? 1 : tmp33939);
  assign tmp34052 = s0 ? 1 : tmp34053;
  assign tmp34056 = l2 ? tmp33932 : tmp33938;
  assign tmp34055 = l1 ? tmp34056 : 1;
  assign tmp34057 = ~(l1 ? tmp34050 : tmp33937);
  assign tmp34054 = s0 ? tmp34055 : tmp34057;
  assign tmp34051 = s1 ? tmp34052 : tmp34054;
  assign tmp34042 = s2 ? tmp34043 : tmp34051;
  assign tmp34062 = l2 ? 1 : tmp33932;
  assign tmp34061 = l1 ? 1 : tmp34062;
  assign tmp34060 = s0 ? tmp33939 : tmp34061;
  assign tmp34059 = s1 ? tmp34060 : 1;
  assign tmp34065 = ~(l2 ? 1 : tmp33942);
  assign tmp34064 = s0 ? 1 : tmp34065;
  assign tmp34068 = l2 ? tmp33932 : tmp33920;
  assign tmp34067 = l1 ? tmp34046 : tmp34068;
  assign tmp34066 = ~(s0 ? tmp34067 : tmp34032);
  assign tmp34063 = s1 ? tmp34064 : tmp34066;
  assign tmp34058 = s2 ? tmp34059 : tmp34063;
  assign tmp34041 = s3 ? tmp34042 : tmp34058;
  assign tmp34073 = l1 ? tmp34050 : tmp33932;
  assign tmp34074 = ~(l1 ? tmp34050 : tmp34062);
  assign tmp34072 = s0 ? tmp34073 : tmp34074;
  assign tmp34075 = ~(s0 ? 1 : tmp33985);
  assign tmp34071 = s1 ? tmp34072 : tmp34075;
  assign tmp34079 = l2 ? 1 : tmp33920;
  assign tmp34078 = l1 ? tmp34079 : tmp33939;
  assign tmp34077 = s0 ? tmp34048 : tmp34078;
  assign tmp34081 = l1 ? tmp34050 : tmp33937;
  assign tmp34082 = ~(l2 ? 1 : tmp33938);
  assign tmp34080 = s0 ? tmp34081 : tmp34082;
  assign tmp34076 = s1 ? tmp34077 : tmp34080;
  assign tmp34070 = s2 ? tmp34071 : tmp34076;
  assign tmp34086 = l1 ? tmp34050 : tmp34062;
  assign tmp34085 = s0 ? 1 : tmp34086;
  assign tmp34088 = ~(l1 ? tmp34079 : tmp34034);
  assign tmp34087 = s0 ? 1 : tmp34088;
  assign tmp34084 = s1 ? tmp34085 : tmp34087;
  assign tmp34090 = s0 ? tmp34067 : tmp34073;
  assign tmp34089 = ~(s1 ? tmp34090 : 0);
  assign tmp34083 = ~(s2 ? tmp34084 : tmp34089);
  assign tmp34069 = ~(s3 ? tmp34070 : tmp34083);
  assign tmp34040 = s4 ? tmp34041 : tmp34069;
  assign tmp33988 = s5 ? tmp33989 : tmp34040;
  assign tmp33914 = s6 ? tmp33915 : tmp33988;
  assign tmp34096 = l2 ? tmp33943 : tmp33921;
  assign tmp34095 = l1 ? tmp34096 : tmp33922;
  assign tmp34099 = l2 ? tmp33938 : tmp33921;
  assign tmp34098 = l1 ? tmp34099 : tmp33922;
  assign tmp34097 = s0 ? tmp33926 : tmp34098;
  assign tmp34094 = s1 ? tmp34095 : tmp34097;
  assign tmp34103 = l1 ? tmp34050 : tmp33939;
  assign tmp34105 = l2 ? tmp33942 : tmp33921;
  assign tmp34104 = ~(l1 ? tmp34105 : tmp33941);
  assign tmp34102 = s0 ? tmp34103 : tmp34104;
  assign tmp34108 = l2 ? tmp33932 : tmp33942;
  assign tmp34107 = l1 ? tmp34108 : tmp33947;
  assign tmp34106 = s0 ? tmp34107 : tmp34104;
  assign tmp34101 = s1 ? tmp34102 : tmp34106;
  assign tmp34110 = s0 ? tmp34107 : tmp33952;
  assign tmp34112 = l1 ? tmp34105 : tmp33941;
  assign tmp34113 = l1 ? tmp34105 : tmp33922;
  assign tmp34111 = ~(s0 ? tmp34112 : tmp34113);
  assign tmp34109 = s1 ? tmp34110 : tmp34111;
  assign tmp34100 = ~(s2 ? tmp34101 : tmp34109);
  assign tmp34093 = s3 ? tmp34094 : tmp34100;
  assign tmp34118 = l1 ? tmp34050 : tmp33947;
  assign tmp34117 = s0 ? tmp34118 : tmp33960;
  assign tmp34119 = ~(s0 ? tmp34113 : tmp34112);
  assign tmp34116 = s1 ? tmp34117 : tmp34119;
  assign tmp34121 = s0 ? tmp34095 : tmp33964;
  assign tmp34120 = ~(s1 ? tmp34121 : tmp33966);
  assign tmp34115 = s2 ? tmp34116 : tmp34120;
  assign tmp34123 = s1 ? tmp33926 : tmp33977;
  assign tmp34127 = l2 ? tmp33923 : tmp33920;
  assign tmp34126 = ~(l1 ? tmp34127 : tmp33983);
  assign tmp34125 = s0 ? tmp34112 : tmp34126;
  assign tmp34129 = l1 ? tmp33978 : tmp33987;
  assign tmp34128 = s0 ? tmp34129 : tmp34112;
  assign tmp34124 = s1 ? tmp34125 : tmp34128;
  assign tmp34122 = ~(s2 ? tmp34123 : tmp34124);
  assign tmp34114 = ~(s3 ? tmp34115 : tmp34122);
  assign tmp34092 = s4 ? tmp34093 : tmp34114;
  assign tmp34135 = s0 ? tmp34098 : 0;
  assign tmp34136 = ~(l1 ? tmp34050 : tmp33939);
  assign tmp34134 = s1 ? tmp34135 : tmp34136;
  assign tmp34138 = l1 ? tmp34068 : tmp33939;
  assign tmp34140 = l1 ? tmp34127 : tmp33983;
  assign tmp34139 = s0 ? tmp34140 : tmp34001;
  assign tmp34137 = ~(s1 ? tmp34138 : tmp34139);
  assign tmp34133 = s2 ? tmp34134 : tmp34137;
  assign tmp34144 = l2 ? tmp33942 : tmp33938;
  assign tmp34143 = ~(l1 ? tmp34144 : tmp34010);
  assign tmp34142 = s1 ? tmp34107 : tmp34143;
  assign tmp34146 = s0 ? tmp34129 : tmp34014;
  assign tmp34148 = l1 ? tmp34105 : tmp34010;
  assign tmp34149 = l1 ? tmp34144 : tmp33987;
  assign tmp34147 = s0 ? tmp34148 : tmp34149;
  assign tmp34145 = ~(s1 ? tmp34146 : tmp34147);
  assign tmp34141 = ~(s2 ? tmp34142 : tmp34145);
  assign tmp34132 = s3 ? tmp34133 : tmp34141;
  assign tmp34153 = s0 ? tmp33977 : tmp34148;
  assign tmp34152 = s1 ? tmp34153 : tmp34022;
  assign tmp34155 = s0 ? tmp34103 : tmp33952;
  assign tmp34154 = ~(s1 ? tmp33952 : tmp34155);
  assign tmp34151 = s2 ? tmp34152 : tmp34154;
  assign tmp34159 = l1 ? tmp34108 : tmp34034;
  assign tmp34158 = s0 ? tmp34103 : tmp34159;
  assign tmp34160 = ~(l1 ? tmp34144 : tmp33932);
  assign tmp34157 = s1 ? tmp34158 : tmp34160;
  assign tmp34161 = ~(s1 ? tmp34014 : tmp33977);
  assign tmp34156 = ~(s2 ? tmp34157 : tmp34161);
  assign tmp34150 = s3 ? tmp34151 : tmp34156;
  assign tmp34131 = s4 ? tmp34132 : tmp34150;
  assign tmp34167 = l1 ? tmp34144 : tmp34010;
  assign tmp34166 = s0 ? tmp34167 : tmp34045;
  assign tmp34168 = l1 ? 1 : tmp34024;
  assign tmp34165 = s1 ? tmp34166 : tmp34168;
  assign tmp34169 = ~(s1 ? tmp34103 : tmp34027);
  assign tmp34164 = s2 ? tmp34165 : tmp34169;
  assign tmp34171 = s1 ? tmp34061 : 1;
  assign tmp34172 = ~(s1 ? tmp34046 : tmp34103);
  assign tmp34170 = s2 ? tmp34171 : tmp34172;
  assign tmp34163 = s3 ? tmp34164 : tmp34170;
  assign tmp34175 = s1 ? tmp34061 : tmp34129;
  assign tmp34176 = ~(l1 ? tmp34068 : tmp33939);
  assign tmp34174 = s2 ? tmp34175 : tmp34176;
  assign tmp34178 = ~(l1 ? tmp34068 : tmp34034);
  assign tmp34177 = s1 ? tmp34061 : tmp34178;
  assign tmp34173 = s3 ? tmp34174 : tmp34177;
  assign tmp34162 = s4 ? tmp34163 : tmp34173;
  assign tmp34130 = s5 ? tmp34131 : tmp34162;
  assign tmp34091 = s6 ? tmp34092 : tmp34130;
  assign tmp33913 = s7 ? tmp33914 : tmp34091;
  assign tmp34185 = l1 ? tmp33927 : tmp33922;
  assign tmp34184 = s0 ? tmp33926 : tmp34185;
  assign tmp34183 = s1 ? tmp34113 : tmp34184;
  assign tmp34189 = l1 ? tmp34024 : tmp33939;
  assign tmp34188 = s0 ? tmp34189 : tmp34104;
  assign tmp34192 = l2 ? tmp33923 : tmp33942;
  assign tmp34191 = l1 ? tmp34192 : tmp33947;
  assign tmp34190 = s0 ? tmp34191 : tmp34104;
  assign tmp34187 = s1 ? tmp34188 : tmp34190;
  assign tmp34194 = s0 ? tmp34191 : tmp33952;
  assign tmp34193 = s1 ? tmp34194 : tmp34111;
  assign tmp34186 = ~(s2 ? tmp34187 : tmp34193);
  assign tmp34182 = s3 ? tmp34183 : tmp34186;
  assign tmp34199 = l1 ? tmp34024 : tmp33947;
  assign tmp34198 = s0 ? tmp34199 : tmp33960;
  assign tmp34197 = s1 ? tmp34198 : tmp34119;
  assign tmp34201 = s0 ? tmp34113 : tmp33964;
  assign tmp34200 = ~(s1 ? tmp34201 : tmp33966);
  assign tmp34196 = s2 ? tmp34197 : tmp34200;
  assign tmp34195 = ~(s3 ? tmp34196 : tmp34122);
  assign tmp34181 = s4 ? tmp34182 : tmp34195;
  assign tmp34207 = s0 ? tmp34185 : 0;
  assign tmp34208 = ~(l1 ? tmp34024 : tmp33939);
  assign tmp34206 = s1 ? tmp34207 : tmp34208;
  assign tmp34210 = l1 ? tmp34127 : tmp33939;
  assign tmp34209 = ~(s1 ? tmp34210 : tmp34139);
  assign tmp34205 = s2 ? tmp34206 : tmp34209;
  assign tmp34212 = s1 ? tmp34191 : tmp34143;
  assign tmp34211 = ~(s2 ? tmp34212 : tmp34145);
  assign tmp34204 = s3 ? tmp34205 : tmp34211;
  assign tmp34214 = s2 ? tmp34152 : tmp34208;
  assign tmp34218 = l1 ? tmp34192 : tmp34034;
  assign tmp34217 = s0 ? tmp34103 : tmp34218;
  assign tmp34216 = s1 ? tmp34217 : tmp34160;
  assign tmp34215 = ~(s2 ? tmp34216 : tmp34161);
  assign tmp34213 = s3 ? tmp34214 : tmp34215;
  assign tmp34203 = s4 ? tmp34204 : tmp34213;
  assign tmp34202 = s5 ? tmp34203 : tmp34162;
  assign tmp34180 = s6 ? tmp34181 : tmp34202;
  assign tmp34179 = s7 ? tmp33914 : tmp34180;
  assign tmp33912 = s8 ? tmp33913 : tmp34179;
  assign tmp34227 = ~(l3 ? tmp33920 : 1);
  assign tmp34226 = l2 ? tmp33923 : tmp34227;
  assign tmp34225 = l1 ? tmp34096 : tmp34226;
  assign tmp34229 = l1 ? tmp34099 : tmp33928;
  assign tmp34230 = l1 ? tmp34099 : tmp34226;
  assign tmp34228 = s0 ? tmp34229 : tmp34230;
  assign tmp34224 = s1 ? tmp34225 : tmp34228;
  assign tmp34234 = l1 ? tmp34050 : 1;
  assign tmp34235 = ~(l1 ? tmp34096 : tmp34227);
  assign tmp34233 = s0 ? tmp34234 : tmp34235;
  assign tmp34237 = l1 ? tmp34108 : tmp33973;
  assign tmp34236 = s0 ? tmp34237 : tmp34235;
  assign tmp34232 = s1 ? tmp34233 : tmp34236;
  assign tmp34239 = s0 ? tmp34237 : 1;
  assign tmp34241 = l1 ? tmp34096 : tmp34227;
  assign tmp34240 = ~(s0 ? tmp34241 : tmp34225);
  assign tmp34238 = s1 ? tmp34239 : tmp34240;
  assign tmp34231 = ~(s2 ? tmp34232 : tmp34238);
  assign tmp34223 = s3 ? tmp34224 : tmp34231;
  assign tmp34246 = l1 ? tmp34050 : tmp33973;
  assign tmp34247 = ~(l1 ? tmp34099 : tmp33929);
  assign tmp34245 = s0 ? tmp34246 : tmp34247;
  assign tmp34248 = ~(s0 ? tmp34225 : tmp34241);
  assign tmp34244 = s1 ? tmp34245 : tmp34248;
  assign tmp34252 = l2 ? tmp33938 : tmp33929;
  assign tmp34251 = l1 ? tmp34252 : tmp33964;
  assign tmp34250 = s0 ? tmp34225 : tmp34251;
  assign tmp34253 = l1 ? tmp34099 : tmp33967;
  assign tmp34249 = ~(s1 ? tmp34250 : tmp34253);
  assign tmp34243 = s2 ? tmp34244 : tmp34249;
  assign tmp34255 = s1 ? tmp34229 : tmp33977;
  assign tmp34258 = ~(l1 ? tmp34068 : tmp33942);
  assign tmp34257 = s0 ? tmp34241 : tmp34258;
  assign tmp34259 = s0 ? tmp34129 : tmp34241;
  assign tmp34256 = s1 ? tmp34257 : tmp34259;
  assign tmp34254 = ~(s2 ? tmp34255 : tmp34256);
  assign tmp34242 = ~(s3 ? tmp34243 : tmp34254);
  assign tmp34222 = s4 ? tmp34223 : tmp34242;
  assign tmp34265 = s0 ? tmp34230 : 0;
  assign tmp34266 = ~(l1 ? tmp34050 : 1);
  assign tmp34264 = s1 ? tmp34265 : tmp34266;
  assign tmp34268 = l1 ? tmp34068 : 1;
  assign tmp34270 = l1 ? tmp34068 : tmp33942;
  assign tmp34271 = ~(l1 ? tmp33937 : tmp34002);
  assign tmp34269 = s0 ? tmp34270 : tmp34271;
  assign tmp34267 = ~(s1 ? tmp34268 : tmp34269);
  assign tmp34263 = s2 ? tmp34264 : tmp34267;
  assign tmp34276 = ~(l3 ? 1 : 0);
  assign tmp34275 = ~(l2 ? tmp33942 : tmp34276);
  assign tmp34274 = ~(l1 ? tmp34144 : tmp34275);
  assign tmp34273 = s1 ? tmp34237 : tmp34274;
  assign tmp34279 = l1 ? tmp34096 : tmp34010;
  assign tmp34281 = l2 ? tmp33943 : tmp33938;
  assign tmp34280 = l1 ? tmp34281 : tmp33987;
  assign tmp34278 = s0 ? tmp34279 : tmp34280;
  assign tmp34277 = ~(s1 ? tmp34146 : tmp34278);
  assign tmp34272 = ~(s2 ? tmp34273 : tmp34277);
  assign tmp34262 = s3 ? tmp34263 : tmp34272;
  assign tmp34286 = l1 ? tmp34096 : tmp34275;
  assign tmp34285 = s0 ? tmp33977 : tmp34286;
  assign tmp34288 = ~(l1 ? tmp33938 : tmp34024);
  assign tmp34287 = ~(s0 ? 1 : tmp34288);
  assign tmp34284 = s1 ? tmp34285 : tmp34287;
  assign tmp34283 = s2 ? tmp34284 : tmp34266;
  assign tmp34292 = l1 ? tmp34108 : tmp34046;
  assign tmp34291 = s0 ? tmp34234 : tmp34292;
  assign tmp34290 = s1 ? tmp34291 : tmp34160;
  assign tmp34289 = ~(s2 ? tmp34290 : tmp34161);
  assign tmp34282 = s3 ? tmp34283 : tmp34289;
  assign tmp34261 = s4 ? tmp34262 : tmp34282;
  assign tmp34298 = l1 ? tmp34144 : tmp34275;
  assign tmp34297 = s0 ? tmp34298 : tmp34045;
  assign tmp34296 = s1 ? tmp34297 : tmp34168;
  assign tmp34299 = ~(s1 ? tmp34234 : tmp34027);
  assign tmp34295 = s2 ? tmp34296 : tmp34299;
  assign tmp34301 = ~(s1 ? tmp34046 : tmp34234);
  assign tmp34300 = s2 ? tmp34171 : tmp34301;
  assign tmp34294 = s3 ? tmp34295 : tmp34300;
  assign tmp34304 = ~(l1 ? tmp34068 : 1);
  assign tmp34303 = s2 ? tmp34175 : tmp34304;
  assign tmp34306 = ~(l1 ? tmp34068 : tmp34046);
  assign tmp34305 = s1 ? tmp34061 : tmp34306;
  assign tmp34302 = s3 ? tmp34303 : tmp34305;
  assign tmp34293 = s4 ? tmp34294 : tmp34302;
  assign tmp34260 = s5 ? tmp34261 : tmp34293;
  assign tmp34221 = s6 ? tmp34222 : tmp34260;
  assign tmp34220 = s7 ? tmp33914 : tmp34221;
  assign tmp34219 = s8 ? tmp34179 : tmp34220;
  assign tmp33911 = s9 ? tmp33912 : tmp34219;
  assign tmp34314 = s0 ? tmp34229 : tmp34098;
  assign tmp34313 = s1 ? tmp34095 : tmp34314;
  assign tmp34318 = ~(l1 ? tmp34096 : tmp33941);
  assign tmp34317 = s0 ? tmp34103 : tmp34318;
  assign tmp34319 = s0 ? tmp34107 : tmp34318;
  assign tmp34316 = s1 ? tmp34317 : tmp34319;
  assign tmp34321 = s0 ? tmp34107 : 1;
  assign tmp34323 = l1 ? tmp34096 : tmp33941;
  assign tmp34322 = ~(s0 ? tmp34323 : tmp34095);
  assign tmp34320 = s1 ? tmp34321 : tmp34322;
  assign tmp34315 = ~(s2 ? tmp34316 : tmp34320);
  assign tmp34312 = s3 ? tmp34313 : tmp34315;
  assign tmp34327 = s0 ? tmp34118 : tmp34247;
  assign tmp34328 = ~(s0 ? tmp34095 : tmp34323);
  assign tmp34326 = s1 ? tmp34327 : tmp34328;
  assign tmp34330 = s0 ? tmp34095 : tmp34251;
  assign tmp34329 = ~(s1 ? tmp34330 : tmp34253);
  assign tmp34325 = s2 ? tmp34326 : tmp34329;
  assign tmp34334 = ~(l1 ? tmp34068 : tmp33983);
  assign tmp34333 = s0 ? tmp34323 : tmp34334;
  assign tmp34335 = s0 ? tmp34129 : tmp34323;
  assign tmp34332 = s1 ? tmp34333 : tmp34335;
  assign tmp34331 = ~(s2 ? tmp34255 : tmp34332);
  assign tmp34324 = ~(s3 ? tmp34325 : tmp34331);
  assign tmp34311 = s4 ? tmp34312 : tmp34324;
  assign tmp34342 = l1 ? tmp34068 : tmp33983;
  assign tmp34341 = s0 ? tmp34342 : tmp34271;
  assign tmp34340 = ~(s1 ? tmp34138 : tmp34341);
  assign tmp34339 = s2 ? tmp34134 : tmp34340;
  assign tmp34343 = ~(s2 ? tmp34142 : tmp34277);
  assign tmp34338 = s3 ? tmp34339 : tmp34343;
  assign tmp34347 = s0 ? tmp33977 : tmp34279;
  assign tmp34346 = s1 ? tmp34347 : tmp34287;
  assign tmp34345 = s2 ? tmp34346 : tmp34136;
  assign tmp34344 = s3 ? tmp34345 : tmp34156;
  assign tmp34337 = s4 ? tmp34338 : tmp34344;
  assign tmp34336 = s5 ? tmp34337 : tmp34162;
  assign tmp34310 = s6 ? tmp34311 : tmp34336;
  assign tmp34309 = s7 ? tmp33914 : tmp34310;
  assign tmp34308 = s8 ? tmp34309 : tmp33914;
  assign tmp34355 = ~(s1 ? tmp33952 : tmp34103);
  assign tmp34354 = s2 ? tmp34152 : tmp34355;
  assign tmp34353 = s3 ? tmp34354 : tmp34156;
  assign tmp34352 = s4 ? tmp34132 : tmp34353;
  assign tmp34351 = s5 ? tmp34352 : tmp34162;
  assign tmp34350 = s6 ? tmp34092 : tmp34351;
  assign tmp34349 = s7 ? tmp34350 : tmp34221;
  assign tmp34356 = s7 ? tmp34180 : tmp34310;
  assign tmp34348 = s8 ? tmp34349 : tmp34356;
  assign tmp34307 = s9 ? tmp34308 : tmp34348;
  assign tmp33910 = s10 ? tmp33911 : tmp34307;
  assign tmp34360 = s7 ? tmp34091 : tmp34221;
  assign tmp34359 = s8 ? tmp34360 : tmp34356;
  assign tmp34358 = s9 ? tmp34308 : tmp34359;
  assign tmp34357 = s10 ? tmp33911 : tmp34358;
  assign tmp33909 = s11 ? tmp33910 : tmp34357;
  assign tmp34373 = ~(l1 ? tmp34105 : tmp34227);
  assign tmp34372 = s0 ? tmp34234 : tmp34373;
  assign tmp34374 = s0 ? tmp34237 : tmp34373;
  assign tmp34371 = s1 ? tmp34372 : tmp34374;
  assign tmp34376 = s0 ? tmp34237 : tmp33952;
  assign tmp34378 = l1 ? tmp34105 : tmp34227;
  assign tmp34377 = ~(s0 ? tmp34378 : tmp34225);
  assign tmp34375 = s1 ? tmp34376 : tmp34377;
  assign tmp34370 = ~(s2 ? tmp34371 : tmp34375);
  assign tmp34369 = s3 ? tmp34224 : tmp34370;
  assign tmp34382 = ~(s0 ? tmp34225 : tmp34378);
  assign tmp34381 = s1 ? tmp34245 : tmp34382;
  assign tmp34384 = s0 ? tmp34225 : tmp33964;
  assign tmp34385 = s0 ? tmp34253 : tmp33968;
  assign tmp34383 = ~(s1 ? tmp34384 : tmp34385);
  assign tmp34380 = s2 ? tmp34381 : tmp34383;
  assign tmp34387 = s1 ? tmp34229 : tmp33976;
  assign tmp34390 = ~(l1 ? tmp34127 : tmp33942);
  assign tmp34389 = s0 ? tmp34378 : tmp34390;
  assign tmp34391 = s0 ? tmp34129 : tmp34378;
  assign tmp34388 = s1 ? tmp34389 : tmp34391;
  assign tmp34386 = ~(s2 ? tmp34387 : tmp34388);
  assign tmp34379 = ~(s3 ? tmp34380 : tmp34386);
  assign tmp34368 = s4 ? tmp34369 : tmp34379;
  assign tmp34397 = ~(s0 ? tmp33995 : tmp34234);
  assign tmp34396 = s1 ? tmp34265 : tmp34397;
  assign tmp34399 = s0 ? tmp33995 : tmp34268;
  assign tmp34401 = l1 ? tmp34127 : tmp33942;
  assign tmp34400 = s0 ? tmp34401 : tmp34001;
  assign tmp34398 = ~(s1 ? tmp34399 : tmp34400);
  assign tmp34395 = s2 ? tmp34396 : tmp34398;
  assign tmp34405 = ~(l1 ? tmp34108 : tmp33973);
  assign tmp34404 = s0 ? 1 : tmp34405;
  assign tmp34406 = s0 ? 1 : tmp34298;
  assign tmp34403 = s1 ? tmp34404 : tmp34406;
  assign tmp34409 = l1 ? tmp34105 : tmp34275;
  assign tmp34410 = l1 ? tmp34144 : tmp33923;
  assign tmp34408 = s0 ? tmp34409 : tmp34410;
  assign tmp34407 = s1 ? tmp34146 : tmp34408;
  assign tmp34402 = s2 ? tmp34403 : tmp34407;
  assign tmp34394 = s3 ? tmp34395 : tmp34402;
  assign tmp34415 = l2 ? tmp33932 : tmp33923;
  assign tmp34414 = ~(l1 ? tmp34144 : tmp34415);
  assign tmp34413 = s1 ? tmp34291 : tmp34414;
  assign tmp34412 = ~(s2 ? tmp34413 : tmp34161);
  assign tmp34411 = s3 ? tmp34283 : tmp34412;
  assign tmp34393 = s4 ? tmp34394 : tmp34411;
  assign tmp34419 = ~(s1 ? tmp34234 : tmp34082);
  assign tmp34418 = s2 ? tmp34296 : tmp34419;
  assign tmp34417 = s3 ? tmp34418 : tmp34300;
  assign tmp34416 = s4 ? tmp34417 : tmp34302;
  assign tmp34392 = s5 ? tmp34393 : tmp34416;
  assign tmp34367 = s6 ? tmp34368 : tmp34392;
  assign tmp34366 = s7 ? tmp33914 : tmp34367;
  assign tmp34425 = l1 ? tmp34105 : tmp34226;
  assign tmp34427 = l1 ? tmp33927 : tmp34226;
  assign tmp34426 = s0 ? tmp33926 : tmp34427;
  assign tmp34424 = s1 ? tmp34425 : tmp34426;
  assign tmp34431 = l1 ? tmp34024 : 1;
  assign tmp34430 = s0 ? tmp34431 : tmp34373;
  assign tmp34433 = l1 ? tmp34192 : tmp33973;
  assign tmp34432 = s0 ? tmp34433 : tmp34373;
  assign tmp34429 = s1 ? tmp34430 : tmp34432;
  assign tmp34435 = s0 ? tmp34433 : tmp33952;
  assign tmp34436 = ~(s0 ? tmp34378 : tmp34425);
  assign tmp34434 = s1 ? tmp34435 : tmp34436;
  assign tmp34428 = ~(s2 ? tmp34429 : tmp34434);
  assign tmp34423 = s3 ? tmp34424 : tmp34428;
  assign tmp34441 = l1 ? tmp34024 : tmp33973;
  assign tmp34440 = s0 ? tmp34441 : tmp33960;
  assign tmp34442 = ~(s0 ? tmp34425 : tmp34378);
  assign tmp34439 = s1 ? tmp34440 : tmp34442;
  assign tmp34444 = s0 ? tmp34425 : tmp33964;
  assign tmp34443 = ~(s1 ? tmp34444 : tmp33966);
  assign tmp34438 = s2 ? tmp34439 : tmp34443;
  assign tmp34445 = ~(s2 ? tmp34123 : tmp34388);
  assign tmp34437 = ~(s3 ? tmp34438 : tmp34445);
  assign tmp34422 = s4 ? tmp34423 : tmp34437;
  assign tmp34451 = s0 ? tmp34427 : 0;
  assign tmp34452 = ~(s0 ? tmp33995 : tmp34431);
  assign tmp34450 = s1 ? tmp34451 : tmp34452;
  assign tmp34455 = l1 ? tmp34127 : 1;
  assign tmp34454 = s0 ? tmp33995 : tmp34455;
  assign tmp34453 = ~(s1 ? tmp34454 : tmp34400);
  assign tmp34449 = s2 ? tmp34450 : tmp34453;
  assign tmp34457 = s1 ? tmp34433 : tmp34274;
  assign tmp34458 = ~(s1 ? tmp34146 : tmp34408);
  assign tmp34456 = ~(s2 ? tmp34457 : tmp34458);
  assign tmp34448 = s3 ? tmp34449 : tmp34456;
  assign tmp34462 = s0 ? tmp33977 : tmp34409;
  assign tmp34461 = s1 ? tmp34462 : tmp34022;
  assign tmp34463 = ~(l1 ? tmp34024 : 1);
  assign tmp34460 = s2 ? tmp34461 : tmp34463;
  assign tmp34467 = l1 ? tmp34192 : tmp34046;
  assign tmp34466 = s0 ? tmp34234 : tmp34467;
  assign tmp34465 = s1 ? tmp34466 : tmp34414;
  assign tmp34464 = ~(s2 ? tmp34465 : tmp34161);
  assign tmp34459 = s3 ? tmp34460 : tmp34464;
  assign tmp34447 = s4 ? tmp34448 : tmp34459;
  assign tmp34446 = s5 ? tmp34447 : tmp34416;
  assign tmp34421 = s6 ? tmp34422 : tmp34446;
  assign tmp34420 = s7 ? tmp33914 : tmp34421;
  assign tmp34365 = s8 ? tmp34366 : tmp34420;
  assign tmp34473 = s1 ? tmp34095 : tmp34228;
  assign tmp34472 = s3 ? tmp34473 : tmp34315;
  assign tmp34476 = s1 ? tmp34245 : tmp34328;
  assign tmp34475 = s2 ? tmp34476 : tmp34329;
  assign tmp34474 = ~(s3 ? tmp34475 : tmp34331);
  assign tmp34471 = s4 ? tmp34472 : tmp34474;
  assign tmp34482 = ~(s0 ? tmp33995 : tmp34103);
  assign tmp34481 = s1 ? tmp34265 : tmp34482;
  assign tmp34483 = ~(s1 ? tmp34399 : tmp34341);
  assign tmp34480 = s2 ? tmp34481 : tmp34483;
  assign tmp34485 = s1 ? tmp34107 : tmp34274;
  assign tmp34488 = l1 ? tmp34281 : tmp33923;
  assign tmp34487 = s0 ? tmp34286 : tmp34488;
  assign tmp34486 = ~(s1 ? tmp34146 : tmp34487);
  assign tmp34484 = ~(s2 ? tmp34485 : tmp34486);
  assign tmp34479 = s3 ? tmp34480 : tmp34484;
  assign tmp34478 = s4 ? tmp34479 : tmp34411;
  assign tmp34477 = s5 ? tmp34478 : tmp34416;
  assign tmp34470 = s6 ? tmp34471 : tmp34477;
  assign tmp34469 = s7 ? tmp33914 : tmp34470;
  assign tmp34468 = s8 ? tmp34420 : tmp34469;
  assign tmp34364 = s9 ? tmp34365 : tmp34468;
  assign tmp34497 = ~(s1 ? tmp34399 : tmp34269);
  assign tmp34496 = s2 ? tmp34396 : tmp34497;
  assign tmp34498 = ~(s2 ? tmp34273 : tmp34486);
  assign tmp34495 = s3 ? tmp34496 : tmp34498;
  assign tmp34494 = s4 ? tmp34495 : tmp34411;
  assign tmp34493 = s5 ? tmp34494 : tmp34416;
  assign tmp34492 = s6 ? tmp34222 : tmp34493;
  assign tmp34491 = s7 ? tmp33914 : tmp34492;
  assign tmp34490 = s8 ? tmp34491 : tmp33914;
  assign tmp34504 = ~(s2 ? tmp34255 : tmp34388);
  assign tmp34503 = ~(s3 ? tmp34380 : tmp34504);
  assign tmp34502 = s4 ? tmp34369 : tmp34503;
  assign tmp34509 = ~(s1 ? tmp34268 : tmp34400);
  assign tmp34508 = s2 ? tmp34396 : tmp34509;
  assign tmp34511 = s1 ? tmp34404 : tmp34298;
  assign tmp34510 = s2 ? tmp34511 : tmp34407;
  assign tmp34507 = s3 ? tmp34508 : tmp34510;
  assign tmp34506 = s4 ? tmp34507 : tmp34411;
  assign tmp34505 = s5 ? tmp34506 : tmp34416;
  assign tmp34501 = s6 ? tmp34502 : tmp34505;
  assign tmp34517 = ~(s1 ? tmp34268 : tmp34341);
  assign tmp34516 = s2 ? tmp34481 : tmp34517;
  assign tmp34515 = s3 ? tmp34516 : tmp34484;
  assign tmp34514 = s4 ? tmp34515 : tmp34411;
  assign tmp34513 = s5 ? tmp34514 : tmp34416;
  assign tmp34512 = s6 ? tmp34471 : tmp34513;
  assign tmp34500 = s7 ? tmp34501 : tmp34512;
  assign tmp34524 = ~(s1 ? tmp34455 : tmp34400);
  assign tmp34523 = s2 ? tmp34450 : tmp34524;
  assign tmp34522 = s3 ? tmp34523 : tmp34456;
  assign tmp34521 = s4 ? tmp34522 : tmp34459;
  assign tmp34520 = s5 ? tmp34521 : tmp34416;
  assign tmp34519 = s6 ? tmp34422 : tmp34520;
  assign tmp34529 = s2 ? tmp34396 : tmp34267;
  assign tmp34528 = s3 ? tmp34529 : tmp34498;
  assign tmp34527 = s4 ? tmp34528 : tmp34411;
  assign tmp34526 = s5 ? tmp34527 : tmp34416;
  assign tmp34525 = s6 ? tmp34222 : tmp34526;
  assign tmp34518 = s7 ? tmp34519 : tmp34525;
  assign tmp34499 = s8 ? tmp34500 : tmp34518;
  assign tmp34489 = s9 ? tmp34490 : tmp34499;
  assign tmp34363 = s10 ? tmp34364 : tmp34489;
  assign tmp34533 = s7 ? tmp34367 : tmp34470;
  assign tmp34534 = s7 ? tmp34421 : tmp34492;
  assign tmp34532 = s8 ? tmp34533 : tmp34534;
  assign tmp34531 = s9 ? tmp34490 : tmp34532;
  assign tmp34530 = s10 ? tmp34364 : tmp34531;
  assign tmp34362 = s11 ? tmp34363 : tmp34530;
  assign tmp34545 = l1 ? tmp34099 : tmp33975;
  assign tmp34546 = l1 ? tmp34099 : tmp34227;
  assign tmp34544 = s0 ? tmp34545 : tmp34546;
  assign tmp34543 = s1 ? tmp34241 : tmp34544;
  assign tmp34550 = l1 ? tmp34108 : 1;
  assign tmp34549 = s0 ? tmp34550 : tmp34235;
  assign tmp34548 = s1 ? tmp34233 : tmp34549;
  assign tmp34552 = s0 ? tmp34550 : tmp33952;
  assign tmp34551 = s1 ? tmp34552 : tmp34235;
  assign tmp34547 = ~(s2 ? tmp34548 : tmp34551);
  assign tmp34542 = s3 ? tmp34543 : tmp34547;
  assign tmp34556 = s0 ? tmp34234 : tmp34247;
  assign tmp34555 = s1 ? tmp34556 : tmp34235;
  assign tmp34558 = s0 ? tmp34241 : tmp33964;
  assign tmp34557 = ~(s1 ? tmp34558 : tmp34385);
  assign tmp34554 = s2 ? tmp34555 : tmp34557;
  assign tmp34560 = s1 ? tmp34545 : tmp33976;
  assign tmp34559 = ~(s2 ? tmp34560 : tmp34256);
  assign tmp34553 = ~(s3 ? tmp34554 : tmp34559);
  assign tmp34541 = s4 ? tmp34542 : tmp34553;
  assign tmp34566 = s0 ? tmp34546 : 0;
  assign tmp34565 = s1 ? tmp34566 : tmp34266;
  assign tmp34564 = s2 ? tmp34565 : tmp34267;
  assign tmp34568 = s1 ? tmp34550 : tmp34274;
  assign tmp34567 = ~(s2 ? tmp34568 : tmp34486);
  assign tmp34563 = s3 ? tmp34564 : tmp34567;
  assign tmp34562 = s4 ? tmp34563 : tmp34411;
  assign tmp34561 = s5 ? tmp34562 : tmp34416;
  assign tmp34540 = s6 ? tmp34541 : tmp34561;
  assign tmp34539 = s7 ? tmp33914 : tmp34540;
  assign tmp34575 = l1 ? tmp33927 : tmp34227;
  assign tmp34574 = s0 ? tmp33974 : tmp34575;
  assign tmp34573 = s1 ? tmp34378 : tmp34574;
  assign tmp34579 = l1 ? tmp34192 : 1;
  assign tmp34578 = s0 ? tmp34579 : tmp34373;
  assign tmp34577 = s1 ? tmp34430 : tmp34578;
  assign tmp34581 = s0 ? tmp34579 : tmp33952;
  assign tmp34580 = s1 ? tmp34581 : tmp34373;
  assign tmp34576 = ~(s2 ? tmp34577 : tmp34580);
  assign tmp34572 = s3 ? tmp34573 : tmp34576;
  assign tmp34585 = s0 ? tmp34431 : tmp33960;
  assign tmp34584 = s1 ? tmp34585 : tmp34373;
  assign tmp34587 = s0 ? tmp34378 : tmp33964;
  assign tmp34586 = ~(s1 ? tmp34587 : tmp33966);
  assign tmp34583 = s2 ? tmp34584 : tmp34586;
  assign tmp34589 = s1 ? tmp33974 : tmp33977;
  assign tmp34588 = ~(s2 ? tmp34589 : tmp34388);
  assign tmp34582 = ~(s3 ? tmp34583 : tmp34588);
  assign tmp34571 = s4 ? tmp34572 : tmp34582;
  assign tmp34595 = s0 ? tmp34575 : 0;
  assign tmp34594 = s1 ? tmp34595 : tmp34463;
  assign tmp34593 = s2 ? tmp34594 : tmp34524;
  assign tmp34597 = s1 ? tmp34579 : tmp34274;
  assign tmp34596 = ~(s2 ? tmp34597 : tmp34458);
  assign tmp34592 = s3 ? tmp34593 : tmp34596;
  assign tmp34591 = s4 ? tmp34592 : tmp34459;
  assign tmp34590 = s5 ? tmp34591 : tmp34416;
  assign tmp34570 = s6 ? tmp34571 : tmp34590;
  assign tmp34569 = s7 ? tmp33914 : tmp34570;
  assign tmp34538 = s8 ? tmp34539 : tmp34569;
  assign tmp34603 = s1 ? tmp34323 : tmp34544;
  assign tmp34607 = l1 ? tmp34108 : tmp33939;
  assign tmp34606 = s0 ? tmp34607 : tmp34318;
  assign tmp34605 = s1 ? tmp34317 : tmp34606;
  assign tmp34609 = s0 ? tmp34607 : 1;
  assign tmp34608 = s1 ? tmp34609 : tmp34318;
  assign tmp34604 = ~(s2 ? tmp34605 : tmp34608);
  assign tmp34602 = s3 ? tmp34603 : tmp34604;
  assign tmp34612 = s1 ? tmp34556 : tmp34318;
  assign tmp34614 = s0 ? tmp34323 : tmp34251;
  assign tmp34613 = ~(s1 ? tmp34614 : tmp34253);
  assign tmp34611 = s2 ? tmp34612 : tmp34613;
  assign tmp34616 = s1 ? tmp34545 : tmp33977;
  assign tmp34615 = ~(s2 ? tmp34616 : tmp34332);
  assign tmp34610 = ~(s3 ? tmp34611 : tmp34615);
  assign tmp34601 = s4 ? tmp34602 : tmp34610;
  assign tmp34621 = s1 ? tmp34566 : tmp34136;
  assign tmp34620 = s2 ? tmp34621 : tmp34517;
  assign tmp34623 = s1 ? tmp34607 : tmp34274;
  assign tmp34622 = ~(s2 ? tmp34623 : tmp34486);
  assign tmp34619 = s3 ? tmp34620 : tmp34622;
  assign tmp34618 = s4 ? tmp34619 : tmp34411;
  assign tmp34617 = s5 ? tmp34618 : tmp34416;
  assign tmp34600 = s6 ? tmp34601 : tmp34617;
  assign tmp34599 = s7 ? tmp33914 : tmp34600;
  assign tmp34598 = s8 ? tmp34569 : tmp34599;
  assign tmp34537 = s9 ? tmp34538 : tmp34598;
  assign tmp34632 = s0 ? tmp34550 : 1;
  assign tmp34631 = s1 ? tmp34632 : tmp34235;
  assign tmp34630 = ~(s2 ? tmp34548 : tmp34631);
  assign tmp34629 = s3 ? tmp34543 : tmp34630;
  assign tmp34636 = s0 ? tmp34241 : tmp34251;
  assign tmp34635 = ~(s1 ? tmp34636 : tmp34253);
  assign tmp34634 = s2 ? tmp34555 : tmp34635;
  assign tmp34637 = ~(s2 ? tmp34616 : tmp34256);
  assign tmp34633 = ~(s3 ? tmp34634 : tmp34637);
  assign tmp34628 = s4 ? tmp34629 : tmp34633;
  assign tmp34627 = s6 ? tmp34628 : tmp34561;
  assign tmp34626 = s7 ? tmp33914 : tmp34627;
  assign tmp34625 = s8 ? tmp34626 : tmp33914;
  assign tmp34642 = ~(s3 ? tmp34554 : tmp34637);
  assign tmp34641 = s4 ? tmp34542 : tmp34642;
  assign tmp34640 = s6 ? tmp34641 : tmp34561;
  assign tmp34639 = s7 ? tmp34640 : tmp34600;
  assign tmp34643 = s7 ? tmp34570 : tmp34627;
  assign tmp34638 = s8 ? tmp34639 : tmp34643;
  assign tmp34624 = s9 ? tmp34625 : tmp34638;
  assign tmp34536 = s10 ? tmp34537 : tmp34624;
  assign tmp34647 = s7 ? tmp34540 : tmp34600;
  assign tmp34646 = s8 ? tmp34647 : tmp34643;
  assign tmp34645 = s9 ? tmp34625 : tmp34646;
  assign tmp34644 = s10 ? tmp34537 : tmp34645;
  assign tmp34535 = s11 ? tmp34536 : tmp34644;
  assign tmp34361 = s12 ? tmp34362 : tmp34535;
  assign tmp33908 = s13 ? tmp33909 : tmp34361;
  assign tmp34659 = s0 ? tmp34241 : tmp34390;
  assign tmp34658 = s1 ? tmp34659 : tmp34259;
  assign tmp34657 = ~(s2 ? tmp34255 : tmp34658);
  assign tmp34656 = ~(s3 ? tmp34243 : tmp34657);
  assign tmp34655 = s4 ? tmp34223 : tmp34656;
  assign tmp34663 = s2 ? tmp34264 : tmp34509;
  assign tmp34665 = s1 ? tmp34146 : tmp34487;
  assign tmp34664 = s2 ? tmp34403 : tmp34665;
  assign tmp34662 = s3 ? tmp34663 : tmp34664;
  assign tmp34661 = s4 ? tmp34662 : tmp34411;
  assign tmp34660 = s5 ? tmp34661 : tmp34416;
  assign tmp34654 = s6 ? tmp34655 : tmp34660;
  assign tmp34653 = s7 ? tmp33914 : tmp34654;
  assign tmp34670 = s3 ? tmp34263 : tmp34498;
  assign tmp34669 = s4 ? tmp34670 : tmp34411;
  assign tmp34668 = s5 ? tmp34669 : tmp34416;
  assign tmp34667 = s6 ? tmp34222 : tmp34668;
  assign tmp34666 = s7 ? tmp33914 : tmp34667;
  assign tmp34652 = s8 ? tmp34653 : tmp34666;
  assign tmp34677 = s2 ? tmp34284 : tmp34136;
  assign tmp34680 = s0 ? tmp34103 : tmp34292;
  assign tmp34679 = s1 ? tmp34680 : tmp34414;
  assign tmp34678 = ~(s2 ? tmp34679 : tmp34161);
  assign tmp34676 = s3 ? tmp34677 : tmp34678;
  assign tmp34675 = s4 ? tmp34338 : tmp34676;
  assign tmp34684 = ~(s1 ? tmp34103 : tmp34082);
  assign tmp34683 = s2 ? tmp34165 : tmp34684;
  assign tmp34682 = s3 ? tmp34683 : tmp34300;
  assign tmp34685 = s3 ? tmp34174 : tmp34305;
  assign tmp34681 = s4 ? tmp34682 : tmp34685;
  assign tmp34674 = s5 ? tmp34675 : tmp34681;
  assign tmp34673 = s6 ? tmp34311 : tmp34674;
  assign tmp34672 = s7 ? tmp33914 : tmp34673;
  assign tmp34671 = s8 ? tmp34666 : tmp34672;
  assign tmp34651 = s9 ? tmp34652 : tmp34671;
  assign tmp34687 = s8 ? tmp34666 : tmp33914;
  assign tmp34689 = s7 ? tmp34654 : tmp34673;
  assign tmp34688 = s8 ? tmp34689 : tmp34667;
  assign tmp34686 = s9 ? tmp34687 : tmp34688;
  assign tmp34650 = s10 ? tmp34651 : tmp34686;
  assign tmp34700 = l1 ? tmp34099 : tmp33941;
  assign tmp34699 = s0 ? tmp33974 : tmp34700;
  assign tmp34698 = s1 ? tmp34323 : tmp34699;
  assign tmp34697 = s3 ? tmp34698 : tmp34604;
  assign tmp34704 = s0 ? tmp34103 : tmp33960;
  assign tmp34703 = s1 ? tmp34704 : tmp34318;
  assign tmp34705 = ~(s1 ? tmp34614 : tmp33966);
  assign tmp34702 = s2 ? tmp34703 : tmp34705;
  assign tmp34708 = s0 ? tmp34323 : tmp34126;
  assign tmp34707 = s1 ? tmp34708 : tmp34335;
  assign tmp34706 = ~(s2 ? tmp34589 : tmp34707);
  assign tmp34701 = ~(s3 ? tmp34702 : tmp34706);
  assign tmp34696 = s4 ? tmp34697 : tmp34701;
  assign tmp34714 = s0 ? tmp34700 : 0;
  assign tmp34713 = s1 ? tmp34714 : tmp34136;
  assign tmp34716 = s0 ? tmp34140 : tmp34271;
  assign tmp34715 = ~(s1 ? tmp34138 : tmp34716);
  assign tmp34712 = s2 ? tmp34713 : tmp34715;
  assign tmp34718 = s1 ? tmp34607 : tmp34143;
  assign tmp34720 = s0 ? tmp34279 : tmp34149;
  assign tmp34719 = ~(s1 ? tmp34146 : tmp34720);
  assign tmp34717 = ~(s2 ? tmp34718 : tmp34719);
  assign tmp34711 = s3 ? tmp34712 : tmp34717;
  assign tmp34723 = s1 ? tmp34347 : tmp34022;
  assign tmp34724 = s1 ? tmp34036 : tmp34136;
  assign tmp34722 = s2 ? tmp34723 : tmp34724;
  assign tmp34728 = l1 ? tmp34144 : tmp33932;
  assign tmp34727 = ~(s0 ? tmp34036 : tmp34728);
  assign tmp34726 = s1 ? tmp34158 : tmp34727;
  assign tmp34725 = ~(s2 ? tmp34726 : tmp34161);
  assign tmp34721 = s3 ? tmp34722 : tmp34725;
  assign tmp34710 = s4 ? tmp34711 : tmp34721;
  assign tmp34709 = s5 ? tmp34710 : tmp34162;
  assign tmp34695 = s6 ? tmp34696 : tmp34709;
  assign tmp34694 = s7 ? tmp33914 : tmp34695;
  assign tmp34734 = s0 ? tmp34545 : tmp34700;
  assign tmp34733 = s1 ? tmp34323 : tmp34734;
  assign tmp34732 = s3 ? tmp34733 : tmp34604;
  assign tmp34738 = s0 ? tmp34103 : tmp34247;
  assign tmp34737 = s1 ? tmp34738 : tmp34318;
  assign tmp34736 = s2 ? tmp34737 : tmp34613;
  assign tmp34735 = ~(s3 ? tmp34736 : tmp34615);
  assign tmp34731 = s4 ? tmp34732 : tmp34735;
  assign tmp34742 = s2 ? tmp34713 : tmp34340;
  assign tmp34743 = ~(s2 ? tmp34718 : tmp34277);
  assign tmp34741 = s3 ? tmp34742 : tmp34743;
  assign tmp34740 = s4 ? tmp34741 : tmp34344;
  assign tmp34739 = s5 ? tmp34740 : tmp34162;
  assign tmp34730 = s6 ? tmp34731 : tmp34739;
  assign tmp34729 = s7 ? tmp33914 : tmp34730;
  assign tmp34693 = s8 ? tmp34694 : tmp34729;
  assign tmp34692 = s9 ? tmp34693 : tmp34729;
  assign tmp34745 = s8 ? tmp34729 : tmp33914;
  assign tmp34751 = s3 ? tmp34722 : tmp34156;
  assign tmp34750 = s4 ? tmp34711 : tmp34751;
  assign tmp34749 = s5 ? tmp34750 : tmp34162;
  assign tmp34748 = s6 ? tmp34696 : tmp34749;
  assign tmp34753 = s5 ? tmp34562 : tmp34293;
  assign tmp34752 = s6 ? tmp34628 : tmp34753;
  assign tmp34747 = s7 ? tmp34748 : tmp34752;
  assign tmp34746 = s8 ? tmp34747 : tmp34730;
  assign tmp34744 = s9 ? tmp34745 : tmp34746;
  assign tmp34691 = s10 ? tmp34692 : tmp34744;
  assign tmp34757 = s7 ? tmp34695 : tmp34752;
  assign tmp34756 = s8 ? tmp34757 : tmp34730;
  assign tmp34755 = s9 ? tmp34745 : tmp34756;
  assign tmp34754 = s10 ? tmp34692 : tmp34755;
  assign tmp34690 = s11 ? tmp34691 : tmp34754;
  assign tmp34649 = s12 ? tmp34650 : tmp34690;
  assign tmp34769 = s0 ? tmp33918 : tmp34251;
  assign tmp34768 = ~(s1 ? tmp34769 : tmp33966);
  assign tmp34767 = s2 ? tmp33957 : tmp34768;
  assign tmp34770 = ~(s2 ? tmp34123 : tmp33979);
  assign tmp34766 = ~(s3 ? tmp34767 : tmp34770);
  assign tmp34765 = s4 ? tmp33916 : tmp34766;
  assign tmp34776 = ~(l1 ? tmp33937 : tmp33939);
  assign tmp34775 = s1 ? tmp33993 : tmp34776;
  assign tmp34777 = ~(s1 ? tmp33998 : tmp33999);
  assign tmp34774 = s2 ? tmp34775 : tmp34777;
  assign tmp34780 = ~(l1 ? tmp34009 : tmp34010);
  assign tmp34779 = s1 ? tmp33945 : tmp34780;
  assign tmp34781 = ~(s1 ? tmp34013 : tmp34015);
  assign tmp34778 = ~(s2 ? tmp34779 : tmp34781);
  assign tmp34773 = s3 ? tmp34774 : tmp34778;
  assign tmp34783 = s2 ? tmp34020 : tmp34776;
  assign tmp34786 = ~(l1 ? tmp34009 : tmp33932);
  assign tmp34785 = s1 ? tmp34031 : tmp34786;
  assign tmp34784 = ~(s2 ? tmp34785 : tmp34161);
  assign tmp34782 = s3 ? tmp34783 : tmp34784;
  assign tmp34772 = s4 ? tmp34773 : tmp34782;
  assign tmp34791 = l1 ? tmp34050 : tmp34024;
  assign tmp34790 = s1 ? tmp34044 : tmp34791;
  assign tmp34793 = ~(s0 ? tmp34055 : tmp34057);
  assign tmp34792 = ~(s1 ? tmp34032 : tmp34793);
  assign tmp34789 = s2 ? tmp34790 : tmp34792;
  assign tmp34795 = ~(s1 ? tmp34046 : tmp34032);
  assign tmp34794 = s2 ? tmp34059 : tmp34795;
  assign tmp34788 = s3 ? tmp34789 : tmp34794;
  assign tmp34798 = s1 ? tmp34086 : tmp33985;
  assign tmp34799 = ~(s1 ? tmp34078 : tmp34080);
  assign tmp34797 = s2 ? tmp34798 : tmp34799;
  assign tmp34800 = s1 ? tmp34086 : tmp34088;
  assign tmp34796 = s3 ? tmp34797 : tmp34800;
  assign tmp34787 = s4 ? tmp34788 : tmp34796;
  assign tmp34771 = s5 ? tmp34772 : tmp34787;
  assign tmp34764 = s6 ? tmp34765 : tmp34771;
  assign tmp34763 = s7 ? tmp33914 : tmp34764;
  assign tmp34807 = l2 ? tmp33948 : tmp33921;
  assign tmp34806 = l1 ? tmp34807 : tmp33922;
  assign tmp34810 = l2 ? tmp33923 : tmp33921;
  assign tmp34809 = l1 ? tmp34810 : tmp33922;
  assign tmp34808 = s0 ? tmp34229 : tmp34809;
  assign tmp34805 = s1 ? tmp34806 : tmp34808;
  assign tmp34814 = ~(l1 ? tmp34807 : tmp33941);
  assign tmp34813 = s0 ? tmp34032 : tmp34814;
  assign tmp34816 = l1 ? tmp34046 : tmp33947;
  assign tmp34815 = s0 ? tmp34816 : tmp34814;
  assign tmp34812 = s1 ? tmp34813 : tmp34815;
  assign tmp34818 = s0 ? tmp34816 : 1;
  assign tmp34820 = l1 ? tmp34807 : tmp33941;
  assign tmp34819 = ~(s0 ? tmp34820 : tmp34806);
  assign tmp34817 = s1 ? tmp34818 : tmp34819;
  assign tmp34811 = ~(s2 ? tmp34812 : tmp34817);
  assign tmp34804 = s3 ? tmp34805 : tmp34811;
  assign tmp34825 = l1 ? 1 : tmp33947;
  assign tmp34824 = s0 ? tmp34825 : tmp34247;
  assign tmp34826 = ~(s0 ? tmp34806 : tmp34820);
  assign tmp34823 = s1 ? tmp34824 : tmp34826;
  assign tmp34828 = s0 ? tmp34806 : tmp34251;
  assign tmp34827 = ~(s1 ? tmp34828 : tmp34253);
  assign tmp34822 = s2 ? tmp34823 : tmp34827;
  assign tmp34832 = ~(l1 ? tmp34079 : tmp33983);
  assign tmp34831 = s0 ? tmp34820 : tmp34832;
  assign tmp34833 = s0 ? tmp33985 : tmp34820;
  assign tmp34830 = s1 ? tmp34831 : tmp34833;
  assign tmp34829 = ~(s2 ? tmp34255 : tmp34830);
  assign tmp34821 = ~(s3 ? tmp34822 : tmp34829);
  assign tmp34803 = s4 ? tmp34804 : tmp34821;
  assign tmp34839 = s0 ? tmp34809 : 0;
  assign tmp34838 = s1 ? tmp34839 : tmp34053;
  assign tmp34842 = l1 ? tmp34079 : tmp33983;
  assign tmp34841 = s0 ? tmp34842 : tmp34271;
  assign tmp34840 = ~(s1 ? tmp34078 : tmp34841);
  assign tmp34837 = s2 ? tmp34838 : tmp34840;
  assign tmp34844 = s1 ? tmp34816 : tmp34780;
  assign tmp34847 = l1 ? tmp34807 : tmp34010;
  assign tmp34849 = l2 ? tmp33948 : tmp33938;
  assign tmp34848 = l1 ? tmp34849 : tmp33987;
  assign tmp34846 = s0 ? tmp34847 : tmp34848;
  assign tmp34845 = ~(s1 ? tmp34013 : tmp34846);
  assign tmp34843 = ~(s2 ? tmp34844 : tmp34845);
  assign tmp34836 = s3 ? tmp34837 : tmp34843;
  assign tmp34853 = s0 ? tmp33977 : tmp34847;
  assign tmp34852 = s1 ? tmp34853 : tmp34287;
  assign tmp34851 = s2 ? tmp34852 : tmp34053;
  assign tmp34857 = l1 ? tmp34046 : tmp34034;
  assign tmp34856 = s0 ? tmp34032 : tmp34857;
  assign tmp34855 = s1 ? tmp34856 : tmp34786;
  assign tmp34854 = ~(s2 ? tmp34855 : tmp34161);
  assign tmp34850 = s3 ? tmp34851 : tmp34854;
  assign tmp34835 = s4 ? tmp34836 : tmp34850;
  assign tmp34862 = ~(l1 ? tmp34056 : 1);
  assign tmp34861 = ~(s1 ? tmp34032 : tmp34862);
  assign tmp34860 = s2 ? tmp34790 : tmp34861;
  assign tmp34859 = s3 ? tmp34860 : tmp34794;
  assign tmp34865 = ~(s1 ? tmp34078 : tmp34082);
  assign tmp34864 = s2 ? tmp34798 : tmp34865;
  assign tmp34863 = s3 ? tmp34864 : tmp34800;
  assign tmp34858 = s4 ? tmp34859 : tmp34863;
  assign tmp34834 = s5 ? tmp34835 : tmp34858;
  assign tmp34802 = s6 ? tmp34803 : tmp34834;
  assign tmp34801 = s7 ? tmp33914 : tmp34802;
  assign tmp34762 = s8 ? tmp34763 : tmp34801;
  assign tmp34872 = l1 ? tmp34807 : tmp34226;
  assign tmp34874 = l1 ? tmp34810 : tmp34226;
  assign tmp34873 = s0 ? tmp34229 : tmp34874;
  assign tmp34871 = s1 ? tmp34872 : tmp34873;
  assign tmp34878 = ~(l1 ? tmp34807 : tmp34227);
  assign tmp34877 = s0 ? tmp34032 : tmp34878;
  assign tmp34880 = l1 ? tmp34046 : tmp33973;
  assign tmp34879 = s0 ? tmp34880 : tmp34878;
  assign tmp34876 = s1 ? tmp34877 : tmp34879;
  assign tmp34882 = s0 ? tmp34880 : 1;
  assign tmp34884 = l1 ? tmp34807 : tmp34227;
  assign tmp34883 = ~(s0 ? tmp34884 : tmp34872);
  assign tmp34881 = s1 ? tmp34882 : tmp34883;
  assign tmp34875 = ~(s2 ? tmp34876 : tmp34881);
  assign tmp34870 = s3 ? tmp34871 : tmp34875;
  assign tmp34889 = l1 ? 1 : tmp33973;
  assign tmp34888 = s0 ? tmp34889 : tmp34247;
  assign tmp34890 = ~(s0 ? tmp34872 : tmp34884);
  assign tmp34887 = s1 ? tmp34888 : tmp34890;
  assign tmp34892 = s0 ? tmp34872 : tmp34251;
  assign tmp34891 = ~(s1 ? tmp34892 : tmp34253);
  assign tmp34886 = s2 ? tmp34887 : tmp34891;
  assign tmp34896 = ~(l1 ? tmp34079 : tmp33942);
  assign tmp34895 = s0 ? tmp34884 : tmp34896;
  assign tmp34897 = s0 ? tmp33985 : tmp34884;
  assign tmp34894 = s1 ? tmp34895 : tmp34897;
  assign tmp34893 = ~(s2 ? tmp34255 : tmp34894);
  assign tmp34885 = ~(s3 ? tmp34886 : tmp34893);
  assign tmp34869 = s4 ? tmp34870 : tmp34885;
  assign tmp34903 = s0 ? tmp34874 : 0;
  assign tmp34902 = s1 ? tmp34903 : tmp34053;
  assign tmp34905 = l1 ? tmp34079 : 1;
  assign tmp34907 = l1 ? tmp34079 : tmp33942;
  assign tmp34906 = s0 ? tmp34907 : tmp34271;
  assign tmp34904 = ~(s1 ? tmp34905 : tmp34906);
  assign tmp34901 = s2 ? tmp34902 : tmp34904;
  assign tmp34910 = ~(l1 ? tmp34009 : tmp34275);
  assign tmp34909 = s1 ? tmp34880 : tmp34910;
  assign tmp34913 = l1 ? tmp34807 : tmp34275;
  assign tmp34914 = l1 ? tmp34849 : tmp33923;
  assign tmp34912 = s0 ? tmp34913 : tmp34914;
  assign tmp34911 = ~(s1 ? tmp34013 : tmp34912);
  assign tmp34908 = ~(s2 ? tmp34909 : tmp34911);
  assign tmp34900 = s3 ? tmp34901 : tmp34908;
  assign tmp34918 = s0 ? tmp33977 : tmp34913;
  assign tmp34917 = s1 ? tmp34918 : tmp34287;
  assign tmp34916 = s2 ? tmp34917 : 0;
  assign tmp34921 = s0 ? 1 : tmp34046;
  assign tmp34922 = ~(l1 ? tmp34009 : tmp34415);
  assign tmp34920 = s1 ? tmp34921 : tmp34922;
  assign tmp34919 = ~(s2 ? tmp34920 : tmp34161);
  assign tmp34915 = s3 ? tmp34916 : tmp34919;
  assign tmp34899 = s4 ? tmp34900 : tmp34915;
  assign tmp34928 = l1 ? tmp34009 : tmp34275;
  assign tmp34927 = s0 ? tmp34928 : tmp34045;
  assign tmp34926 = s1 ? tmp34927 : tmp34791;
  assign tmp34929 = ~(s1 ? 1 : tmp34862);
  assign tmp34925 = s2 ? tmp34926 : tmp34929;
  assign tmp34931 = ~(s1 ? tmp34046 : 1);
  assign tmp34930 = s2 ? tmp34059 : tmp34931;
  assign tmp34924 = s3 ? tmp34925 : tmp34930;
  assign tmp34934 = ~(s1 ? tmp34905 : tmp34082);
  assign tmp34933 = s2 ? tmp34798 : tmp34934;
  assign tmp34936 = ~(l1 ? tmp34079 : tmp34046);
  assign tmp34935 = s1 ? tmp34086 : tmp34936;
  assign tmp34932 = s3 ? tmp34933 : tmp34935;
  assign tmp34923 = s4 ? tmp34924 : tmp34932;
  assign tmp34898 = s5 ? tmp34899 : tmp34923;
  assign tmp34868 = s6 ? tmp34869 : tmp34898;
  assign tmp34867 = s7 ? tmp33914 : tmp34868;
  assign tmp34866 = s8 ? tmp34801 : tmp34867;
  assign tmp34761 = s9 ? tmp34762 : tmp34866;
  assign tmp34938 = s8 ? tmp34801 : tmp33914;
  assign tmp34946 = ~(l1 ? tmp34079 : tmp33939);
  assign tmp34945 = s2 ? tmp34798 : tmp34946;
  assign tmp34944 = s3 ? tmp34945 : tmp34800;
  assign tmp34943 = s4 ? tmp34788 : tmp34944;
  assign tmp34942 = s5 ? tmp34772 : tmp34943;
  assign tmp34941 = s6 ? tmp34765 : tmp34942;
  assign tmp34952 = ~(l1 ? tmp34079 : 1);
  assign tmp34951 = s2 ? tmp34798 : tmp34952;
  assign tmp34950 = s3 ? tmp34951 : tmp34935;
  assign tmp34949 = s4 ? tmp34924 : tmp34950;
  assign tmp34948 = s5 ? tmp34899 : tmp34949;
  assign tmp34947 = s6 ? tmp34869 : tmp34948;
  assign tmp34940 = s7 ? tmp34941 : tmp34947;
  assign tmp34955 = s4 ? tmp34859 : tmp34944;
  assign tmp34954 = s5 ? tmp34835 : tmp34955;
  assign tmp34953 = s6 ? tmp34803 : tmp34954;
  assign tmp34939 = s8 ? tmp34940 : tmp34953;
  assign tmp34937 = s9 ? tmp34938 : tmp34939;
  assign tmp34760 = s10 ? tmp34761 : tmp34937;
  assign tmp34959 = s7 ? tmp34764 : tmp34868;
  assign tmp34958 = s8 ? tmp34959 : tmp34802;
  assign tmp34957 = s9 ? tmp34938 : tmp34958;
  assign tmp34956 = s10 ? tmp34761 : tmp34957;
  assign tmp34759 = s11 ? tmp34760 : tmp34956;
  assign tmp34970 = l1 ? tmp33931 : tmp33941;
  assign tmp34969 = s0 ? tmp33974 : tmp34970;
  assign tmp34968 = s1 ? tmp33954 : tmp34969;
  assign tmp34974 = l1 ? tmp33946 : tmp33939;
  assign tmp34973 = s0 ? tmp34974 : tmp33940;
  assign tmp34972 = s1 ? tmp33935 : tmp34973;
  assign tmp34976 = s0 ? tmp34974 : 1;
  assign tmp34975 = s1 ? tmp34976 : tmp33940;
  assign tmp34971 = ~(s2 ? tmp34972 : tmp34975);
  assign tmp34967 = s3 ? tmp34968 : tmp34971;
  assign tmp34980 = s0 ? tmp33936 : tmp33960;
  assign tmp34979 = s1 ? tmp34980 : tmp33940;
  assign tmp34982 = s0 ? tmp33954 : tmp34251;
  assign tmp34981 = ~(s1 ? tmp34982 : tmp33966);
  assign tmp34978 = s2 ? tmp34979 : tmp34981;
  assign tmp34983 = ~(s2 ? tmp34589 : tmp33979);
  assign tmp34977 = ~(s3 ? tmp34978 : tmp34983);
  assign tmp34966 = s4 ? tmp34967 : tmp34977;
  assign tmp34989 = s0 ? tmp34970 : 0;
  assign tmp34988 = s1 ? tmp34989 : tmp34776;
  assign tmp34991 = s0 ? tmp34000 : tmp34271;
  assign tmp34990 = ~(s1 ? tmp33998 : tmp34991);
  assign tmp34987 = s2 ? tmp34988 : tmp34990;
  assign tmp34993 = s1 ? tmp34974 : tmp34780;
  assign tmp34992 = ~(s2 ? tmp34993 : tmp34781);
  assign tmp34986 = s3 ? tmp34987 : tmp34992;
  assign tmp34985 = s4 ? tmp34986 : tmp34782;
  assign tmp34984 = s5 ? tmp34985 : tmp34858;
  assign tmp34965 = s6 ? tmp34966 : tmp34984;
  assign tmp34964 = s7 ? tmp33914 : tmp34965;
  assign tmp35000 = l1 ? tmp34810 : tmp33941;
  assign tmp34999 = s0 ? tmp34545 : tmp35000;
  assign tmp34998 = s1 ? tmp34820 : tmp34999;
  assign tmp35004 = l1 ? tmp34046 : tmp33939;
  assign tmp35003 = s0 ? tmp35004 : tmp34814;
  assign tmp35002 = s1 ? tmp34813 : tmp35003;
  assign tmp35006 = s0 ? tmp35004 : 1;
  assign tmp35005 = s1 ? tmp35006 : tmp34814;
  assign tmp35001 = ~(s2 ? tmp35002 : tmp35005);
  assign tmp34997 = s3 ? tmp34998 : tmp35001;
  assign tmp35010 = s0 ? tmp34032 : tmp34247;
  assign tmp35009 = s1 ? tmp35010 : tmp34814;
  assign tmp35012 = s0 ? tmp34820 : tmp34251;
  assign tmp35011 = ~(s1 ? tmp35012 : tmp34253);
  assign tmp35008 = s2 ? tmp35009 : tmp35011;
  assign tmp35013 = ~(s2 ? tmp34616 : tmp34830);
  assign tmp35007 = ~(s3 ? tmp35008 : tmp35013);
  assign tmp34996 = s4 ? tmp34997 : tmp35007;
  assign tmp35019 = s0 ? tmp35000 : 0;
  assign tmp35018 = s1 ? tmp35019 : tmp34053;
  assign tmp35017 = s2 ? tmp35018 : tmp34840;
  assign tmp35021 = s1 ? tmp35004 : tmp34780;
  assign tmp35020 = ~(s2 ? tmp35021 : tmp34845);
  assign tmp35016 = s3 ? tmp35017 : tmp35020;
  assign tmp35015 = s4 ? tmp35016 : tmp34850;
  assign tmp35014 = s5 ? tmp35015 : tmp34858;
  assign tmp34995 = s6 ? tmp34996 : tmp35014;
  assign tmp34994 = s7 ? tmp33914 : tmp34995;
  assign tmp34963 = s8 ? tmp34964 : tmp34994;
  assign tmp35029 = l1 ? tmp34810 : tmp34227;
  assign tmp35028 = s0 ? tmp34545 : tmp35029;
  assign tmp35027 = s1 ? tmp34884 : tmp35028;
  assign tmp35032 = s0 ? 1 : tmp34878;
  assign tmp35034 = l1 ? tmp34046 : 1;
  assign tmp35033 = s0 ? tmp35034 : tmp34878;
  assign tmp35031 = s1 ? tmp35032 : tmp35033;
  assign tmp35036 = s0 ? tmp35034 : 1;
  assign tmp35035 = s1 ? tmp35036 : tmp34878;
  assign tmp35030 = ~(s2 ? tmp35031 : tmp35035);
  assign tmp35026 = s3 ? tmp35027 : tmp35030;
  assign tmp35040 = s0 ? 1 : tmp34247;
  assign tmp35039 = s1 ? tmp35040 : tmp34878;
  assign tmp35042 = s0 ? tmp34884 : tmp34251;
  assign tmp35041 = ~(s1 ? tmp35042 : tmp34253);
  assign tmp35038 = s2 ? tmp35039 : tmp35041;
  assign tmp35043 = ~(s2 ? tmp34616 : tmp34894);
  assign tmp35037 = ~(s3 ? tmp35038 : tmp35043);
  assign tmp35025 = s4 ? tmp35026 : tmp35037;
  assign tmp35049 = s0 ? tmp35029 : 0;
  assign tmp35048 = s1 ? tmp35049 : 0;
  assign tmp35047 = s2 ? tmp35048 : tmp34904;
  assign tmp35051 = s1 ? tmp35034 : tmp34910;
  assign tmp35050 = ~(s2 ? tmp35051 : tmp34911);
  assign tmp35046 = s3 ? tmp35047 : tmp35050;
  assign tmp35045 = s4 ? tmp35046 : tmp34915;
  assign tmp35044 = s5 ? tmp35045 : tmp34923;
  assign tmp35024 = s6 ? tmp35025 : tmp35044;
  assign tmp35023 = s7 ? tmp33914 : tmp35024;
  assign tmp35022 = s8 ? tmp34994 : tmp35023;
  assign tmp34962 = s9 ? tmp34963 : tmp35022;
  assign tmp35053 = s8 ? tmp34994 : tmp33914;
  assign tmp35057 = s5 ? tmp34985 : tmp34955;
  assign tmp35056 = s6 ? tmp34966 : tmp35057;
  assign tmp35059 = s5 ? tmp35045 : tmp34949;
  assign tmp35058 = s6 ? tmp35025 : tmp35059;
  assign tmp35055 = s7 ? tmp35056 : tmp35058;
  assign tmp35061 = s5 ? tmp35015 : tmp34955;
  assign tmp35060 = s6 ? tmp34996 : tmp35061;
  assign tmp35054 = s8 ? tmp35055 : tmp35060;
  assign tmp35052 = s9 ? tmp35053 : tmp35054;
  assign tmp34961 = s10 ? tmp34962 : tmp35052;
  assign tmp35065 = s7 ? tmp34965 : tmp35024;
  assign tmp35064 = s8 ? tmp35065 : tmp34995;
  assign tmp35063 = s9 ? tmp35053 : tmp35064;
  assign tmp35062 = s10 ? tmp34962 : tmp35063;
  assign tmp34960 = s11 ? tmp34961 : tmp35062;
  assign tmp34758 = s12 ? tmp34759 : tmp34960;
  assign tmp34648 = s13 ? tmp34649 : tmp34758;
  assign tmp33907 = s14 ? tmp33908 : tmp34648;
  assign tmp35079 = ~(l1 ? 1 : tmp34024);
  assign tmp35078 = ~(s0 ? tmp34048 : tmp35079);
  assign tmp35077 = s1 ? tmp34297 : tmp35078;
  assign tmp35076 = s2 ? tmp35077 : tmp34419;
  assign tmp35075 = s3 ? tmp35076 : tmp34300;
  assign tmp35082 = ~(s0 ? tmp34048 : tmp34268);
  assign tmp35081 = s2 ? tmp34175 : tmp35082;
  assign tmp35080 = s3 ? tmp35081 : tmp34305;
  assign tmp35074 = s4 ? tmp35075 : tmp35080;
  assign tmp35073 = s5 ? tmp34562 : tmp35074;
  assign tmp35072 = s6 ? tmp34628 : tmp35073;
  assign tmp35071 = s7 ? tmp33914 : tmp35072;
  assign tmp35084 = s8 ? tmp35071 : tmp33914;
  assign tmp35087 = s4 ? tmp35075 : tmp34302;
  assign tmp35086 = s5 ? tmp34562 : tmp35087;
  assign tmp35085 = s6 ? tmp34628 : tmp35086;
  assign tmp35083 = s9 ? tmp35084 : tmp35085;
  assign tmp35070 = s10 ? tmp35071 : tmp35083;
  assign tmp35089 = s9 ? tmp35084 : tmp35072;
  assign tmp35088 = s10 ? tmp35071 : tmp35089;
  assign tmp35069 = s11 ? tmp35070 : tmp35088;
  assign tmp35097 = ~(s2 ? tmp34413 : tmp34038);
  assign tmp35096 = s3 ? tmp34283 : tmp35097;
  assign tmp35095 = s4 ? tmp34563 : tmp35096;
  assign tmp35094 = s5 ? tmp35095 : tmp34416;
  assign tmp35093 = s6 ? tmp34628 : tmp35094;
  assign tmp35092 = s7 ? tmp33914 : tmp35093;
  assign tmp35099 = s8 ? tmp35092 : tmp33914;
  assign tmp35098 = s9 ? tmp35099 : tmp34627;
  assign tmp35091 = s10 ? tmp35092 : tmp35098;
  assign tmp35101 = s9 ? tmp35099 : tmp35093;
  assign tmp35100 = s10 ? tmp35092 : tmp35101;
  assign tmp35090 = s11 ? tmp35091 : tmp35100;
  assign tmp35068 = s12 ? tmp35069 : tmp35090;
  assign tmp35113 = s0 ? tmp34067 : tmp34234;
  assign tmp35112 = ~(s1 ? tmp34046 : tmp35113);
  assign tmp35111 = s2 ? tmp34171 : tmp35112;
  assign tmp35110 = s3 ? tmp34418 : tmp35111;
  assign tmp35116 = ~(l1 ? tmp34046 : tmp34068);
  assign tmp35115 = s2 ? tmp34305 : tmp35116;
  assign tmp35114 = s3 ? tmp34303 : tmp35115;
  assign tmp35109 = s4 ? tmp35110 : tmp35114;
  assign tmp35108 = s5 ? tmp34562 : tmp35109;
  assign tmp35107 = s6 ? tmp34628 : tmp35108;
  assign tmp35106 = s7 ? tmp33914 : tmp35107;
  assign tmp35124 = s0 ? tmp34234 : tmp34318;
  assign tmp35125 = s0 ? tmp34550 : tmp34318;
  assign tmp35123 = s1 ? tmp35124 : tmp35125;
  assign tmp35126 = s1 ? tmp34632 : tmp34318;
  assign tmp35122 = ~(s2 ? tmp35123 : tmp35126);
  assign tmp35121 = s3 ? tmp34733 : tmp35122;
  assign tmp35120 = s4 ? tmp35121 : tmp34735;
  assign tmp35131 = s1 ? tmp34714 : tmp34266;
  assign tmp35130 = s2 ? tmp35131 : tmp34340;
  assign tmp35133 = s1 ? tmp34550 : tmp34143;
  assign tmp35132 = ~(s2 ? tmp35133 : tmp34277);
  assign tmp35129 = s3 ? tmp35130 : tmp35132;
  assign tmp35128 = s4 ? tmp35129 : tmp34344;
  assign tmp35136 = s2 ? tmp34165 : tmp34419;
  assign tmp35139 = s0 ? tmp34067 : tmp34103;
  assign tmp35138 = ~(s1 ? tmp34046 : tmp35139);
  assign tmp35137 = s2 ? tmp34171 : tmp35138;
  assign tmp35135 = s3 ? tmp35136 : tmp35137;
  assign tmp35141 = s2 ? tmp34177 : tmp35116;
  assign tmp35140 = s3 ? tmp34174 : tmp35141;
  assign tmp35134 = s4 ? tmp35135 : tmp35140;
  assign tmp35127 = s5 ? tmp35128 : tmp35134;
  assign tmp35119 = s6 ? tmp35120 : tmp35127;
  assign tmp35118 = s7 ? tmp33914 : tmp35119;
  assign tmp35117 = s8 ? tmp35106 : tmp35118;
  assign tmp35105 = s9 ? tmp35106 : tmp35117;
  assign tmp35143 = s8 ? tmp35106 : tmp33914;
  assign tmp35148 = s4 ? tmp35110 : tmp34302;
  assign tmp35147 = s5 ? tmp34562 : tmp35148;
  assign tmp35146 = s6 ? tmp34628 : tmp35147;
  assign tmp35151 = s4 ? tmp35135 : tmp34173;
  assign tmp35150 = s5 ? tmp35128 : tmp35151;
  assign tmp35149 = s6 ? tmp35120 : tmp35150;
  assign tmp35145 = s7 ? tmp35146 : tmp35149;
  assign tmp35144 = s8 ? tmp35145 : tmp35146;
  assign tmp35142 = s9 ? tmp35143 : tmp35144;
  assign tmp35104 = s10 ? tmp35105 : tmp35142;
  assign tmp35155 = s7 ? tmp35107 : tmp35119;
  assign tmp35154 = s8 ? tmp35155 : tmp35107;
  assign tmp35153 = s9 ? tmp35143 : tmp35154;
  assign tmp35152 = s10 ? tmp35105 : tmp35153;
  assign tmp35103 = s11 ? tmp35104 : tmp35152;
  assign tmp35163 = s1 ? tmp34064 : tmp34266;
  assign tmp35162 = s2 ? tmp34171 : tmp35163;
  assign tmp35161 = s3 ? tmp34418 : tmp35162;
  assign tmp35166 = s0 ? 1 : tmp34306;
  assign tmp35165 = s1 ? tmp34061 : tmp35166;
  assign tmp35164 = s3 ? tmp34303 : tmp35165;
  assign tmp35160 = s4 ? tmp35161 : tmp35164;
  assign tmp35159 = s5 ? tmp34562 : tmp35160;
  assign tmp35158 = s6 ? tmp34628 : tmp35159;
  assign tmp35157 = s7 ? tmp33914 : tmp35158;
  assign tmp35168 = s8 ? tmp35157 : tmp33914;
  assign tmp35167 = s9 ? tmp35168 : tmp35158;
  assign tmp35156 = s10 ? tmp35157 : tmp35167;
  assign tmp35102 = s12 ? tmp35103 : tmp35156;
  assign tmp35067 = s13 ? tmp35068 : tmp35102;
  assign tmp35181 = s1 ? tmp34036 : tmp34776;
  assign tmp35180 = s2 ? tmp34020 : tmp35181;
  assign tmp35182 = ~(s2 ? tmp34030 : tmp34161);
  assign tmp35179 = s3 ? tmp35180 : tmp35182;
  assign tmp35178 = s4 ? tmp34986 : tmp35179;
  assign tmp35187 = ~(l1 ? tmp33986 : tmp33987);
  assign tmp35186 = s1 ? tmp34072 : tmp35187;
  assign tmp35188 = s1 ? tmp34078 : tmp34082;
  assign tmp35185 = s2 ? tmp35186 : tmp35188;
  assign tmp35190 = ~(l1 ? tmp34050 : tmp33932);
  assign tmp35189 = ~(s2 ? tmp34800 : tmp35190);
  assign tmp35184 = ~(s3 ? tmp35185 : tmp35189);
  assign tmp35183 = s4 ? tmp34859 : tmp35184;
  assign tmp35177 = s5 ? tmp35178 : tmp35183;
  assign tmp35176 = s6 ? tmp34966 : tmp35177;
  assign tmp35175 = s7 ? tmp33914 : tmp35176;
  assign tmp35193 = s5 ? tmp35015 : tmp35183;
  assign tmp35192 = s6 ? tmp34996 : tmp35193;
  assign tmp35191 = s7 ? tmp33914 : tmp35192;
  assign tmp35174 = s8 ? tmp35175 : tmp35191;
  assign tmp35201 = s0 ? 1 : tmp34814;
  assign tmp35202 = s0 ? tmp35034 : tmp34814;
  assign tmp35200 = s1 ? tmp35201 : tmp35202;
  assign tmp35203 = s1 ? tmp35036 : tmp34814;
  assign tmp35199 = ~(s2 ? tmp35200 : tmp35203);
  assign tmp35198 = s3 ? tmp34998 : tmp35199;
  assign tmp35197 = s4 ? tmp35198 : tmp35007;
  assign tmp35208 = s1 ? tmp35019 : 0;
  assign tmp35207 = s2 ? tmp35208 : tmp34840;
  assign tmp35210 = s1 ? tmp35034 : tmp34780;
  assign tmp35209 = ~(s2 ? tmp35210 : tmp34845);
  assign tmp35206 = s3 ? tmp35207 : tmp35209;
  assign tmp35205 = s4 ? tmp35206 : tmp34850;
  assign tmp35213 = s2 ? tmp34790 : tmp34929;
  assign tmp35212 = s3 ? tmp35213 : tmp34794;
  assign tmp35211 = s4 ? tmp35212 : tmp35184;
  assign tmp35204 = s5 ? tmp35205 : tmp35211;
  assign tmp35196 = s6 ? tmp35197 : tmp35204;
  assign tmp35195 = s7 ? tmp33914 : tmp35196;
  assign tmp35194 = s8 ? tmp35191 : tmp35195;
  assign tmp35173 = s9 ? tmp35174 : tmp35194;
  assign tmp35215 = s8 ? tmp35191 : tmp33914;
  assign tmp35221 = s3 ? tmp35180 : tmp34784;
  assign tmp35220 = s4 ? tmp34986 : tmp35221;
  assign tmp35224 = s2 ? tmp35186 : tmp34078;
  assign tmp35225 = ~(s1 ? tmp34086 : tmp34088);
  assign tmp35223 = ~(s3 ? tmp35224 : tmp35225);
  assign tmp35222 = s4 ? tmp34859 : tmp35223;
  assign tmp35219 = s5 ? tmp35220 : tmp35222;
  assign tmp35218 = s6 ? tmp34966 : tmp35219;
  assign tmp35228 = s4 ? tmp35212 : tmp35223;
  assign tmp35227 = s5 ? tmp35205 : tmp35228;
  assign tmp35226 = s6 ? tmp35197 : tmp35227;
  assign tmp35217 = s7 ? tmp35218 : tmp35226;
  assign tmp35230 = s5 ? tmp35015 : tmp35222;
  assign tmp35229 = s6 ? tmp34996 : tmp35230;
  assign tmp35216 = s8 ? tmp35217 : tmp35229;
  assign tmp35214 = s9 ? tmp35215 : tmp35216;
  assign tmp35172 = s10 ? tmp35173 : tmp35214;
  assign tmp35234 = s7 ? tmp35176 : tmp35196;
  assign tmp35233 = s8 ? tmp35234 : tmp35192;
  assign tmp35232 = s9 ? tmp35215 : tmp35233;
  assign tmp35231 = s10 ? tmp35173 : tmp35232;
  assign tmp35171 = s11 ? tmp35172 : tmp35231;
  assign tmp35243 = s0 ? tmp34545 : tmp34970;
  assign tmp35242 = s1 ? tmp33954 : tmp35243;
  assign tmp35241 = s3 ? tmp35242 : tmp34971;
  assign tmp35247 = s0 ? tmp33936 : tmp34247;
  assign tmp35246 = s1 ? tmp35247 : tmp33940;
  assign tmp35248 = ~(s1 ? tmp34982 : tmp34253);
  assign tmp35245 = s2 ? tmp35246 : tmp35248;
  assign tmp35249 = ~(s2 ? tmp34616 : tmp33979);
  assign tmp35244 = ~(s3 ? tmp35245 : tmp35249);
  assign tmp35240 = s4 ? tmp35241 : tmp35244;
  assign tmp35254 = s1 ? tmp34021 : tmp34287;
  assign tmp35253 = s2 ? tmp35254 : tmp34776;
  assign tmp35252 = s3 ? tmp35253 : tmp34784;
  assign tmp35251 = s4 ? tmp34986 : tmp35252;
  assign tmp35258 = s1 ? tmp34052 : tmp34055;
  assign tmp35257 = s2 ? tmp34790 : tmp35258;
  assign tmp35259 = s2 ? tmp34171 : tmp34795;
  assign tmp35256 = s3 ? tmp35257 : tmp35259;
  assign tmp35261 = s1 ? tmp34085 : tmp34088;
  assign tmp35260 = s3 ? tmp34945 : tmp35261;
  assign tmp35255 = s4 ? tmp35256 : tmp35260;
  assign tmp35250 = s5 ? tmp35251 : tmp35255;
  assign tmp35239 = s6 ? tmp35240 : tmp35250;
  assign tmp35238 = s7 ? tmp33914 : tmp35239;
  assign tmp35266 = s3 ? tmp34860 : tmp35259;
  assign tmp35265 = s4 ? tmp35266 : tmp34944;
  assign tmp35264 = s5 ? tmp35015 : tmp35265;
  assign tmp35263 = s6 ? tmp34996 : tmp35264;
  assign tmp35262 = s7 ? tmp33914 : tmp35263;
  assign tmp35237 = s8 ? tmp35238 : tmp35262;
  assign tmp35275 = ~(l1 ? tmp34056 : tmp33939);
  assign tmp35274 = ~(s1 ? 1 : tmp35275);
  assign tmp35273 = s2 ? tmp34926 : tmp35274;
  assign tmp35276 = s2 ? tmp34171 : tmp34931;
  assign tmp35272 = s3 ? tmp35273 : tmp35276;
  assign tmp35271 = s4 ? tmp35272 : tmp34950;
  assign tmp35270 = s5 ? tmp35045 : tmp35271;
  assign tmp35269 = s6 ? tmp35025 : tmp35270;
  assign tmp35268 = s7 ? tmp33914 : tmp35269;
  assign tmp35267 = s8 ? tmp35262 : tmp35268;
  assign tmp35236 = s9 ? tmp35237 : tmp35267;
  assign tmp35278 = s8 ? tmp35262 : tmp33914;
  assign tmp35280 = s7 ? tmp35239 : tmp35269;
  assign tmp35279 = s8 ? tmp35280 : tmp35263;
  assign tmp35277 = s9 ? tmp35278 : tmp35279;
  assign tmp35235 = s10 ? tmp35236 : tmp35277;
  assign tmp35170 = s12 ? tmp35171 : tmp35235;
  assign tmp35289 = s2 ? tmp34305 : 1;
  assign tmp35288 = s3 ? tmp34303 : tmp35289;
  assign tmp35287 = s4 ? tmp34417 : tmp35288;
  assign tmp35286 = s5 ? tmp34562 : tmp35287;
  assign tmp35285 = s6 ? tmp34628 : tmp35286;
  assign tmp35284 = s7 ? tmp33914 : tmp35285;
  assign tmp35295 = s3 ? tmp35136 : tmp34170;
  assign tmp35297 = s2 ? tmp34177 : 1;
  assign tmp35296 = s3 ? tmp34174 : tmp35297;
  assign tmp35294 = s4 ? tmp35295 : tmp35296;
  assign tmp35293 = s5 ? tmp35128 : tmp35294;
  assign tmp35292 = s6 ? tmp35120 : tmp35293;
  assign tmp35291 = s7 ? tmp33914 : tmp35292;
  assign tmp35290 = s8 ? tmp35284 : tmp35291;
  assign tmp35283 = s9 ? tmp35284 : tmp35290;
  assign tmp35299 = s8 ? tmp35284 : tmp33914;
  assign tmp35301 = s7 ? tmp35285 : tmp35292;
  assign tmp35300 = s8 ? tmp35301 : tmp35285;
  assign tmp35298 = s9 ? tmp35299 : tmp35300;
  assign tmp35282 = s10 ? tmp35283 : tmp35298;
  assign tmp35307 = s4 ? tmp34967 : tmp35244;
  assign tmp35313 = s0 ? 1 : tmp33985;
  assign tmp35312 = s1 ? tmp34086 : tmp35313;
  assign tmp35311 = s2 ? tmp35312 : tmp34946;
  assign tmp35314 = s2 ? tmp34800 : 1;
  assign tmp35310 = s3 ? tmp35311 : tmp35314;
  assign tmp35309 = s4 ? tmp35266 : tmp35310;
  assign tmp35308 = s5 ? tmp35251 : tmp35309;
  assign tmp35306 = s6 ? tmp35307 : tmp35308;
  assign tmp35305 = s7 ? tmp33914 : tmp35306;
  assign tmp35317 = s5 ? tmp35015 : tmp35309;
  assign tmp35316 = s6 ? tmp34996 : tmp35317;
  assign tmp35315 = s7 ? tmp33914 : tmp35316;
  assign tmp35304 = s8 ? tmp35305 : tmp35315;
  assign tmp35324 = s2 ? tmp34790 : tmp35274;
  assign tmp35323 = s3 ? tmp35324 : tmp35259;
  assign tmp35322 = s4 ? tmp35323 : tmp35310;
  assign tmp35321 = s5 ? tmp35205 : tmp35322;
  assign tmp35320 = s6 ? tmp35197 : tmp35321;
  assign tmp35319 = s7 ? tmp33914 : tmp35320;
  assign tmp35318 = s8 ? tmp35315 : tmp35319;
  assign tmp35303 = s9 ? tmp35304 : tmp35318;
  assign tmp35326 = s8 ? tmp35315 : tmp33914;
  assign tmp35328 = s7 ? tmp35306 : tmp35320;
  assign tmp35327 = s8 ? tmp35328 : tmp35316;
  assign tmp35325 = s9 ? tmp35326 : tmp35327;
  assign tmp35302 = s10 ? tmp35303 : tmp35325;
  assign tmp35281 = s12 ? tmp35282 : tmp35302;
  assign tmp35169 = s13 ? tmp35170 : tmp35281;
  assign tmp35066 = s14 ? tmp35067 : tmp35169;
  assign tmp33906 = s15 ? tmp33907 : tmp35066;
  assign tmp35343 = s0 ? tmp34189 : tmp33952;
  assign tmp35342 = ~(s1 ? tmp33952 : tmp35343);
  assign tmp35341 = s2 ? tmp34152 : tmp35342;
  assign tmp35340 = s3 ? tmp35341 : tmp34215;
  assign tmp35339 = s4 ? tmp34204 : tmp35340;
  assign tmp35338 = s5 ? tmp35339 : tmp34162;
  assign tmp35337 = s6 ? tmp34181 : tmp35338;
  assign tmp35336 = s7 ? tmp33914 : tmp35337;
  assign tmp35335 = s8 ? tmp33913 : tmp35336;
  assign tmp35334 = s9 ? tmp35335 : tmp35336;
  assign tmp35345 = s8 ? tmp35336 : tmp33914;
  assign tmp35353 = s1 ? tmp34451 : tmp34463;
  assign tmp35352 = s2 ? tmp35353 : tmp34524;
  assign tmp35351 = s3 ? tmp35352 : tmp34456;
  assign tmp35356 = ~(s1 ? tmp33952 : tmp34431);
  assign tmp35355 = s2 ? tmp34461 : tmp35356;
  assign tmp35358 = s1 ? tmp34466 : tmp34160;
  assign tmp35357 = ~(s2 ? tmp35358 : tmp34161);
  assign tmp35354 = s3 ? tmp35355 : tmp35357;
  assign tmp35350 = s4 ? tmp35351 : tmp35354;
  assign tmp35349 = s5 ? tmp35350 : tmp34293;
  assign tmp35348 = s6 ? tmp34422 : tmp35349;
  assign tmp35347 = s7 ? tmp34350 : tmp35348;
  assign tmp35364 = ~(s1 ? tmp33952 : tmp34189);
  assign tmp35363 = s2 ? tmp34152 : tmp35364;
  assign tmp35362 = s3 ? tmp35363 : tmp34215;
  assign tmp35361 = s4 ? tmp34204 : tmp35362;
  assign tmp35360 = s5 ? tmp35361 : tmp34162;
  assign tmp35359 = s6 ? tmp34181 : tmp35360;
  assign tmp35346 = s8 ? tmp35347 : tmp35359;
  assign tmp35344 = s9 ? tmp35345 : tmp35346;
  assign tmp35333 = s10 ? tmp35334 : tmp35344;
  assign tmp35375 = s0 ? tmp34431 : tmp33952;
  assign tmp35374 = ~(s1 ? tmp33952 : tmp35375);
  assign tmp35373 = s2 ? tmp34461 : tmp35374;
  assign tmp35372 = s3 ? tmp35373 : tmp35357;
  assign tmp35371 = s4 ? tmp35351 : tmp35372;
  assign tmp35370 = s5 ? tmp35371 : tmp34293;
  assign tmp35369 = s6 ? tmp34422 : tmp35370;
  assign tmp35368 = s7 ? tmp34091 : tmp35369;
  assign tmp35367 = s8 ? tmp35368 : tmp35337;
  assign tmp35366 = s9 ? tmp35345 : tmp35367;
  assign tmp35365 = s10 ? tmp35334 : tmp35366;
  assign tmp35332 = s11 ? tmp35333 : tmp35365;
  assign tmp35386 = ~(s1 ? tmp34587 : tmp33965);
  assign tmp35385 = s2 ? tmp34584 : tmp35386;
  assign tmp35388 = s1 ? tmp33974 : tmp33976;
  assign tmp35387 = ~(s2 ? tmp35388 : tmp34388);
  assign tmp35384 = ~(s3 ? tmp35385 : tmp35387);
  assign tmp35383 = s4 ? tmp34572 : tmp35384;
  assign tmp35382 = s6 ? tmp35383 : tmp34590;
  assign tmp35381 = s7 ? tmp33914 : tmp35382;
  assign tmp35380 = s8 ? tmp34539 : tmp35381;
  assign tmp35394 = s1 ? tmp34112 : tmp34574;
  assign tmp35398 = l1 ? tmp34192 : tmp33939;
  assign tmp35397 = s0 ? tmp35398 : tmp34104;
  assign tmp35396 = s1 ? tmp34188 : tmp35397;
  assign tmp35400 = s0 ? tmp35398 : tmp33952;
  assign tmp35399 = s1 ? tmp35400 : tmp34104;
  assign tmp35395 = ~(s2 ? tmp35396 : tmp35399);
  assign tmp35393 = s3 ? tmp35394 : tmp35395;
  assign tmp35403 = s1 ? tmp34585 : tmp34104;
  assign tmp35405 = s0 ? tmp34112 : tmp33964;
  assign tmp35404 = ~(s1 ? tmp35405 : tmp33965);
  assign tmp35402 = s2 ? tmp35403 : tmp35404;
  assign tmp35406 = ~(s2 ? tmp35388 : tmp34124);
  assign tmp35401 = ~(s3 ? tmp35402 : tmp35406);
  assign tmp35392 = s4 ? tmp35393 : tmp35401;
  assign tmp35411 = s1 ? tmp34595 : tmp34208;
  assign tmp35412 = ~(s1 ? tmp34455 : tmp34139);
  assign tmp35410 = s2 ? tmp35411 : tmp35412;
  assign tmp35414 = s1 ? tmp35398 : tmp34274;
  assign tmp35413 = ~(s2 ? tmp35414 : tmp34458);
  assign tmp35409 = s3 ? tmp35410 : tmp35413;
  assign tmp35408 = s4 ? tmp35409 : tmp34459;
  assign tmp35407 = s5 ? tmp35408 : tmp34416;
  assign tmp35391 = s6 ? tmp35392 : tmp35407;
  assign tmp35390 = s7 ? tmp33914 : tmp35391;
  assign tmp35389 = s8 ? tmp35381 : tmp35390;
  assign tmp35379 = s9 ? tmp35380 : tmp35389;
  assign tmp35416 = s8 ? tmp35381 : tmp33914;
  assign tmp35422 = ~(s2 ? tmp34589 : tmp34124);
  assign tmp35421 = ~(s3 ? tmp35402 : tmp35422);
  assign tmp35420 = s4 ? tmp35393 : tmp35421;
  assign tmp35419 = s6 ? tmp35420 : tmp35407;
  assign tmp35418 = s7 ? tmp34640 : tmp35419;
  assign tmp35425 = ~(s3 ? tmp35385 : tmp34588);
  assign tmp35424 = s4 ? tmp34572 : tmp35425;
  assign tmp35423 = s6 ? tmp35424 : tmp34590;
  assign tmp35417 = s8 ? tmp35418 : tmp35423;
  assign tmp35415 = s9 ? tmp35416 : tmp35417;
  assign tmp35378 = s10 ? tmp35379 : tmp35415;
  assign tmp35429 = s7 ? tmp34540 : tmp35391;
  assign tmp35428 = s8 ? tmp35429 : tmp35382;
  assign tmp35427 = s9 ? tmp35416 : tmp35428;
  assign tmp35426 = s10 ? tmp35379 : tmp35427;
  assign tmp35377 = s11 ? tmp35378 : tmp35426;
  assign tmp35376 = s12 ? tmp34362 : tmp35377;
  assign tmp35331 = s13 ? tmp35332 : tmp35376;
  assign tmp35442 = ~(l1 ? tmp34192 : tmp33973);
  assign tmp35441 = s0 ? 1 : tmp35442;
  assign tmp35440 = s1 ? tmp35441 : tmp34406;
  assign tmp35439 = s2 ? tmp35440 : tmp34407;
  assign tmp35438 = s3 ? tmp35352 : tmp35439;
  assign tmp35437 = s4 ? tmp35438 : tmp34459;
  assign tmp35436 = s5 ? tmp35437 : tmp34416;
  assign tmp35435 = s6 ? tmp34422 : tmp35436;
  assign tmp35434 = s7 ? tmp33914 : tmp35435;
  assign tmp35452 = ~(l1 ? tmp34192 : tmp33947);
  assign tmp35451 = s0 ? 1 : tmp35452;
  assign tmp35453 = s0 ? 1 : tmp34167;
  assign tmp35450 = s1 ? tmp35451 : tmp35453;
  assign tmp35454 = s1 ? tmp34146 : tmp34147;
  assign tmp35449 = s2 ? tmp35450 : tmp35454;
  assign tmp35448 = s3 ? tmp34205 : tmp35449;
  assign tmp35456 = s2 ? tmp34461 : tmp34208;
  assign tmp35459 = s0 ? tmp34103 : tmp34467;
  assign tmp35458 = s1 ? tmp35459 : tmp34414;
  assign tmp35457 = ~(s2 ? tmp35458 : tmp34161);
  assign tmp35455 = s3 ? tmp35456 : tmp35457;
  assign tmp35447 = s4 ? tmp35448 : tmp35455;
  assign tmp35446 = s5 ? tmp35447 : tmp34681;
  assign tmp35445 = s6 ? tmp34181 : tmp35446;
  assign tmp35444 = s7 ? tmp33914 : tmp35445;
  assign tmp35443 = s8 ? tmp35434 : tmp35444;
  assign tmp35433 = s9 ? tmp35434 : tmp35443;
  assign tmp35461 = s8 ? tmp35434 : tmp33914;
  assign tmp35463 = s7 ? tmp34654 : tmp35445;
  assign tmp35462 = s8 ? tmp35463 : tmp35435;
  assign tmp35460 = s9 ? tmp35461 : tmp35462;
  assign tmp35432 = s10 ? tmp35433 : tmp35460;
  assign tmp35472 = l1 ? tmp33927 : tmp33941;
  assign tmp35471 = s0 ? tmp33974 : tmp35472;
  assign tmp35470 = s1 ? tmp34112 : tmp35471;
  assign tmp35469 = s3 ? tmp35470 : tmp35395;
  assign tmp35476 = s0 ? tmp34189 : tmp33960;
  assign tmp35475 = s1 ? tmp35476 : tmp34104;
  assign tmp35477 = ~(s1 ? tmp35405 : tmp33966);
  assign tmp35474 = s2 ? tmp35475 : tmp35477;
  assign tmp35473 = ~(s3 ? tmp35474 : tmp35422);
  assign tmp35468 = s4 ? tmp35469 : tmp35473;
  assign tmp35483 = s0 ? tmp35472 : 0;
  assign tmp35482 = s1 ? tmp35483 : tmp34208;
  assign tmp35481 = s2 ? tmp35482 : tmp34209;
  assign tmp35485 = s1 ? tmp35398 : tmp34143;
  assign tmp35484 = ~(s2 ? tmp35485 : tmp34145);
  assign tmp35480 = s3 ? tmp35481 : tmp35484;
  assign tmp35488 = s1 ? tmp34036 : tmp34208;
  assign tmp35487 = s2 ? tmp34152 : tmp35488;
  assign tmp35490 = s1 ? tmp34217 : tmp34727;
  assign tmp35489 = ~(s2 ? tmp35490 : tmp34161);
  assign tmp35486 = s3 ? tmp35487 : tmp35489;
  assign tmp35479 = s4 ? tmp35480 : tmp35486;
  assign tmp35478 = s5 ? tmp35479 : tmp34162;
  assign tmp35467 = s6 ? tmp35468 : tmp35478;
  assign tmp35466 = s7 ? tmp33914 : tmp35467;
  assign tmp35492 = s8 ? tmp35466 : tmp33914;
  assign tmp35496 = s3 ? tmp35487 : tmp34215;
  assign tmp35495 = s4 ? tmp35480 : tmp35496;
  assign tmp35494 = s5 ? tmp35495 : tmp34162;
  assign tmp35493 = s6 ? tmp35468 : tmp35494;
  assign tmp35491 = s9 ? tmp35492 : tmp35493;
  assign tmp35465 = s10 ? tmp35466 : tmp35491;
  assign tmp35498 = s9 ? tmp35492 : tmp35467;
  assign tmp35497 = s10 ? tmp35466 : tmp35498;
  assign tmp35464 = s11 ? tmp35465 : tmp35497;
  assign tmp35431 = s12 ? tmp35432 : tmp35464;
  assign tmp35506 = s5 ? tmp34772 : tmp35265;
  assign tmp35505 = s6 ? tmp34765 : tmp35506;
  assign tmp35504 = s7 ? tmp33914 : tmp35505;
  assign tmp35509 = s5 ? tmp34835 : tmp35265;
  assign tmp35508 = s6 ? tmp34803 : tmp35509;
  assign tmp35507 = s7 ? tmp33914 : tmp35508;
  assign tmp35503 = s8 ? tmp35504 : tmp35507;
  assign tmp35513 = s5 ? tmp34835 : tmp34787;
  assign tmp35512 = s6 ? tmp34803 : tmp35513;
  assign tmp35511 = s7 ? tmp33914 : tmp35512;
  assign tmp35510 = s8 ? tmp35507 : tmp35511;
  assign tmp35502 = s9 ? tmp35503 : tmp35510;
  assign tmp35515 = s8 ? tmp35507 : tmp33914;
  assign tmp35522 = s1 ? tmp35032 : tmp34879;
  assign tmp35521 = ~(s2 ? tmp35522 : tmp34881);
  assign tmp35520 = s3 ? tmp34871 : tmp35521;
  assign tmp35519 = s4 ? tmp35520 : tmp34885;
  assign tmp35527 = s1 ? tmp34903 : 0;
  assign tmp35528 = ~(s1 ? tmp34078 : tmp34906);
  assign tmp35526 = s2 ? tmp35527 : tmp35528;
  assign tmp35530 = s1 ? tmp34880 : tmp34780;
  assign tmp35529 = ~(s2 ? tmp35530 : tmp34845);
  assign tmp35525 = s3 ? tmp35526 : tmp35529;
  assign tmp35532 = s2 ? tmp34917 : tmp34053;
  assign tmp35535 = s0 ? tmp34032 : tmp34046;
  assign tmp35534 = s1 ? tmp35535 : tmp34922;
  assign tmp35533 = ~(s2 ? tmp35534 : tmp34161);
  assign tmp35531 = s3 ? tmp35532 : tmp35533;
  assign tmp35524 = s4 ? tmp35525 : tmp35531;
  assign tmp35537 = s3 ? tmp34789 : tmp34930;
  assign tmp35538 = s3 ? tmp34945 : tmp34935;
  assign tmp35536 = s4 ? tmp35537 : tmp35538;
  assign tmp35523 = s5 ? tmp35524 : tmp35536;
  assign tmp35518 = s6 ? tmp35519 : tmp35523;
  assign tmp35517 = s7 ? tmp35505 : tmp35518;
  assign tmp35516 = s8 ? tmp35517 : tmp35508;
  assign tmp35514 = s9 ? tmp35515 : tmp35516;
  assign tmp35501 = s10 ? tmp35502 : tmp35514;
  assign tmp35546 = s3 ? tmp34797 : tmp34935;
  assign tmp35545 = s4 ? tmp35537 : tmp35546;
  assign tmp35544 = s5 ? tmp35524 : tmp35545;
  assign tmp35543 = s6 ? tmp35519 : tmp35544;
  assign tmp35542 = s7 ? tmp35505 : tmp35543;
  assign tmp35541 = s8 ? tmp35542 : tmp35508;
  assign tmp35540 = s9 ? tmp35515 : tmp35541;
  assign tmp35539 = s10 ? tmp35502 : tmp35540;
  assign tmp35500 = s11 ? tmp35501 : tmp35539;
  assign tmp35553 = s5 ? tmp34985 : tmp35265;
  assign tmp35552 = s6 ? tmp34966 : tmp35553;
  assign tmp35551 = s7 ? tmp33914 : tmp35552;
  assign tmp35550 = s8 ? tmp35551 : tmp35262;
  assign tmp35554 = s8 ? tmp35262 : tmp35023;
  assign tmp35549 = s9 ? tmp35550 : tmp35554;
  assign tmp35557 = s7 ? tmp35552 : tmp35058;
  assign tmp35556 = s8 ? tmp35557 : tmp35263;
  assign tmp35555 = s9 ? tmp35278 : tmp35556;
  assign tmp35548 = s10 ? tmp35549 : tmp35555;
  assign tmp35561 = s7 ? tmp35552 : tmp35024;
  assign tmp35560 = s8 ? tmp35561 : tmp35263;
  assign tmp35559 = s9 ? tmp35278 : tmp35560;
  assign tmp35558 = s10 ? tmp35549 : tmp35559;
  assign tmp35547 = s11 ? tmp35548 : tmp35558;
  assign tmp35499 = s12 ? tmp35500 : tmp35547;
  assign tmp35430 = s13 ? tmp35431 : tmp35499;
  assign tmp35330 = s14 ? tmp35331 : tmp35430;
  assign tmp35571 = s5 ? tmp35178 : tmp35265;
  assign tmp35570 = s6 ? tmp34966 : tmp35571;
  assign tmp35569 = s7 ? tmp33914 : tmp35570;
  assign tmp35568 = s8 ? tmp35569 : tmp35262;
  assign tmp35572 = s8 ? tmp35262 : tmp35195;
  assign tmp35567 = s9 ? tmp35568 : tmp35572;
  assign tmp35577 = s5 ? tmp35220 : tmp35265;
  assign tmp35576 = s6 ? tmp34966 : tmp35577;
  assign tmp35575 = s7 ? tmp35576 : tmp35226;
  assign tmp35574 = s8 ? tmp35575 : tmp35263;
  assign tmp35573 = s9 ? tmp35278 : tmp35574;
  assign tmp35566 = s10 ? tmp35567 : tmp35573;
  assign tmp35581 = s7 ? tmp35570 : tmp35196;
  assign tmp35580 = s8 ? tmp35581 : tmp35263;
  assign tmp35579 = s9 ? tmp35278 : tmp35580;
  assign tmp35578 = s10 ? tmp35567 : tmp35579;
  assign tmp35565 = s11 ? tmp35566 : tmp35578;
  assign tmp35587 = s5 ? tmp35015 : tmp35255;
  assign tmp35586 = s6 ? tmp34996 : tmp35587;
  assign tmp35585 = s7 ? tmp33914 : tmp35586;
  assign tmp35584 = s8 ? tmp35238 : tmp35585;
  assign tmp35583 = s9 ? tmp35584 : tmp35585;
  assign tmp35589 = s8 ? tmp35585 : tmp33914;
  assign tmp35597 = s0 ? tmp35004 : tmp34878;
  assign tmp35596 = s1 ? tmp34877 : tmp35597;
  assign tmp35598 = s1 ? tmp35006 : tmp34878;
  assign tmp35595 = ~(s2 ? tmp35596 : tmp35598);
  assign tmp35594 = s3 ? tmp35027 : tmp35595;
  assign tmp35593 = s4 ? tmp35594 : tmp35037;
  assign tmp35603 = s1 ? tmp35049 : tmp34053;
  assign tmp35602 = s2 ? tmp35603 : tmp34904;
  assign tmp35605 = s1 ? tmp35004 : tmp34910;
  assign tmp35604 = ~(s2 ? tmp35605 : tmp34911);
  assign tmp35601 = s3 ? tmp35602 : tmp35604;
  assign tmp35600 = s4 ? tmp35601 : tmp34915;
  assign tmp35610 = l1 ? tmp34056 : tmp33939;
  assign tmp35609 = s1 ? tmp34052 : tmp35610;
  assign tmp35608 = s2 ? tmp34926 : tmp35609;
  assign tmp35607 = s3 ? tmp35608 : tmp35276;
  assign tmp35612 = s1 ? tmp34085 : tmp34936;
  assign tmp35611 = s3 ? tmp34951 : tmp35612;
  assign tmp35606 = s4 ? tmp35607 : tmp35611;
  assign tmp35599 = s5 ? tmp35600 : tmp35606;
  assign tmp35592 = s6 ? tmp35593 : tmp35599;
  assign tmp35591 = s7 ? tmp35239 : tmp35592;
  assign tmp35590 = s8 ? tmp35591 : tmp35586;
  assign tmp35588 = s9 ? tmp35589 : tmp35590;
  assign tmp35582 = s10 ? tmp35583 : tmp35588;
  assign tmp35564 = s12 ? tmp35565 : tmp35582;
  assign tmp35563 = s13 ? tmp35564 : tmp35281;
  assign tmp35562 = s14 ? tmp35067 : tmp35563;
  assign tmp35329 = s15 ? tmp35330 : tmp35562;
  assign tmp33905 = s16 ? tmp33906 : tmp35329;
  assign tmp35620 = s8 ? tmp35336 : tmp34220;
  assign tmp35619 = s9 ? tmp35335 : tmp35620;
  assign tmp35623 = s7 ? tmp35359 : tmp34310;
  assign tmp35622 = s8 ? tmp34349 : tmp35623;
  assign tmp35621 = s9 ? tmp34308 : tmp35622;
  assign tmp35618 = s10 ? tmp35619 : tmp35621;
  assign tmp35627 = s7 ? tmp35337 : tmp34310;
  assign tmp35626 = s8 ? tmp34360 : tmp35627;
  assign tmp35625 = s9 ? tmp34308 : tmp35626;
  assign tmp35624 = s10 ? tmp35619 : tmp35625;
  assign tmp35617 = s11 ? tmp35618 : tmp35624;
  assign tmp35632 = s8 ? tmp35381 : tmp34599;
  assign tmp35631 = s9 ? tmp35380 : tmp35632;
  assign tmp35635 = s7 ? tmp35423 : tmp34627;
  assign tmp35634 = s8 ? tmp34639 : tmp35635;
  assign tmp35633 = s9 ? tmp34625 : tmp35634;
  assign tmp35630 = s10 ? tmp35631 : tmp35633;
  assign tmp35639 = s7 ? tmp35382 : tmp34627;
  assign tmp35638 = s8 ? tmp34647 : tmp35639;
  assign tmp35637 = s9 ? tmp34625 : tmp35638;
  assign tmp35636 = s10 ? tmp35631 : tmp35637;
  assign tmp35629 = s11 ? tmp35630 : tmp35636;
  assign tmp35628 = s12 ? tmp34362 : tmp35629;
  assign tmp35616 = s13 ? tmp35617 : tmp35628;
  assign tmp35644 = s8 ? tmp35434 : tmp34672;
  assign tmp35643 = s9 ? tmp35434 : tmp35644;
  assign tmp35647 = s7 ? tmp35435 : tmp34667;
  assign tmp35646 = s8 ? tmp34689 : tmp35647;
  assign tmp35645 = s9 ? tmp34687 : tmp35646;
  assign tmp35642 = s10 ? tmp35643 : tmp35645;
  assign tmp35652 = s7 ? tmp33914 : tmp34752;
  assign tmp35651 = s8 ? tmp35466 : tmp35652;
  assign tmp35650 = s9 ? tmp35466 : tmp35651;
  assign tmp35654 = s7 ? tmp35493 : tmp34730;
  assign tmp35653 = s9 ? tmp34745 : tmp35654;
  assign tmp35649 = s10 ? tmp35650 : tmp35653;
  assign tmp35657 = s7 ? tmp35467 : tmp34730;
  assign tmp35656 = s9 ? tmp34745 : tmp35657;
  assign tmp35655 = s10 ? tmp35650 : tmp35656;
  assign tmp35648 = s11 ? tmp35649 : tmp35655;
  assign tmp35641 = s12 ? tmp35642 : tmp35648;
  assign tmp35662 = s8 ? tmp34763 : tmp35511;
  assign tmp35663 = s8 ? tmp35511 : tmp34867;
  assign tmp35661 = s9 ? tmp35662 : tmp35663;
  assign tmp35668 = s5 ? tmp34835 : tmp34943;
  assign tmp35667 = s6 ? tmp34803 : tmp35668;
  assign tmp35666 = s7 ? tmp35667 : tmp34953;
  assign tmp35665 = s8 ? tmp34940 : tmp35666;
  assign tmp35664 = s9 ? tmp34938 : tmp35665;
  assign tmp35660 = s10 ? tmp35661 : tmp35664;
  assign tmp35672 = s7 ? tmp35512 : tmp34802;
  assign tmp35671 = s8 ? tmp34959 : tmp35672;
  assign tmp35670 = s9 ? tmp34938 : tmp35671;
  assign tmp35669 = s10 ? tmp35661 : tmp35670;
  assign tmp35659 = s11 ? tmp35660 : tmp35669;
  assign tmp35658 = s12 ? tmp35659 : tmp34960;
  assign tmp35640 = s13 ? tmp35641 : tmp35658;
  assign tmp35615 = s14 ? tmp35616 : tmp35640;
  assign tmp35678 = s8 ? tmp35585 : tmp35268;
  assign tmp35677 = s9 ? tmp35584 : tmp35678;
  assign tmp35680 = s8 ? tmp35280 : tmp35586;
  assign tmp35679 = s9 ? tmp35278 : tmp35680;
  assign tmp35676 = s10 ? tmp35677 : tmp35679;
  assign tmp35675 = s12 ? tmp35171 : tmp35676;
  assign tmp35674 = s13 ? tmp35675 : tmp35281;
  assign tmp35673 = s14 ? tmp35067 : tmp35674;
  assign tmp35614 = s15 ? tmp35615 : tmp35673;
  assign tmp35687 = s9 ? tmp35662 : tmp35511;
  assign tmp35689 = s8 ? tmp35511 : tmp33914;
  assign tmp35691 = s7 ? tmp34941 : tmp35518;
  assign tmp35690 = s8 ? tmp35691 : tmp35667;
  assign tmp35688 = s9 ? tmp35689 : tmp35690;
  assign tmp35686 = s10 ? tmp35687 : tmp35688;
  assign tmp35695 = s7 ? tmp34764 : tmp35543;
  assign tmp35694 = s8 ? tmp35695 : tmp35512;
  assign tmp35693 = s9 ? tmp35689 : tmp35694;
  assign tmp35692 = s10 ? tmp35687 : tmp35693;
  assign tmp35685 = s11 ? tmp35686 : tmp35692;
  assign tmp35684 = s12 ? tmp35685 : tmp34960;
  assign tmp35683 = s13 ? tmp35431 : tmp35684;
  assign tmp35682 = s14 ? tmp35331 : tmp35683;
  assign tmp35698 = s12 ? tmp35171 : tmp35582;
  assign tmp35697 = s13 ? tmp35698 : tmp35281;
  assign tmp35696 = s14 ? tmp35067 : tmp35697;
  assign tmp35681 = s15 ? tmp35682 : tmp35696;
  assign tmp35613 = s16 ? tmp35614 : tmp35681;
  assign tmp33904 = ~(s17 ? tmp33905 : tmp35613);
  assign s3n = tmp33904;

  assign tmp35716 = l4 ? 1 : 0;
  assign tmp35717 = ~(l4 ? 1 : 0);
  assign tmp35715 = l3 ? tmp35716 : tmp35717;
  assign tmp35714 = l2 ? 1 : tmp35715;
  assign tmp35719 = l3 ? 1 : 0;
  assign tmp35720 = ~(l3 ? 1 : 0);
  assign tmp35718 = l2 ? tmp35719 : tmp35720;
  assign tmp35713 = l1 ? tmp35714 : tmp35718;
  assign tmp35724 = l3 ? 1 : tmp35717;
  assign tmp35725 = ~(l3 ? tmp35716 : 0);
  assign tmp35723 = l2 ? tmp35724 : tmp35725;
  assign tmp35727 = l3 ? tmp35716 : 0;
  assign tmp35726 = ~(l2 ? tmp35727 : 0);
  assign tmp35722 = l1 ? tmp35723 : tmp35726;
  assign tmp35730 = ~(l3 ? tmp35716 : tmp35717);
  assign tmp35729 = l2 ? tmp35719 : tmp35730;
  assign tmp35731 = ~(l2 ? tmp35727 : tmp35720);
  assign tmp35728 = l1 ? tmp35729 : tmp35731;
  assign tmp35721 = ~(s0 ? tmp35722 : tmp35728);
  assign tmp35712 = s1 ? tmp35713 : tmp35721;
  assign tmp35736 = l2 ? 1 : tmp35724;
  assign tmp35737 = ~(l2 ? tmp35716 : tmp35727);
  assign tmp35735 = l1 ? tmp35736 : tmp35737;
  assign tmp35739 = l2 ? tmp35727 : tmp35730;
  assign tmp35740 = l2 ? 1 : tmp35719;
  assign tmp35738 = ~(l1 ? tmp35739 : tmp35740);
  assign tmp35734 = s0 ? tmp35735 : tmp35738;
  assign tmp35743 = l2 ? tmp35719 : tmp35725;
  assign tmp35745 = ~(l3 ? 1 : tmp35717);
  assign tmp35744 = ~(l2 ? tmp35727 : tmp35745);
  assign tmp35742 = l1 ? tmp35743 : tmp35744;
  assign tmp35746 = l1 ? tmp35739 : tmp35740;
  assign tmp35741 = ~(s0 ? tmp35742 : tmp35746);
  assign tmp35733 = s1 ? tmp35734 : tmp35741;
  assign tmp35749 = l1 ? tmp35723 : 1;
  assign tmp35748 = s0 ? tmp35742 : tmp35749;
  assign tmp35751 = ~(l1 ? tmp35714 : tmp35718);
  assign tmp35750 = s0 ? tmp35746 : tmp35751;
  assign tmp35747 = ~(s1 ? tmp35748 : tmp35750);
  assign tmp35732 = s2 ? tmp35733 : tmp35747;
  assign tmp35711 = s3 ? tmp35712 : tmp35732;
  assign tmp35756 = l1 ? tmp35743 : tmp35731;
  assign tmp35757 = ~(l1 ? tmp35736 : tmp35725);
  assign tmp35755 = s0 ? tmp35756 : tmp35757;
  assign tmp35758 = ~(s0 ? tmp35713 : tmp35738);
  assign tmp35754 = s1 ? tmp35755 : tmp35758;
  assign tmp35761 = ~(l1 ? tmp35723 : 1);
  assign tmp35760 = s0 ? tmp35713 : tmp35761;
  assign tmp35765 = l3 ? tmp35716 : 1;
  assign tmp35764 = ~(l2 ? tmp35765 : 0);
  assign tmp35763 = l1 ? tmp35736 : tmp35764;
  assign tmp35767 = l2 ? tmp35724 : 1;
  assign tmp35768 = l2 ? 1 : tmp35725;
  assign tmp35766 = ~(l1 ? tmp35767 : tmp35768);
  assign tmp35762 = s0 ? tmp35763 : tmp35766;
  assign tmp35759 = ~(s1 ? tmp35760 : tmp35762);
  assign tmp35753 = s2 ? tmp35754 : tmp35759;
  assign tmp35773 = l2 ? 1 : tmp35717;
  assign tmp35772 = l1 ? tmp35773 : tmp35726;
  assign tmp35771 = s0 ? tmp35772 : tmp35761;
  assign tmp35775 = l1 ? tmp35767 : tmp35768;
  assign tmp35778 = l3 ? 1 : tmp35716;
  assign tmp35777 = l2 ? tmp35765 : tmp35778;
  assign tmp35779 = l2 ? 1 : tmp35778;
  assign tmp35776 = l1 ? tmp35777 : tmp35779;
  assign tmp35774 = ~(s0 ? tmp35775 : tmp35776);
  assign tmp35770 = s1 ? tmp35771 : tmp35774;
  assign tmp35783 = ~(l2 ? 1 : tmp35719);
  assign tmp35782 = ~(l1 ? tmp35714 : tmp35783);
  assign tmp35781 = s0 ? tmp35746 : tmp35782;
  assign tmp35786 = l2 ? tmp35716 : tmp35778;
  assign tmp35785 = l1 ? tmp35786 : tmp35779;
  assign tmp35784 = s0 ? tmp35785 : tmp35746;
  assign tmp35780 = ~(s1 ? tmp35781 : tmp35784);
  assign tmp35769 = ~(s2 ? tmp35770 : tmp35780);
  assign tmp35752 = ~(s3 ? tmp35753 : tmp35769);
  assign tmp35710 = s4 ? tmp35711 : tmp35752;
  assign tmp35793 = ~(l1 ? 1 : tmp35725);
  assign tmp35792 = s0 ? tmp35728 : tmp35793;
  assign tmp35795 = l1 ? tmp35768 : tmp35726;
  assign tmp35794 = ~(s0 ? tmp35795 : tmp35735);
  assign tmp35791 = s1 ? tmp35792 : tmp35794;
  assign tmp35798 = l1 ? tmp35714 : tmp35764;
  assign tmp35797 = s0 ? tmp35795 : tmp35798;
  assign tmp35800 = l1 ? tmp35714 : tmp35783;
  assign tmp35801 = l1 ? 1 : tmp35737;
  assign tmp35799 = s0 ? tmp35800 : tmp35801;
  assign tmp35796 = ~(s1 ? tmp35797 : tmp35799);
  assign tmp35790 = s2 ? tmp35791 : tmp35796;
  assign tmp35806 = l2 ? tmp35719 : 1;
  assign tmp35805 = ~(l1 ? tmp35806 : tmp35744);
  assign tmp35804 = s0 ? 1 : tmp35805;
  assign tmp35808 = ~(l1 ? tmp35786 : tmp35740);
  assign tmp35807 = s0 ? 1 : tmp35808;
  assign tmp35803 = s1 ? tmp35804 : tmp35807;
  assign tmp35812 = l2 ? 1 : tmp35765;
  assign tmp35811 = ~(l1 ? tmp35812 : tmp35765);
  assign tmp35810 = s0 ? tmp35785 : tmp35811;
  assign tmp35815 = l2 ? tmp35727 : tmp35778;
  assign tmp35814 = l1 ? tmp35815 : tmp35740;
  assign tmp35813 = s0 ? tmp35746 : tmp35814;
  assign tmp35809 = ~(s1 ? tmp35810 : tmp35813);
  assign tmp35802 = ~(s2 ? tmp35803 : tmp35809);
  assign tmp35789 = s3 ? tmp35790 : tmp35802;
  assign tmp35821 = l2 ? tmp35765 : 1;
  assign tmp35820 = l1 ? tmp35821 : tmp35779;
  assign tmp35819 = s0 ? tmp35820 : tmp35746;
  assign tmp35823 = l1 ? tmp35736 : tmp35726;
  assign tmp35824 = l1 ? tmp35736 : tmp35806;
  assign tmp35822 = ~(s0 ? tmp35823 : tmp35824);
  assign tmp35818 = s1 ? tmp35819 : tmp35822;
  assign tmp35827 = l1 ? tmp35736 : 1;
  assign tmp35826 = s0 ? tmp35772 : tmp35827;
  assign tmp35828 = s0 ? tmp35763 : tmp35772;
  assign tmp35825 = ~(s1 ? tmp35826 : tmp35828);
  assign tmp35817 = s2 ? tmp35818 : tmp35825;
  assign tmp35833 = l2 ? tmp35778 : 1;
  assign tmp35832 = l1 ? tmp35833 : tmp35740;
  assign tmp35835 = l2 ? tmp35727 : 1;
  assign tmp35834 = l1 ? tmp35835 : tmp35740;
  assign tmp35831 = s0 ? tmp35832 : tmp35834;
  assign tmp35838 = l2 ? tmp35716 : tmp35765;
  assign tmp35837 = l1 ? tmp35714 : tmp35838;
  assign tmp35836 = ~(s0 ? tmp35827 : tmp35837);
  assign tmp35830 = s1 ? tmp35831 : tmp35836;
  assign tmp35841 = l1 ? tmp35821 : 1;
  assign tmp35842 = l1 ? 1 : tmp35812;
  assign tmp35840 = s0 ? tmp35841 : tmp35842;
  assign tmp35843 = s0 ? tmp35776 : tmp35842;
  assign tmp35839 = s1 ? tmp35840 : tmp35843;
  assign tmp35829 = s2 ? tmp35830 : tmp35839;
  assign tmp35816 = s3 ? tmp35817 : tmp35829;
  assign tmp35788 = s4 ? tmp35789 : tmp35816;
  assign tmp35849 = l1 ? tmp35786 : tmp35740;
  assign tmp35850 = ~(l1 ? tmp35812 : tmp35821);
  assign tmp35848 = s0 ? tmp35849 : tmp35850;
  assign tmp35852 = l1 ? tmp35765 : tmp35821;
  assign tmp35853 = l1 ? tmp35812 : tmp35806;
  assign tmp35851 = ~(s0 ? tmp35852 : tmp35853);
  assign tmp35847 = s1 ? tmp35848 : tmp35851;
  assign tmp35857 = l2 ? tmp35778 : tmp35765;
  assign tmp35856 = l1 ? tmp35857 : 1;
  assign tmp35858 = ~(l1 ? tmp35833 : tmp35736);
  assign tmp35855 = s0 ? tmp35856 : tmp35858;
  assign tmp35860 = ~(l1 ? 1 : tmp35767);
  assign tmp35859 = s0 ? tmp35827 : tmp35860;
  assign tmp35854 = ~(s1 ? tmp35855 : tmp35859);
  assign tmp35846 = s2 ? tmp35847 : tmp35854;
  assign tmp35865 = l2 ? tmp35778 : tmp35724;
  assign tmp35864 = l1 ? tmp35865 : tmp35736;
  assign tmp35863 = s0 ? tmp35864 : tmp35842;
  assign tmp35867 = ~(l1 ? tmp35779 : 1);
  assign tmp35866 = s0 ? tmp35779 : tmp35867;
  assign tmp35862 = s1 ? tmp35863 : tmp35866;
  assign tmp35870 = ~(l1 ? tmp35812 : tmp35857);
  assign tmp35869 = s0 ? tmp35842 : tmp35870;
  assign tmp35872 = l1 ? tmp35765 : tmp35779;
  assign tmp35873 = ~(l1 ? tmp35833 : tmp35740);
  assign tmp35871 = ~(s0 ? tmp35872 : tmp35873);
  assign tmp35868 = ~(s1 ? tmp35869 : tmp35871);
  assign tmp35861 = ~(s2 ? tmp35862 : tmp35868);
  assign tmp35845 = s3 ? tmp35846 : tmp35861;
  assign tmp35878 = l1 ? 1 : tmp35833;
  assign tmp35879 = ~(l1 ? tmp35812 : 1);
  assign tmp35877 = s0 ? tmp35878 : tmp35879;
  assign tmp35882 = l2 ? tmp35778 : tmp35716;
  assign tmp35881 = l1 ? tmp35882 : tmp35779;
  assign tmp35883 = ~(l1 ? tmp35786 : tmp35779);
  assign tmp35880 = ~(s0 ? tmp35881 : tmp35883);
  assign tmp35876 = s1 ? tmp35877 : tmp35880;
  assign tmp35885 = s0 ? tmp35852 : tmp35798;
  assign tmp35887 = l1 ? 1 : tmp35767;
  assign tmp35888 = ~(l1 ? tmp35865 : tmp35736);
  assign tmp35886 = ~(s0 ? tmp35887 : tmp35888);
  assign tmp35884 = ~(s1 ? tmp35885 : tmp35886);
  assign tmp35875 = s2 ? tmp35876 : tmp35884;
  assign tmp35892 = l1 ? tmp35812 : tmp35765;
  assign tmp35891 = s0 ? tmp35856 : tmp35892;
  assign tmp35894 = ~(l1 ? tmp35714 : tmp35857);
  assign tmp35893 = ~(s0 ? tmp35842 : tmp35894);
  assign tmp35890 = s1 ? tmp35891 : tmp35893;
  assign tmp35897 = ~(l1 ? 1 : tmp35833);
  assign tmp35896 = s0 ? tmp35872 : tmp35897;
  assign tmp35898 = s0 ? tmp35779 : tmp35881;
  assign tmp35895 = s1 ? tmp35896 : tmp35898;
  assign tmp35889 = ~(s2 ? tmp35890 : tmp35895);
  assign tmp35874 = s3 ? tmp35875 : tmp35889;
  assign tmp35844 = s4 ? tmp35845 : tmp35874;
  assign tmp35787 = ~(s5 ? tmp35788 : tmp35844);
  assign tmp35709 = s6 ? tmp35710 : tmp35787;
  assign tmp35904 = l2 ? tmp35719 : tmp35715;
  assign tmp35903 = l1 ? tmp35904 : tmp35768;
  assign tmp35906 = l1 ? tmp35723 : tmp35764;
  assign tmp35908 = l2 ? 1 : tmp35730;
  assign tmp35909 = ~(l2 ? tmp35765 : tmp35720);
  assign tmp35907 = l1 ? tmp35908 : tmp35909;
  assign tmp35905 = ~(s0 ? tmp35906 : tmp35907);
  assign tmp35902 = s1 ? tmp35903 : tmp35905;
  assign tmp35914 = l2 ? tmp35719 : tmp35724;
  assign tmp35913 = l1 ? tmp35914 : tmp35737;
  assign tmp35916 = l2 ? tmp35715 : tmp35730;
  assign tmp35917 = l2 ? tmp35778 : tmp35727;
  assign tmp35915 = ~(l1 ? tmp35916 : tmp35917);
  assign tmp35912 = s0 ? tmp35913 : tmp35915;
  assign tmp35920 = ~(l2 ? tmp35765 : tmp35745);
  assign tmp35919 = l1 ? tmp35768 : tmp35920;
  assign tmp35921 = l1 ? tmp35916 : tmp35917;
  assign tmp35918 = ~(s0 ? tmp35919 : tmp35921);
  assign tmp35911 = s1 ? tmp35912 : tmp35918;
  assign tmp35923 = s0 ? tmp35919 : tmp35749;
  assign tmp35926 = l2 ? tmp35778 : tmp35715;
  assign tmp35925 = ~(l1 ? tmp35926 : tmp35768);
  assign tmp35924 = s0 ? tmp35921 : tmp35925;
  assign tmp35922 = ~(s1 ? tmp35923 : tmp35924);
  assign tmp35910 = s2 ? tmp35911 : tmp35922;
  assign tmp35901 = s3 ? tmp35902 : tmp35910;
  assign tmp35931 = l1 ? tmp35768 : tmp35909;
  assign tmp35930 = s0 ? tmp35931 : tmp35757;
  assign tmp35933 = l1 ? tmp35926 : tmp35768;
  assign tmp35932 = ~(s0 ? tmp35933 : tmp35915);
  assign tmp35929 = s1 ? tmp35930 : tmp35932;
  assign tmp35935 = s0 ? tmp35903 : tmp35761;
  assign tmp35934 = ~(s1 ? tmp35935 : tmp35823);
  assign tmp35928 = s2 ? tmp35929 : tmp35934;
  assign tmp35938 = l1 ? tmp35777 : tmp35882;
  assign tmp35937 = s1 ? tmp35906 : tmp35938;
  assign tmp35942 = ~(l2 ? tmp35778 : tmp35727);
  assign tmp35941 = ~(l1 ? tmp35926 : tmp35942);
  assign tmp35940 = s0 ? tmp35921 : tmp35941;
  assign tmp35945 = l2 ? tmp35719 : tmp35716;
  assign tmp35944 = l1 ? tmp35777 : tmp35945;
  assign tmp35943 = s0 ? tmp35944 : tmp35921;
  assign tmp35939 = s1 ? tmp35940 : tmp35943;
  assign tmp35936 = s2 ? tmp35937 : tmp35939;
  assign tmp35927 = ~(s3 ? tmp35928 : tmp35936);
  assign tmp35900 = s4 ? tmp35901 : tmp35927;
  assign tmp35951 = s0 ? tmp35907 : tmp35793;
  assign tmp35952 = ~(l1 ? tmp35914 : tmp35737);
  assign tmp35950 = s1 ? tmp35951 : tmp35952;
  assign tmp35955 = ~(l2 ? tmp35716 : 0);
  assign tmp35954 = l1 ? tmp35904 : tmp35955;
  assign tmp35957 = l1 ? tmp35926 : tmp35942;
  assign tmp35956 = s0 ? tmp35957 : tmp35801;
  assign tmp35953 = ~(s1 ? tmp35954 : tmp35956);
  assign tmp35949 = s2 ? tmp35950 : tmp35953;
  assign tmp35960 = l1 ? 1 : tmp35920;
  assign tmp35961 = l1 ? tmp35777 : tmp35917;
  assign tmp35959 = s1 ? tmp35960 : tmp35961;
  assign tmp35963 = s0 ? tmp35944 : tmp35850;
  assign tmp35966 = l2 ? tmp35715 : tmp35778;
  assign tmp35965 = l1 ? tmp35966 : tmp35917;
  assign tmp35964 = s0 ? tmp35921 : tmp35965;
  assign tmp35962 = s1 ? tmp35963 : tmp35964;
  assign tmp35958 = s2 ? tmp35959 : tmp35962;
  assign tmp35948 = s3 ? tmp35949 : tmp35958;
  assign tmp35971 = l1 ? tmp35821 : tmp35882;
  assign tmp35973 = l2 ? tmp35719 : tmp35727;
  assign tmp35972 = l1 ? tmp35916 : tmp35973;
  assign tmp35970 = s0 ? tmp35971 : tmp35972;
  assign tmp35974 = ~(s0 ? tmp35823 : tmp35827);
  assign tmp35969 = s1 ? tmp35970 : tmp35974;
  assign tmp35977 = l1 ? tmp35914 : tmp35955;
  assign tmp35976 = s0 ? tmp35977 : tmp35772;
  assign tmp35975 = ~(s1 ? tmp35772 : tmp35976);
  assign tmp35968 = s2 ? tmp35969 : tmp35975;
  assign tmp35982 = l2 ? tmp35778 : tmp35719;
  assign tmp35981 = l1 ? 1 : tmp35982;
  assign tmp35983 = l1 ? tmp35821 : tmp35973;
  assign tmp35980 = s0 ? tmp35981 : tmp35983;
  assign tmp35984 = ~(l1 ? tmp35926 : tmp35821);
  assign tmp35979 = s1 ? tmp35980 : tmp35984;
  assign tmp35986 = l1 ? tmp35821 : tmp35812;
  assign tmp35985 = s1 ? tmp35986 : tmp35938;
  assign tmp35978 = s2 ? tmp35979 : tmp35985;
  assign tmp35967 = s3 ? tmp35968 : tmp35978;
  assign tmp35947 = s4 ? tmp35948 : tmp35967;
  assign tmp35991 = s0 ? tmp35961 : tmp35850;
  assign tmp35992 = ~(l1 ? tmp35857 : 1);
  assign tmp35990 = s1 ? tmp35991 : tmp35992;
  assign tmp35994 = l1 ? 1 : tmp35736;
  assign tmp35995 = ~(l1 ? tmp35865 : 1);
  assign tmp35993 = s1 ? tmp35994 : tmp35995;
  assign tmp35989 = s2 ? tmp35990 : tmp35993;
  assign tmp35998 = ~(l1 ? tmp35779 : tmp35812);
  assign tmp35997 = s1 ? 1 : tmp35998;
  assign tmp36000 = l1 ? tmp35812 : 1;
  assign tmp36001 = ~(l1 ? 1 : tmp35982);
  assign tmp35999 = s1 ? tmp36000 : tmp36001;
  assign tmp35996 = ~(s2 ? tmp35997 : tmp35999);
  assign tmp35988 = s3 ? tmp35989 : tmp35996;
  assign tmp36005 = ~(l1 ? tmp35777 : tmp35945);
  assign tmp36004 = s1 ? tmp35856 : tmp36005;
  assign tmp36006 = l1 ? tmp35926 : tmp35955;
  assign tmp36003 = s2 ? tmp36004 : tmp36006;
  assign tmp36008 = l1 ? tmp35857 : tmp35821;
  assign tmp36009 = l1 ? tmp35926 : 1;
  assign tmp36007 = s1 ? tmp36008 : tmp36009;
  assign tmp36002 = ~(s3 ? tmp36003 : tmp36007);
  assign tmp35987 = s4 ? tmp35988 : tmp36002;
  assign tmp35946 = ~(s5 ? tmp35947 : tmp35987);
  assign tmp35899 = s6 ? tmp35900 : tmp35946;
  assign tmp35708 = s7 ? tmp35709 : tmp35899;
  assign tmp36017 = l2 ? tmp35724 : tmp35730;
  assign tmp36016 = l1 ? tmp36017 : tmp35909;
  assign tmp36015 = ~(s0 ? tmp35906 : tmp36016);
  assign tmp36014 = s1 ? tmp35933 : tmp36015;
  assign tmp36021 = l1 ? tmp35865 : tmp35725;
  assign tmp36022 = ~(l1 ? tmp35916 : tmp35973);
  assign tmp36020 = s0 ? tmp36021 : tmp36022;
  assign tmp36024 = l1 ? tmp35723 : tmp35920;
  assign tmp36023 = ~(s0 ? tmp36024 : tmp35972);
  assign tmp36019 = s1 ? tmp36020 : tmp36023;
  assign tmp36027 = l1 ? tmp35723 : tmp35767;
  assign tmp36026 = s0 ? tmp36024 : tmp36027;
  assign tmp36028 = s0 ? tmp35972 : tmp35925;
  assign tmp36025 = ~(s1 ? tmp36026 : tmp36028);
  assign tmp36018 = s2 ? tmp36019 : tmp36025;
  assign tmp36013 = s3 ? tmp36014 : tmp36018;
  assign tmp36033 = l1 ? tmp35723 : tmp35909;
  assign tmp36032 = s0 ? tmp36033 : tmp35757;
  assign tmp36034 = ~(s0 ? tmp35933 : tmp36022);
  assign tmp36031 = s1 ? tmp36032 : tmp36034;
  assign tmp36036 = s0 ? tmp35933 : tmp35761;
  assign tmp36035 = ~(s1 ? tmp36036 : tmp35823);
  assign tmp36030 = s2 ? tmp36031 : tmp36035;
  assign tmp36041 = ~(l2 ? tmp35719 : tmp35727);
  assign tmp36040 = ~(l1 ? tmp35926 : tmp36041);
  assign tmp36039 = s0 ? tmp35972 : tmp36040;
  assign tmp36042 = s0 ? tmp35944 : tmp35972;
  assign tmp36038 = s1 ? tmp36039 : tmp36042;
  assign tmp36037 = s2 ? tmp35937 : tmp36038;
  assign tmp36029 = ~(s3 ? tmp36030 : tmp36037);
  assign tmp36012 = s4 ? tmp36013 : tmp36029;
  assign tmp36048 = s0 ? tmp36016 : tmp35793;
  assign tmp36049 = ~(l1 ? tmp35865 : tmp35725);
  assign tmp36047 = s1 ? tmp36048 : tmp36049;
  assign tmp36051 = l1 ? tmp35926 : tmp35726;
  assign tmp36053 = l1 ? tmp35926 : tmp36041;
  assign tmp36054 = l1 ? 1 : tmp35725;
  assign tmp36052 = s0 ? tmp36053 : tmp36054;
  assign tmp36050 = ~(s1 ? tmp36051 : tmp36052);
  assign tmp36046 = s2 ? tmp36047 : tmp36050;
  assign tmp36057 = l1 ? tmp35767 : tmp35920;
  assign tmp36058 = l1 ? tmp35777 : tmp35973;
  assign tmp36056 = s1 ? tmp36057 : tmp36058;
  assign tmp36061 = l1 ? tmp35966 : tmp35973;
  assign tmp36060 = s0 ? tmp35972 : tmp36061;
  assign tmp36059 = s1 ? tmp35963 : tmp36060;
  assign tmp36055 = s2 ? tmp36056 : tmp36059;
  assign tmp36045 = s3 ? tmp36046 : tmp36055;
  assign tmp36064 = ~(l1 ? tmp35865 : tmp35726);
  assign tmp36063 = s2 ? tmp35969 : tmp36064;
  assign tmp36068 = l1 ? 1 : tmp35719;
  assign tmp36070 = l2 ? tmp35715 : 1;
  assign tmp36069 = l1 ? tmp36070 : tmp35973;
  assign tmp36067 = s0 ? tmp36068 : tmp36069;
  assign tmp36066 = s1 ? tmp36067 : tmp35984;
  assign tmp36065 = s2 ? tmp36066 : tmp35985;
  assign tmp36062 = s3 ? tmp36063 : tmp36065;
  assign tmp36044 = s4 ? tmp36045 : tmp36062;
  assign tmp36075 = s0 ? tmp36058 : tmp35850;
  assign tmp36074 = s1 ? tmp36075 : tmp35992;
  assign tmp36077 = l1 ? 1 : tmp35724;
  assign tmp36076 = s1 ? tmp36077 : tmp35995;
  assign tmp36073 = s2 ? tmp36074 : tmp36076;
  assign tmp36072 = s3 ? tmp36073 : tmp35996;
  assign tmp36079 = s2 ? tmp36004 : tmp36051;
  assign tmp36078 = ~(s3 ? tmp36079 : tmp36007);
  assign tmp36071 = s4 ? tmp36072 : tmp36078;
  assign tmp36043 = ~(s5 ? tmp36044 : tmp36071);
  assign tmp36011 = s6 ? tmp36012 : tmp36043;
  assign tmp36010 = s7 ? tmp35709 : tmp36011;
  assign tmp35707 = s8 ? tmp35708 : tmp36010;
  assign tmp36086 = l1 ? tmp35904 : tmp35773;
  assign tmp36088 = l1 ? tmp35768 : tmp35764;
  assign tmp36091 = ~(l3 ? 1 : tmp35716);
  assign tmp36090 = ~(l2 ? tmp35765 : tmp36091);
  assign tmp36089 = l1 ? tmp35908 : tmp36090;
  assign tmp36087 = ~(s0 ? tmp36088 : tmp36089);
  assign tmp36085 = s1 ? tmp36086 : tmp36087;
  assign tmp36096 = ~(l2 ? tmp35727 : tmp35716);
  assign tmp36095 = l1 ? tmp35914 : tmp36096;
  assign tmp36098 = l2 ? tmp35765 : tmp35730;
  assign tmp36097 = ~(l1 ? tmp36098 : tmp35945);
  assign tmp36094 = s0 ? tmp36095 : tmp36097;
  assign tmp36100 = l1 ? tmp36098 : tmp35945;
  assign tmp36099 = ~(s0 ? tmp36088 : tmp36100);
  assign tmp36093 = s1 ? tmp36094 : tmp36099;
  assign tmp36103 = l1 ? tmp35768 : tmp35767;
  assign tmp36102 = s0 ? tmp36088 : tmp36103;
  assign tmp36105 = ~(l1 ? tmp35904 : tmp35773);
  assign tmp36104 = s0 ? tmp36100 : tmp36105;
  assign tmp36101 = ~(s1 ? tmp36102 : tmp36104);
  assign tmp36092 = s2 ? tmp36093 : tmp36101;
  assign tmp36084 = s3 ? tmp36085 : tmp36092;
  assign tmp36110 = l1 ? tmp35768 : tmp36090;
  assign tmp36111 = ~(l1 ? tmp35724 : tmp35725);
  assign tmp36109 = s0 ? tmp36110 : tmp36111;
  assign tmp36112 = ~(s0 ? tmp36086 : tmp36097);
  assign tmp36108 = s1 ? tmp36109 : tmp36112;
  assign tmp36115 = ~(l1 ? tmp35768 : 1);
  assign tmp36114 = s0 ? tmp36086 : tmp36115;
  assign tmp36116 = l1 ? tmp35724 : tmp35726;
  assign tmp36113 = ~(s1 ? tmp36114 : tmp36116);
  assign tmp36107 = s2 ? tmp36108 : tmp36113;
  assign tmp36118 = s1 ? tmp36088 : tmp35938;
  assign tmp36122 = ~(l2 ? tmp35719 : tmp35716);
  assign tmp36121 = ~(l1 ? tmp35904 : tmp36122);
  assign tmp36120 = s0 ? tmp36100 : tmp36121;
  assign tmp36123 = s0 ? tmp35944 : tmp36100;
  assign tmp36119 = s1 ? tmp36120 : tmp36123;
  assign tmp36117 = s2 ? tmp36118 : tmp36119;
  assign tmp36106 = ~(s3 ? tmp36107 : tmp36117);
  assign tmp36083 = s4 ? tmp36084 : tmp36106;
  assign tmp36129 = s0 ? tmp36089 : tmp35793;
  assign tmp36130 = ~(l1 ? tmp35914 : tmp36096);
  assign tmp36128 = s1 ? tmp36129 : tmp36130;
  assign tmp36132 = l1 ? tmp35904 : tmp35744;
  assign tmp36134 = l1 ? tmp35904 : tmp36122;
  assign tmp36135 = l1 ? tmp35767 : tmp35725;
  assign tmp36133 = s0 ? tmp36134 : tmp36135;
  assign tmp36131 = ~(s1 ? tmp36132 : tmp36133);
  assign tmp36127 = s2 ? tmp36128 : tmp36131;
  assign tmp36138 = l1 ? 1 : tmp35764;
  assign tmp36137 = s1 ? tmp36138 : tmp35944;
  assign tmp36141 = l1 ? tmp36098 : tmp35973;
  assign tmp36140 = s0 ? tmp36141 : tmp36058;
  assign tmp36139 = s1 ? tmp35963 : tmp36140;
  assign tmp36136 = s2 ? tmp36137 : tmp36139;
  assign tmp36126 = s3 ? tmp36127 : tmp36136;
  assign tmp36145 = s0 ? tmp35971 : tmp36100;
  assign tmp36147 = l1 ? tmp35724 : 1;
  assign tmp36146 = ~(s0 ? tmp36116 : tmp36147);
  assign tmp36144 = s1 ? tmp36145 : tmp36146;
  assign tmp36148 = ~(l1 ? tmp35914 : tmp35744);
  assign tmp36143 = s2 ? tmp36144 : tmp36148;
  assign tmp36153 = l2 ? tmp35719 : tmp35778;
  assign tmp36152 = l1 ? 1 : tmp36153;
  assign tmp36154 = l1 ? tmp35821 : tmp35945;
  assign tmp36151 = s0 ? tmp36152 : tmp36154;
  assign tmp36150 = s1 ? tmp36151 : tmp35984;
  assign tmp36149 = s2 ? tmp36150 : tmp35985;
  assign tmp36142 = s3 ? tmp36143 : tmp36149;
  assign tmp36125 = s4 ? tmp36126 : tmp36142;
  assign tmp36158 = s1 ? tmp35963 : tmp35992;
  assign tmp36159 = s1 ? tmp35887 : tmp35995;
  assign tmp36157 = s2 ? tmp36158 : tmp36159;
  assign tmp36162 = ~(l1 ? 1 : tmp35778);
  assign tmp36161 = s1 ? tmp36000 : tmp36162;
  assign tmp36160 = ~(s2 ? tmp35997 : tmp36161);
  assign tmp36156 = s3 ? tmp36157 : tmp36160;
  assign tmp36165 = l1 ? tmp35926 : tmp35744;
  assign tmp36164 = s2 ? tmp36004 : tmp36165;
  assign tmp36167 = l1 ? tmp35926 : tmp35736;
  assign tmp36166 = s1 ? tmp36008 : tmp36167;
  assign tmp36163 = ~(s3 ? tmp36164 : tmp36166);
  assign tmp36155 = s4 ? tmp36156 : tmp36163;
  assign tmp36124 = ~(s5 ? tmp36125 : tmp36155);
  assign tmp36082 = s6 ? tmp36083 : tmp36124;
  assign tmp36081 = s7 ? tmp35709 : tmp36082;
  assign tmp36080 = s8 ? tmp36010 : tmp36081;
  assign tmp35706 = s9 ? tmp35707 : tmp36080;
  assign tmp36175 = ~(s0 ? tmp36088 : tmp35907);
  assign tmp36174 = s1 ? tmp35903 : tmp36175;
  assign tmp36179 = l1 ? tmp35914 : tmp35725;
  assign tmp36180 = ~(l1 ? tmp36098 : tmp35973);
  assign tmp36178 = s0 ? tmp36179 : tmp36180;
  assign tmp36181 = ~(s0 ? tmp35919 : tmp36141);
  assign tmp36177 = s1 ? tmp36178 : tmp36181;
  assign tmp36183 = s0 ? tmp35919 : tmp36103;
  assign tmp36185 = ~(l1 ? tmp35904 : tmp35768);
  assign tmp36184 = s0 ? tmp36141 : tmp36185;
  assign tmp36182 = ~(s1 ? tmp36183 : tmp36184);
  assign tmp36176 = s2 ? tmp36177 : tmp36182;
  assign tmp36173 = s3 ? tmp36174 : tmp36176;
  assign tmp36189 = s0 ? tmp35931 : tmp36111;
  assign tmp36190 = ~(s0 ? tmp35903 : tmp36180);
  assign tmp36188 = s1 ? tmp36189 : tmp36190;
  assign tmp36192 = s0 ? tmp35903 : tmp36115;
  assign tmp36191 = ~(s1 ? tmp36192 : tmp36116);
  assign tmp36187 = s2 ? tmp36188 : tmp36191;
  assign tmp36196 = ~(l1 ? tmp35904 : tmp36041);
  assign tmp36195 = s0 ? tmp36141 : tmp36196;
  assign tmp36197 = s0 ? tmp35944 : tmp36141;
  assign tmp36194 = s1 ? tmp36195 : tmp36197;
  assign tmp36193 = s2 ? tmp36118 : tmp36194;
  assign tmp36186 = ~(s3 ? tmp36187 : tmp36193);
  assign tmp36172 = s4 ? tmp36173 : tmp36186;
  assign tmp36203 = ~(l1 ? tmp35914 : tmp35725);
  assign tmp36202 = s1 ? tmp35951 : tmp36203;
  assign tmp36205 = l1 ? tmp35904 : tmp35726;
  assign tmp36207 = l1 ? tmp35904 : tmp36041;
  assign tmp36206 = s0 ? tmp36207 : tmp36135;
  assign tmp36204 = ~(s1 ? tmp36205 : tmp36206);
  assign tmp36201 = s2 ? tmp36202 : tmp36204;
  assign tmp36209 = s1 ? tmp35960 : tmp36058;
  assign tmp36208 = s2 ? tmp36209 : tmp36139;
  assign tmp36200 = s3 ? tmp36201 : tmp36208;
  assign tmp36213 = s0 ? tmp35971 : tmp36141;
  assign tmp36212 = s1 ? tmp36213 : tmp36146;
  assign tmp36214 = ~(l1 ? tmp35914 : tmp35726);
  assign tmp36211 = s2 ? tmp36212 : tmp36214;
  assign tmp36217 = s0 ? tmp36068 : tmp35983;
  assign tmp36216 = s1 ? tmp36217 : tmp35984;
  assign tmp36215 = s2 ? tmp36216 : tmp35985;
  assign tmp36210 = s3 ? tmp36211 : tmp36215;
  assign tmp36199 = s4 ? tmp36200 : tmp36210;
  assign tmp36198 = ~(s5 ? tmp36199 : tmp36071);
  assign tmp36171 = s6 ? tmp36172 : tmp36198;
  assign tmp36170 = s7 ? tmp35709 : tmp36171;
  assign tmp36169 = s8 ? tmp36170 : tmp35709;
  assign tmp36225 = ~(s1 ? tmp35772 : tmp35977);
  assign tmp36224 = s2 ? tmp35969 : tmp36225;
  assign tmp36223 = s3 ? tmp36224 : tmp35978;
  assign tmp36222 = s4 ? tmp35948 : tmp36223;
  assign tmp36221 = ~(s5 ? tmp36222 : tmp35987);
  assign tmp36220 = s6 ? tmp35900 : tmp36221;
  assign tmp36219 = s7 ? tmp36220 : tmp36082;
  assign tmp36226 = s7 ? tmp36011 : tmp36171;
  assign tmp36218 = s8 ? tmp36219 : tmp36226;
  assign tmp36168 = s9 ? tmp36169 : tmp36218;
  assign tmp35705 = s10 ? tmp35706 : tmp36168;
  assign tmp36230 = s7 ? tmp35899 : tmp36082;
  assign tmp36229 = s8 ? tmp36230 : tmp36226;
  assign tmp36228 = s9 ? tmp36169 : tmp36229;
  assign tmp36227 = s10 ? tmp35706 : tmp36228;
  assign tmp35704 = s11 ? tmp35705 : tmp36227;
  assign tmp36243 = l1 ? tmp35914 : tmp35717;
  assign tmp36244 = ~(l1 ? tmp35916 : tmp35882);
  assign tmp36242 = s0 ? tmp36243 : tmp36244;
  assign tmp36246 = l1 ? tmp35916 : tmp35882;
  assign tmp36245 = ~(s0 ? tmp36088 : tmp36246);
  assign tmp36241 = s1 ? tmp36242 : tmp36245;
  assign tmp36248 = s0 ? tmp36088 : tmp35749;
  assign tmp36249 = s0 ? tmp36246 : tmp36105;
  assign tmp36247 = ~(s1 ? tmp36248 : tmp36249);
  assign tmp36240 = s2 ? tmp36241 : tmp36247;
  assign tmp36239 = s3 ? tmp36085 : tmp36240;
  assign tmp36253 = ~(s0 ? tmp36086 : tmp36244);
  assign tmp36252 = s1 ? tmp36109 : tmp36253;
  assign tmp36255 = s0 ? tmp36086 : tmp35761;
  assign tmp36256 = s0 ? tmp36116 : tmp35766;
  assign tmp36254 = ~(s1 ? tmp36255 : tmp36256);
  assign tmp36251 = s2 ? tmp36252 : tmp36254;
  assign tmp36259 = s0 ? tmp35775 : tmp35938;
  assign tmp36258 = s1 ? tmp36088 : tmp36259;
  assign tmp36263 = ~(l2 ? tmp35778 : tmp35716);
  assign tmp36262 = ~(l1 ? tmp35926 : tmp36263);
  assign tmp36261 = s0 ? tmp36246 : tmp36262;
  assign tmp36264 = s0 ? tmp35944 : tmp36246;
  assign tmp36260 = s1 ? tmp36261 : tmp36264;
  assign tmp36257 = s2 ? tmp36258 : tmp36260;
  assign tmp36250 = ~(s3 ? tmp36251 : tmp36257);
  assign tmp36238 = s4 ? tmp36239 : tmp36250;
  assign tmp36270 = ~(s0 ? tmp35795 : tmp36243);
  assign tmp36269 = s1 ? tmp36129 : tmp36270;
  assign tmp36272 = s0 ? tmp35795 : tmp36132;
  assign tmp36274 = l1 ? tmp35926 : tmp36263;
  assign tmp36273 = s0 ? tmp36274 : tmp35801;
  assign tmp36271 = ~(s1 ? tmp36272 : tmp36273);
  assign tmp36268 = s2 ? tmp36269 : tmp36271;
  assign tmp36278 = ~(l1 ? 1 : tmp35764);
  assign tmp36277 = s0 ? 1 : tmp36278;
  assign tmp36280 = ~(l1 ? tmp35777 : tmp35882);
  assign tmp36279 = s0 ? 1 : tmp36280;
  assign tmp36276 = s1 ? tmp36277 : tmp36279;
  assign tmp36283 = l1 ? tmp35966 : tmp35882;
  assign tmp36282 = s0 ? tmp36246 : tmp36283;
  assign tmp36281 = ~(s1 ? tmp35963 : tmp36282);
  assign tmp36275 = ~(s2 ? tmp36276 : tmp36281);
  assign tmp36267 = s3 ? tmp36268 : tmp36275;
  assign tmp36288 = l2 ? tmp35765 : tmp35724;
  assign tmp36287 = ~(l1 ? tmp35926 : tmp36288);
  assign tmp36286 = s1 ? tmp36151 : tmp36287;
  assign tmp36285 = s2 ? tmp36286 : tmp35985;
  assign tmp36284 = s3 ? tmp36143 : tmp36285;
  assign tmp36266 = s4 ? tmp36267 : tmp36284;
  assign tmp36293 = s0 ? tmp35938 : tmp35850;
  assign tmp36292 = s1 ? tmp36293 : tmp35992;
  assign tmp36294 = s1 ? 1 : tmp35888;
  assign tmp36291 = s2 ? tmp36292 : tmp36294;
  assign tmp36290 = s3 ? tmp36291 : tmp36160;
  assign tmp36289 = s4 ? tmp36290 : tmp36163;
  assign tmp36265 = ~(s5 ? tmp36266 : tmp36289);
  assign tmp36237 = s6 ? tmp36238 : tmp36265;
  assign tmp36236 = s7 ? tmp35709 : tmp36237;
  assign tmp36300 = l1 ? tmp35926 : tmp35773;
  assign tmp36302 = l1 ? tmp36017 : tmp36090;
  assign tmp36301 = ~(s0 ? tmp35906 : tmp36302);
  assign tmp36299 = s1 ? tmp36300 : tmp36301;
  assign tmp36306 = l1 ? tmp35865 : tmp36096;
  assign tmp36307 = ~(l1 ? tmp35916 : tmp35945);
  assign tmp36305 = s0 ? tmp36306 : tmp36307;
  assign tmp36309 = l1 ? tmp35916 : tmp35945;
  assign tmp36308 = ~(s0 ? tmp35906 : tmp36309);
  assign tmp36304 = s1 ? tmp36305 : tmp36308;
  assign tmp36311 = s0 ? tmp35906 : tmp36027;
  assign tmp36313 = ~(l1 ? tmp35926 : tmp35773);
  assign tmp36312 = s0 ? tmp36309 : tmp36313;
  assign tmp36310 = ~(s1 ? tmp36311 : tmp36312);
  assign tmp36303 = s2 ? tmp36304 : tmp36310;
  assign tmp36298 = s3 ? tmp36299 : tmp36303;
  assign tmp36318 = l1 ? tmp35723 : tmp36090;
  assign tmp36317 = s0 ? tmp36318 : tmp35757;
  assign tmp36319 = ~(s0 ? tmp36300 : tmp36307);
  assign tmp36316 = s1 ? tmp36317 : tmp36319;
  assign tmp36321 = s0 ? tmp36300 : tmp35761;
  assign tmp36320 = ~(s1 ? tmp36321 : tmp35823);
  assign tmp36315 = s2 ? tmp36316 : tmp36320;
  assign tmp36325 = ~(l1 ? tmp35926 : tmp36122);
  assign tmp36324 = s0 ? tmp36309 : tmp36325;
  assign tmp36326 = s0 ? tmp35944 : tmp36309;
  assign tmp36323 = s1 ? tmp36324 : tmp36326;
  assign tmp36322 = s2 ? tmp35937 : tmp36323;
  assign tmp36314 = ~(s3 ? tmp36315 : tmp36322);
  assign tmp36297 = s4 ? tmp36298 : tmp36314;
  assign tmp36332 = s0 ? tmp36302 : tmp35793;
  assign tmp36333 = ~(s0 ? tmp35795 : tmp36306);
  assign tmp36331 = s1 ? tmp36332 : tmp36333;
  assign tmp36335 = s0 ? tmp35795 : tmp36165;
  assign tmp36337 = l1 ? tmp35926 : tmp36122;
  assign tmp36336 = s0 ? tmp36337 : tmp36054;
  assign tmp36334 = ~(s1 ? tmp36335 : tmp36336);
  assign tmp36330 = s2 ? tmp36331 : tmp36334;
  assign tmp36340 = l1 ? tmp35767 : tmp35764;
  assign tmp36339 = s1 ? tmp36340 : tmp35944;
  assign tmp36343 = l1 ? tmp35966 : tmp35945;
  assign tmp36342 = s0 ? tmp36309 : tmp36343;
  assign tmp36341 = s1 ? tmp35963 : tmp36342;
  assign tmp36338 = s2 ? tmp36339 : tmp36341;
  assign tmp36329 = s3 ? tmp36330 : tmp36338;
  assign tmp36347 = s0 ? tmp35971 : tmp36309;
  assign tmp36346 = s1 ? tmp36347 : tmp35974;
  assign tmp36348 = ~(l1 ? tmp35865 : tmp35744);
  assign tmp36345 = s2 ? tmp36346 : tmp36348;
  assign tmp36352 = l1 ? tmp36070 : tmp35945;
  assign tmp36351 = s0 ? tmp36152 : tmp36352;
  assign tmp36350 = s1 ? tmp36351 : tmp36287;
  assign tmp36349 = s2 ? tmp36350 : tmp35985;
  assign tmp36344 = s3 ? tmp36345 : tmp36349;
  assign tmp36328 = s4 ? tmp36329 : tmp36344;
  assign tmp36356 = s1 ? tmp35887 : tmp35888;
  assign tmp36355 = s2 ? tmp36158 : tmp36356;
  assign tmp36354 = s3 ? tmp36355 : tmp36160;
  assign tmp36353 = s4 ? tmp36354 : tmp36163;
  assign tmp36327 = ~(s5 ? tmp36328 : tmp36353);
  assign tmp36296 = s6 ? tmp36297 : tmp36327;
  assign tmp36295 = s7 ? tmp35709 : tmp36296;
  assign tmp36235 = s8 ? tmp36236 : tmp36295;
  assign tmp36362 = s1 ? tmp35903 : tmp36087;
  assign tmp36361 = s3 ? tmp36362 : tmp36176;
  assign tmp36365 = s1 ? tmp36109 : tmp36190;
  assign tmp36364 = s2 ? tmp36365 : tmp36191;
  assign tmp36363 = ~(s3 ? tmp36364 : tmp36193);
  assign tmp36360 = s4 ? tmp36361 : tmp36363;
  assign tmp36371 = ~(s0 ? tmp35795 : tmp36179);
  assign tmp36370 = s1 ? tmp36129 : tmp36371;
  assign tmp36372 = ~(s1 ? tmp36272 : tmp36206);
  assign tmp36369 = s2 ? tmp36370 : tmp36372;
  assign tmp36374 = s1 ? tmp35960 : tmp35944;
  assign tmp36376 = s0 ? tmp36100 : tmp35944;
  assign tmp36375 = s1 ? tmp35963 : tmp36376;
  assign tmp36373 = s2 ? tmp36374 : tmp36375;
  assign tmp36368 = s3 ? tmp36369 : tmp36373;
  assign tmp36367 = s4 ? tmp36368 : tmp36284;
  assign tmp36366 = ~(s5 ? tmp36367 : tmp36353);
  assign tmp36359 = s6 ? tmp36360 : tmp36366;
  assign tmp36358 = s7 ? tmp35709 : tmp36359;
  assign tmp36357 = s8 ? tmp36295 : tmp36358;
  assign tmp36234 = s9 ? tmp36235 : tmp36357;
  assign tmp36386 = ~(s0 ? tmp35795 : tmp36095);
  assign tmp36385 = s1 ? tmp36129 : tmp36386;
  assign tmp36387 = ~(s1 ? tmp36272 : tmp36133);
  assign tmp36384 = s2 ? tmp36385 : tmp36387;
  assign tmp36388 = s2 ? tmp36137 : tmp36375;
  assign tmp36383 = s3 ? tmp36384 : tmp36388;
  assign tmp36382 = s4 ? tmp36383 : tmp36284;
  assign tmp36381 = ~(s5 ? tmp36382 : tmp36353);
  assign tmp36380 = s6 ? tmp36083 : tmp36381;
  assign tmp36379 = s7 ? tmp35709 : tmp36380;
  assign tmp36378 = s8 ? tmp36379 : tmp35709;
  assign tmp36394 = s2 ? tmp36118 : tmp36260;
  assign tmp36393 = ~(s3 ? tmp36251 : tmp36394);
  assign tmp36392 = s4 ? tmp36239 : tmp36393;
  assign tmp36399 = ~(s1 ? tmp36132 : tmp36273);
  assign tmp36398 = s2 ? tmp36269 : tmp36399;
  assign tmp36401 = s1 ? tmp36277 : tmp36280;
  assign tmp36400 = ~(s2 ? tmp36401 : tmp36281);
  assign tmp36397 = s3 ? tmp36398 : tmp36400;
  assign tmp36396 = s4 ? tmp36397 : tmp36284;
  assign tmp36395 = ~(s5 ? tmp36396 : tmp36289);
  assign tmp36391 = s6 ? tmp36392 : tmp36395;
  assign tmp36407 = ~(s1 ? tmp36132 : tmp36206);
  assign tmp36406 = s2 ? tmp36370 : tmp36407;
  assign tmp36405 = s3 ? tmp36406 : tmp36373;
  assign tmp36404 = s4 ? tmp36405 : tmp36284;
  assign tmp36403 = ~(s5 ? tmp36404 : tmp36353);
  assign tmp36402 = s6 ? tmp36360 : tmp36403;
  assign tmp36390 = s7 ? tmp36391 : tmp36402;
  assign tmp36414 = ~(s1 ? tmp36165 : tmp36336);
  assign tmp36413 = s2 ? tmp36331 : tmp36414;
  assign tmp36412 = s3 ? tmp36413 : tmp36338;
  assign tmp36411 = s4 ? tmp36412 : tmp36344;
  assign tmp36410 = ~(s5 ? tmp36411 : tmp36353);
  assign tmp36409 = s6 ? tmp36297 : tmp36410;
  assign tmp36419 = s2 ? tmp36385 : tmp36131;
  assign tmp36418 = s3 ? tmp36419 : tmp36388;
  assign tmp36417 = s4 ? tmp36418 : tmp36284;
  assign tmp36416 = ~(s5 ? tmp36417 : tmp36353);
  assign tmp36415 = s6 ? tmp36083 : tmp36416;
  assign tmp36408 = s7 ? tmp36409 : tmp36415;
  assign tmp36389 = s8 ? tmp36390 : tmp36408;
  assign tmp36377 = s9 ? tmp36378 : tmp36389;
  assign tmp36233 = s10 ? tmp36234 : tmp36377;
  assign tmp36423 = s7 ? tmp36237 : tmp36359;
  assign tmp36424 = s7 ? tmp36296 : tmp36380;
  assign tmp36422 = s8 ? tmp36423 : tmp36424;
  assign tmp36421 = s9 ? tmp36378 : tmp36422;
  assign tmp36420 = s10 ? tmp36234 : tmp36421;
  assign tmp36232 = s11 ? tmp36233 : tmp36420;
  assign tmp36434 = l1 ? tmp35904 : tmp36096;
  assign tmp36436 = l1 ? tmp35768 : tmp35806;
  assign tmp36437 = l1 ? tmp35908 : tmp36153;
  assign tmp36435 = ~(s0 ? tmp36436 : tmp36437);
  assign tmp36433 = s1 ? tmp36434 : tmp36435;
  assign tmp36441 = l1 ? tmp35914 : tmp35773;
  assign tmp36443 = ~(l2 ? tmp35765 : tmp35717);
  assign tmp36442 = ~(l1 ? tmp36098 : tmp36443);
  assign tmp36440 = s0 ? tmp36441 : tmp36442;
  assign tmp36445 = l1 ? tmp36098 : tmp36443;
  assign tmp36444 = ~(s0 ? tmp36436 : tmp36445);
  assign tmp36439 = s1 ? tmp36440 : tmp36444;
  assign tmp36448 = l1 ? tmp35723 : tmp35955;
  assign tmp36447 = s0 ? tmp36436 : tmp36448;
  assign tmp36450 = ~(l1 ? tmp35904 : tmp36096);
  assign tmp36449 = s0 ? tmp36445 : tmp36450;
  assign tmp36446 = ~(s1 ? tmp36447 : tmp36449);
  assign tmp36438 = s2 ? tmp36439 : tmp36446;
  assign tmp36432 = s3 ? tmp36433 : tmp36438;
  assign tmp36455 = l1 ? tmp35768 : tmp36153;
  assign tmp36456 = ~(l1 ? tmp35724 : tmp35768);
  assign tmp36454 = s0 ? tmp36455 : tmp36456;
  assign tmp36457 = ~(s0 ? tmp36434 : tmp36442);
  assign tmp36453 = s1 ? tmp36454 : tmp36457;
  assign tmp36459 = s0 ? tmp36434 : tmp35761;
  assign tmp36460 = s0 ? tmp36147 : tmp35766;
  assign tmp36458 = ~(s1 ? tmp36459 : tmp36460);
  assign tmp36452 = s2 ? tmp36453 : tmp36458;
  assign tmp36462 = s1 ? tmp36436 : tmp36259;
  assign tmp36466 = l2 ? tmp35765 : tmp35717;
  assign tmp36465 = ~(l1 ? tmp35904 : tmp36466);
  assign tmp36464 = s0 ? tmp36445 : tmp36465;
  assign tmp36467 = s0 ? tmp35944 : tmp36445;
  assign tmp36463 = s1 ? tmp36464 : tmp36467;
  assign tmp36461 = s2 ? tmp36462 : tmp36463;
  assign tmp36451 = ~(s3 ? tmp36452 : tmp36461);
  assign tmp36431 = s4 ? tmp36432 : tmp36451;
  assign tmp36474 = ~(l1 ? 1 : tmp35768);
  assign tmp36473 = s0 ? tmp36437 : tmp36474;
  assign tmp36475 = ~(l1 ? tmp35914 : tmp35773);
  assign tmp36472 = s1 ? tmp36473 : tmp36475;
  assign tmp36477 = l1 ? tmp35904 : tmp35736;
  assign tmp36479 = l1 ? tmp35904 : tmp36466;
  assign tmp36478 = s0 ? tmp36479 : tmp35775;
  assign tmp36476 = ~(s1 ? tmp36477 : tmp36478);
  assign tmp36471 = s2 ? tmp36472 : tmp36476;
  assign tmp36482 = l1 ? 1 : tmp35806;
  assign tmp36483 = l1 ? tmp35777 : tmp36443;
  assign tmp36481 = s1 ? tmp36482 : tmp36483;
  assign tmp36485 = s0 ? tmp36445 : tmp35944;
  assign tmp36484 = s1 ? tmp35963 : tmp36485;
  assign tmp36480 = s2 ? tmp36481 : tmp36484;
  assign tmp36470 = s3 ? tmp36471 : tmp36480;
  assign tmp36489 = s0 ? tmp35971 : tmp36445;
  assign tmp36490 = ~(l1 ? tmp35724 : 1);
  assign tmp36488 = s1 ? tmp36489 : tmp36490;
  assign tmp36491 = ~(l1 ? tmp35914 : tmp35736);
  assign tmp36487 = s2 ? tmp36488 : tmp36491;
  assign tmp36495 = l1 ? 1 : tmp36090;
  assign tmp36494 = s0 ? tmp36495 : tmp36154;
  assign tmp36493 = s1 ? tmp36494 : tmp36287;
  assign tmp36492 = s2 ? tmp36493 : tmp35985;
  assign tmp36486 = s3 ? tmp36487 : tmp36492;
  assign tmp36469 = s4 ? tmp36470 : tmp36486;
  assign tmp36500 = s0 ? tmp36483 : tmp35850;
  assign tmp36499 = s1 ? tmp36500 : tmp35992;
  assign tmp36502 = l1 ? 1 : tmp35955;
  assign tmp36501 = s1 ? tmp36502 : tmp35888;
  assign tmp36498 = s2 ? tmp36499 : tmp36501;
  assign tmp36497 = s3 ? tmp36498 : tmp36160;
  assign tmp36504 = s2 ? tmp36004 : tmp36167;
  assign tmp36503 = ~(s3 ? tmp36504 : tmp36166);
  assign tmp36496 = s4 ? tmp36497 : tmp36503;
  assign tmp36468 = ~(s5 ? tmp36469 : tmp36496);
  assign tmp36430 = s6 ? tmp36431 : tmp36468;
  assign tmp36429 = s7 ? tmp35709 : tmp36430;
  assign tmp36510 = l1 ? tmp35926 : tmp36096;
  assign tmp36512 = l1 ? tmp35723 : tmp35806;
  assign tmp36513 = l1 ? tmp36017 : tmp36153;
  assign tmp36511 = ~(s0 ? tmp36512 : tmp36513);
  assign tmp36509 = s1 ? tmp36510 : tmp36511;
  assign tmp36517 = l1 ? tmp35865 : tmp35773;
  assign tmp36518 = ~(l1 ? tmp35916 : tmp36443);
  assign tmp36516 = s0 ? tmp36517 : tmp36518;
  assign tmp36520 = l1 ? tmp35916 : tmp36443;
  assign tmp36519 = ~(s0 ? tmp36512 : tmp36520);
  assign tmp36515 = s1 ? tmp36516 : tmp36519;
  assign tmp36522 = s0 ? tmp36512 : tmp36448;
  assign tmp36524 = ~(l1 ? tmp35926 : tmp36096);
  assign tmp36523 = s0 ? tmp36520 : tmp36524;
  assign tmp36521 = ~(s1 ? tmp36522 : tmp36523);
  assign tmp36514 = s2 ? tmp36515 : tmp36521;
  assign tmp36508 = s3 ? tmp36509 : tmp36514;
  assign tmp36529 = l1 ? tmp35723 : tmp36153;
  assign tmp36530 = ~(l1 ? tmp35736 : tmp35768);
  assign tmp36528 = s0 ? tmp36529 : tmp36530;
  assign tmp36531 = ~(s0 ? tmp36510 : tmp36518);
  assign tmp36527 = s1 ? tmp36528 : tmp36531;
  assign tmp36533 = s0 ? tmp36510 : tmp35761;
  assign tmp36532 = ~(s1 ? tmp36533 : tmp35827);
  assign tmp36526 = s2 ? tmp36527 : tmp36532;
  assign tmp36535 = s1 ? tmp36512 : tmp35938;
  assign tmp36538 = ~(l1 ? tmp35926 : tmp36466);
  assign tmp36537 = s0 ? tmp36520 : tmp36538;
  assign tmp36539 = s0 ? tmp35944 : tmp36520;
  assign tmp36536 = s1 ? tmp36537 : tmp36539;
  assign tmp36534 = s2 ? tmp36535 : tmp36536;
  assign tmp36525 = ~(s3 ? tmp36526 : tmp36534);
  assign tmp36507 = s4 ? tmp36508 : tmp36525;
  assign tmp36545 = s0 ? tmp36513 : tmp36474;
  assign tmp36546 = ~(l1 ? tmp35865 : tmp35773);
  assign tmp36544 = s1 ? tmp36545 : tmp36546;
  assign tmp36549 = l1 ? tmp35926 : tmp36466;
  assign tmp36550 = l1 ? 1 : tmp35768;
  assign tmp36548 = s0 ? tmp36549 : tmp36550;
  assign tmp36547 = ~(s1 ? tmp36167 : tmp36548);
  assign tmp36543 = s2 ? tmp36544 : tmp36547;
  assign tmp36553 = l1 ? tmp35767 : tmp35806;
  assign tmp36552 = s1 ? tmp36553 : tmp36483;
  assign tmp36555 = s0 ? tmp36520 : tmp36343;
  assign tmp36554 = s1 ? tmp35963 : tmp36555;
  assign tmp36551 = s2 ? tmp36552 : tmp36554;
  assign tmp36542 = s3 ? tmp36543 : tmp36551;
  assign tmp36559 = s0 ? tmp35971 : tmp36520;
  assign tmp36560 = ~(l1 ? tmp35736 : 1);
  assign tmp36558 = s1 ? tmp36559 : tmp36560;
  assign tmp36557 = s2 ? tmp36558 : tmp35888;
  assign tmp36563 = s0 ? tmp36495 : tmp36352;
  assign tmp36562 = s1 ? tmp36563 : tmp36287;
  assign tmp36561 = s2 ? tmp36562 : tmp35985;
  assign tmp36556 = s3 ? tmp36557 : tmp36561;
  assign tmp36541 = s4 ? tmp36542 : tmp36556;
  assign tmp36540 = ~(s5 ? tmp36541 : tmp36496);
  assign tmp36506 = s6 ? tmp36507 : tmp36540;
  assign tmp36505 = s7 ? tmp35709 : tmp36506;
  assign tmp36428 = s8 ? tmp36429 : tmp36505;
  assign tmp36570 = l1 ? tmp35904 : tmp35725;
  assign tmp36569 = s1 ? tmp36570 : tmp36435;
  assign tmp36574 = l1 ? tmp35914 : tmp35768;
  assign tmp36576 = ~(l2 ? tmp35765 : tmp35725);
  assign tmp36575 = ~(l1 ? tmp36098 : tmp36576);
  assign tmp36573 = s0 ? tmp36574 : tmp36575;
  assign tmp36578 = l1 ? tmp35768 : tmp35914;
  assign tmp36579 = l1 ? tmp36098 : tmp36576;
  assign tmp36577 = ~(s0 ? tmp36578 : tmp36579);
  assign tmp36572 = s1 ? tmp36573 : tmp36577;
  assign tmp36582 = l1 ? tmp35768 : tmp35955;
  assign tmp36581 = s0 ? tmp36578 : tmp36582;
  assign tmp36584 = ~(l1 ? tmp35904 : tmp35725);
  assign tmp36583 = s0 ? tmp36579 : tmp36584;
  assign tmp36580 = ~(s1 ? tmp36581 : tmp36583);
  assign tmp36571 = s2 ? tmp36572 : tmp36580;
  assign tmp36568 = s3 ? tmp36569 : tmp36571;
  assign tmp36588 = ~(s0 ? tmp36570 : tmp36575);
  assign tmp36587 = s1 ? tmp36454 : tmp36588;
  assign tmp36590 = s0 ? tmp36570 : tmp36115;
  assign tmp36589 = ~(s1 ? tmp36590 : tmp36147);
  assign tmp36586 = s2 ? tmp36587 : tmp36589;
  assign tmp36592 = s1 ? tmp36436 : tmp35938;
  assign tmp36596 = l2 ? tmp35765 : tmp35725;
  assign tmp36595 = ~(l1 ? tmp35904 : tmp36596);
  assign tmp36594 = s0 ? tmp36579 : tmp36595;
  assign tmp36597 = s0 ? tmp35944 : tmp36579;
  assign tmp36593 = s1 ? tmp36594 : tmp36597;
  assign tmp36591 = s2 ? tmp36592 : tmp36593;
  assign tmp36585 = ~(s3 ? tmp36586 : tmp36591);
  assign tmp36567 = s4 ? tmp36568 : tmp36585;
  assign tmp36603 = ~(l1 ? tmp35914 : tmp35768);
  assign tmp36602 = s1 ? tmp36473 : tmp36603;
  assign tmp36606 = l1 ? tmp35904 : tmp36596;
  assign tmp36605 = s0 ? tmp36606 : tmp35775;
  assign tmp36604 = ~(s1 ? tmp36477 : tmp36605);
  assign tmp36601 = s2 ? tmp36602 : tmp36604;
  assign tmp36609 = l1 ? 1 : tmp35914;
  assign tmp36608 = s1 ? tmp36609 : tmp36483;
  assign tmp36607 = s2 ? tmp36608 : tmp36484;
  assign tmp36600 = s3 ? tmp36601 : tmp36607;
  assign tmp36599 = s4 ? tmp36600 : tmp36486;
  assign tmp36598 = ~(s5 ? tmp36599 : tmp36496);
  assign tmp36566 = s6 ? tmp36567 : tmp36598;
  assign tmp36565 = s7 ? tmp35709 : tmp36566;
  assign tmp36564 = s8 ? tmp36505 : tmp36565;
  assign tmp36427 = s9 ? tmp36428 : tmp36564;
  assign tmp36618 = s0 ? tmp36436 : tmp36582;
  assign tmp36617 = ~(s1 ? tmp36618 : tmp36449);
  assign tmp36616 = s2 ? tmp36439 : tmp36617;
  assign tmp36615 = s3 ? tmp36433 : tmp36616;
  assign tmp36622 = s0 ? tmp36434 : tmp36115;
  assign tmp36621 = ~(s1 ? tmp36622 : tmp36147);
  assign tmp36620 = s2 ? tmp36453 : tmp36621;
  assign tmp36623 = s2 ? tmp36592 : tmp36463;
  assign tmp36619 = ~(s3 ? tmp36620 : tmp36623);
  assign tmp36614 = s4 ? tmp36615 : tmp36619;
  assign tmp36613 = s6 ? tmp36614 : tmp36468;
  assign tmp36612 = s7 ? tmp35709 : tmp36613;
  assign tmp36611 = s8 ? tmp36612 : tmp35709;
  assign tmp36628 = ~(s3 ? tmp36452 : tmp36623);
  assign tmp36627 = s4 ? tmp36432 : tmp36628;
  assign tmp36626 = s6 ? tmp36627 : tmp36468;
  assign tmp36625 = s7 ? tmp36626 : tmp36566;
  assign tmp36629 = s7 ? tmp36506 : tmp36613;
  assign tmp36624 = s8 ? tmp36625 : tmp36629;
  assign tmp36610 = s9 ? tmp36611 : tmp36624;
  assign tmp36426 = s10 ? tmp36427 : tmp36610;
  assign tmp36633 = s7 ? tmp36430 : tmp36566;
  assign tmp36632 = s8 ? tmp36633 : tmp36629;
  assign tmp36631 = s9 ? tmp36611 : tmp36632;
  assign tmp36630 = s10 ? tmp36427 : tmp36631;
  assign tmp36425 = s11 ? tmp36426 : tmp36630;
  assign tmp36231 = s12 ? tmp36232 : tmp36425;
  assign tmp35703 = s13 ? tmp35704 : tmp36231;
  assign tmp36647 = ~(l1 ? tmp36098 : tmp35882);
  assign tmp36646 = s0 ? tmp36243 : tmp36647;
  assign tmp36649 = l1 ? tmp36098 : tmp35882;
  assign tmp36648 = ~(s0 ? tmp36088 : tmp36649);
  assign tmp36645 = s1 ? tmp36646 : tmp36648;
  assign tmp36652 = l1 ? tmp35768 : 1;
  assign tmp36651 = s0 ? tmp36088 : tmp36652;
  assign tmp36653 = s0 ? tmp36649 : tmp36105;
  assign tmp36650 = ~(s1 ? tmp36651 : tmp36653);
  assign tmp36644 = s2 ? tmp36645 : tmp36650;
  assign tmp36643 = s3 ? tmp36085 : tmp36644;
  assign tmp36657 = ~(s0 ? tmp36086 : tmp36647);
  assign tmp36656 = s1 ? tmp36109 : tmp36657;
  assign tmp36655 = s2 ? tmp36656 : tmp36113;
  assign tmp36660 = s0 ? tmp36649 : tmp36262;
  assign tmp36661 = s0 ? tmp35944 : tmp36649;
  assign tmp36659 = s1 ? tmp36660 : tmp36661;
  assign tmp36658 = s2 ? tmp36118 : tmp36659;
  assign tmp36654 = ~(s3 ? tmp36655 : tmp36658);
  assign tmp36642 = s4 ? tmp36643 : tmp36654;
  assign tmp36667 = ~(l1 ? tmp35914 : tmp35717);
  assign tmp36666 = s1 ? tmp36129 : tmp36667;
  assign tmp36665 = s2 ? tmp36666 : tmp36399;
  assign tmp36670 = s0 ? tmp36649 : tmp35944;
  assign tmp36669 = ~(s1 ? tmp35963 : tmp36670);
  assign tmp36668 = ~(s2 ? tmp36276 : tmp36669);
  assign tmp36664 = s3 ? tmp36665 : tmp36668;
  assign tmp36663 = s4 ? tmp36664 : tmp36284;
  assign tmp36662 = ~(s5 ? tmp36663 : tmp36289);
  assign tmp36641 = s6 ? tmp36642 : tmp36662;
  assign tmp36640 = s7 ? tmp35709 : tmp36641;
  assign tmp36677 = l2 ? tmp35724 : tmp35717;
  assign tmp36676 = l1 ? tmp35904 : tmp36677;
  assign tmp36680 = ~(l2 ? tmp35715 : 0);
  assign tmp36679 = l1 ? tmp35768 : tmp36680;
  assign tmp36682 = ~(l2 ? tmp35715 : tmp36091);
  assign tmp36681 = l1 ? tmp35908 : tmp36682;
  assign tmp36678 = ~(s0 ? tmp36679 : tmp36681);
  assign tmp36675 = s1 ? tmp36676 : tmp36678;
  assign tmp36685 = ~(s0 ? tmp36679 : tmp36649);
  assign tmp36684 = s1 ? tmp36646 : tmp36685;
  assign tmp36687 = s0 ? tmp36679 : tmp36652;
  assign tmp36689 = ~(l1 ? tmp35904 : tmp36677);
  assign tmp36688 = s0 ? tmp36649 : tmp36689;
  assign tmp36686 = ~(s1 ? tmp36687 : tmp36688);
  assign tmp36683 = s2 ? tmp36684 : tmp36686;
  assign tmp36674 = s3 ? tmp36675 : tmp36683;
  assign tmp36694 = l1 ? tmp35768 : tmp36682;
  assign tmp36693 = s0 ? tmp36694 : tmp36111;
  assign tmp36695 = ~(s0 ? tmp36676 : tmp36647);
  assign tmp36692 = s1 ? tmp36693 : tmp36695;
  assign tmp36697 = s0 ? tmp36676 : tmp36115;
  assign tmp36698 = l1 ? tmp35724 : tmp35955;
  assign tmp36696 = ~(s1 ? tmp36697 : tmp36698);
  assign tmp36691 = s2 ? tmp36692 : tmp36696;
  assign tmp36700 = s1 ? tmp36679 : tmp35938;
  assign tmp36703 = ~(l1 ? tmp35904 : tmp36263);
  assign tmp36702 = s0 ? tmp36649 : tmp36703;
  assign tmp36704 = s0 ? tmp35938 : tmp36649;
  assign tmp36701 = s1 ? tmp36702 : tmp36704;
  assign tmp36699 = s2 ? tmp36700 : tmp36701;
  assign tmp36690 = ~(s3 ? tmp36691 : tmp36699);
  assign tmp36673 = s4 ? tmp36674 : tmp36690;
  assign tmp36710 = s0 ? tmp36681 : tmp35793;
  assign tmp36709 = s1 ? tmp36710 : tmp36667;
  assign tmp36713 = ~(l2 ? tmp35716 : tmp35745);
  assign tmp36712 = l1 ? tmp35904 : tmp36713;
  assign tmp36715 = l1 ? tmp35904 : tmp36263;
  assign tmp36716 = l1 ? tmp35767 : tmp35737;
  assign tmp36714 = s0 ? tmp36715 : tmp36716;
  assign tmp36711 = ~(s1 ? tmp36712 : tmp36714);
  assign tmp36708 = s2 ? tmp36709 : tmp36711;
  assign tmp36719 = l1 ? 1 : tmp36680;
  assign tmp36718 = s1 ? tmp36719 : tmp35938;
  assign tmp36721 = s0 ? tmp36649 : tmp35938;
  assign tmp36720 = s1 ? tmp36293 : tmp36721;
  assign tmp36717 = s2 ? tmp36718 : tmp36720;
  assign tmp36707 = s3 ? tmp36708 : tmp36717;
  assign tmp36725 = s0 ? tmp35971 : tmp36649;
  assign tmp36727 = l1 ? tmp35724 : tmp35767;
  assign tmp36726 = ~(s0 ? tmp36116 : tmp36727);
  assign tmp36724 = s1 ? tmp36725 : tmp36726;
  assign tmp36728 = ~(l1 ? tmp35914 : tmp36713);
  assign tmp36723 = s2 ? tmp36724 : tmp36728;
  assign tmp36732 = l1 ? 1 : tmp35778;
  assign tmp36731 = s0 ? tmp36732 : tmp35971;
  assign tmp36730 = s1 ? tmp36731 : tmp36287;
  assign tmp36729 = s2 ? tmp36730 : tmp35985;
  assign tmp36722 = s3 ? tmp36723 : tmp36729;
  assign tmp36706 = s4 ? tmp36707 : tmp36722;
  assign tmp36737 = ~(l1 ? tmp35857 : tmp35767);
  assign tmp36736 = s1 ? tmp36293 : tmp36737;
  assign tmp36735 = s2 ? tmp36736 : tmp36294;
  assign tmp36734 = s3 ? tmp36735 : tmp36160;
  assign tmp36740 = s1 ? tmp35856 : tmp36280;
  assign tmp36741 = l1 ? tmp35926 : tmp36713;
  assign tmp36739 = s2 ? tmp36740 : tmp36741;
  assign tmp36738 = ~(s3 ? tmp36739 : tmp36166);
  assign tmp36733 = s4 ? tmp36734 : tmp36738;
  assign tmp36705 = ~(s5 ? tmp36706 : tmp36733);
  assign tmp36672 = s6 ? tmp36673 : tmp36705;
  assign tmp36671 = s7 ? tmp35709 : tmp36672;
  assign tmp36639 = s8 ? tmp36640 : tmp36671;
  assign tmp36748 = l1 ? tmp35904 : tmp35723;
  assign tmp36751 = ~(l2 ? tmp35715 : tmp35720);
  assign tmp36750 = l1 ? tmp35908 : tmp36751;
  assign tmp36749 = ~(s0 ? tmp36679 : tmp36750);
  assign tmp36747 = s1 ? tmp36748 : tmp36749;
  assign tmp36755 = ~(l1 ? tmp36098 : tmp35917);
  assign tmp36754 = s0 ? tmp35913 : tmp36755;
  assign tmp36758 = ~(l2 ? tmp35715 : tmp35745);
  assign tmp36757 = l1 ? tmp35768 : tmp36758;
  assign tmp36759 = l1 ? tmp36098 : tmp35917;
  assign tmp36756 = ~(s0 ? tmp36757 : tmp36759);
  assign tmp36753 = s1 ? tmp36754 : tmp36756;
  assign tmp36761 = s0 ? tmp36757 : tmp36652;
  assign tmp36763 = ~(l1 ? tmp35904 : tmp35723);
  assign tmp36762 = s0 ? tmp36759 : tmp36763;
  assign tmp36760 = ~(s1 ? tmp36761 : tmp36762);
  assign tmp36752 = s2 ? tmp36753 : tmp36760;
  assign tmp36746 = s3 ? tmp36747 : tmp36752;
  assign tmp36768 = l1 ? tmp35768 : tmp36751;
  assign tmp36767 = s0 ? tmp36768 : tmp36111;
  assign tmp36769 = ~(s0 ? tmp36748 : tmp36755);
  assign tmp36766 = s1 ? tmp36767 : tmp36769;
  assign tmp36771 = s0 ? tmp36748 : tmp36115;
  assign tmp36770 = ~(s1 ? tmp36771 : tmp36698);
  assign tmp36765 = s2 ? tmp36766 : tmp36770;
  assign tmp36775 = ~(l1 ? tmp35904 : tmp35942);
  assign tmp36774 = s0 ? tmp36759 : tmp36775;
  assign tmp36776 = s0 ? tmp35938 : tmp36759;
  assign tmp36773 = s1 ? tmp36774 : tmp36776;
  assign tmp36772 = s2 ? tmp36700 : tmp36773;
  assign tmp36764 = ~(s3 ? tmp36765 : tmp36772);
  assign tmp36745 = s4 ? tmp36746 : tmp36764;
  assign tmp36782 = s0 ? tmp36750 : tmp35793;
  assign tmp36781 = s1 ? tmp36782 : tmp35952;
  assign tmp36785 = l1 ? tmp35904 : tmp35942;
  assign tmp36784 = s0 ? tmp36785 : tmp36716;
  assign tmp36783 = ~(s1 ? tmp35954 : tmp36784);
  assign tmp36780 = s2 ? tmp36781 : tmp36783;
  assign tmp36788 = l1 ? 1 : tmp36758;
  assign tmp36787 = s1 ? tmp36788 : tmp35961;
  assign tmp36790 = s0 ? tmp36759 : tmp35961;
  assign tmp36789 = s1 ? tmp36293 : tmp36790;
  assign tmp36786 = s2 ? tmp36787 : tmp36789;
  assign tmp36779 = s3 ? tmp36780 : tmp36786;
  assign tmp36793 = ~(l1 ? tmp35914 : tmp35955);
  assign tmp36792 = s2 ? tmp36724 : tmp36793;
  assign tmp36796 = s0 ? tmp35981 : tmp35971;
  assign tmp36795 = s1 ? tmp36796 : tmp36287;
  assign tmp36794 = s2 ? tmp36795 : tmp35985;
  assign tmp36791 = s3 ? tmp36792 : tmp36794;
  assign tmp36778 = s4 ? tmp36779 : tmp36791;
  assign tmp36800 = s1 ? tmp35991 : tmp36737;
  assign tmp36801 = s1 ? tmp35994 : tmp35888;
  assign tmp36799 = s2 ? tmp36800 : tmp36801;
  assign tmp36798 = s3 ? tmp36799 : tmp36160;
  assign tmp36803 = s2 ? tmp36740 : tmp36006;
  assign tmp36802 = ~(s3 ? tmp36803 : tmp36166);
  assign tmp36797 = s4 ? tmp36798 : tmp36802;
  assign tmp36777 = ~(s5 ? tmp36778 : tmp36797);
  assign tmp36744 = s6 ? tmp36745 : tmp36777;
  assign tmp36743 = s7 ? tmp35709 : tmp36744;
  assign tmp36742 = s8 ? tmp36671 : tmp36743;
  assign tmp36638 = s9 ? tmp36639 : tmp36742;
  assign tmp36805 = s8 ? tmp36671 : tmp35709;
  assign tmp36812 = ~(s2 ? tmp36401 : tmp36669);
  assign tmp36811 = s3 ? tmp36665 : tmp36812;
  assign tmp36810 = s4 ? tmp36811 : tmp36284;
  assign tmp36809 = ~(s5 ? tmp36810 : tmp36289);
  assign tmp36808 = s6 ? tmp36642 : tmp36809;
  assign tmp36807 = s7 ? tmp36808 : tmp36744;
  assign tmp36806 = s8 ? tmp36807 : tmp36672;
  assign tmp36804 = s9 ? tmp36805 : tmp36806;
  assign tmp36637 = s10 ? tmp36638 : tmp36804;
  assign tmp36816 = s7 ? tmp36641 : tmp36744;
  assign tmp36815 = s8 ? tmp36816 : tmp36672;
  assign tmp36814 = s9 ? tmp36805 : tmp36815;
  assign tmp36813 = s10 ? tmp36638 : tmp36814;
  assign tmp36636 = s11 ? tmp36637 : tmp36813;
  assign tmp36827 = ~(l2 ? tmp35765 : tmp35727);
  assign tmp36826 = l1 ? tmp35904 : tmp36827;
  assign tmp36829 = l1 ? tmp35908 : tmp35740;
  assign tmp36828 = ~(s0 ? tmp35749 : tmp36829);
  assign tmp36825 = s1 ? tmp36826 : tmp36828;
  assign tmp36833 = l1 ? tmp35914 : tmp35723;
  assign tmp36835 = ~(l2 ? tmp35727 : tmp35725);
  assign tmp36834 = ~(l1 ? tmp36098 : tmp36835);
  assign tmp36832 = s0 ? tmp36833 : tmp36834;
  assign tmp36837 = l1 ? tmp35768 : tmp35736;
  assign tmp36838 = l1 ? tmp36098 : tmp36835;
  assign tmp36836 = ~(s0 ? tmp36837 : tmp36838);
  assign tmp36831 = s1 ? tmp36832 : tmp36836;
  assign tmp36840 = s0 ? tmp36837 : tmp36582;
  assign tmp36842 = ~(l1 ? tmp35904 : tmp36827);
  assign tmp36841 = s0 ? tmp36838 : tmp36842;
  assign tmp36839 = ~(s1 ? tmp36840 : tmp36841);
  assign tmp36830 = s2 ? tmp36831 : tmp36839;
  assign tmp36824 = s3 ? tmp36825 : tmp36830;
  assign tmp36847 = l1 ? tmp35768 : tmp35740;
  assign tmp36846 = s0 ? tmp36847 : tmp36530;
  assign tmp36848 = ~(s0 ? tmp36826 : tmp36834);
  assign tmp36845 = s1 ? tmp36846 : tmp36848;
  assign tmp36850 = s0 ? tmp36826 : tmp36115;
  assign tmp36849 = ~(s1 ? tmp36850 : tmp35824);
  assign tmp36844 = s2 ? tmp36845 : tmp36849;
  assign tmp36854 = l2 ? 1 : tmp35716;
  assign tmp36853 = l1 ? tmp35777 : tmp36854;
  assign tmp36852 = s1 ? tmp35749 : tmp36853;
  assign tmp36858 = l2 ? tmp35727 : tmp35725;
  assign tmp36857 = ~(l1 ? tmp35926 : tmp36858);
  assign tmp36856 = s0 ? tmp36838 : tmp36857;
  assign tmp36859 = s0 ? tmp36853 : tmp36838;
  assign tmp36855 = s1 ? tmp36856 : tmp36859;
  assign tmp36851 = s2 ? tmp36852 : tmp36855;
  assign tmp36843 = ~(s3 ? tmp36844 : tmp36851);
  assign tmp36823 = s4 ? tmp36824 : tmp36843;
  assign tmp36865 = s0 ? tmp36829 : tmp36474;
  assign tmp36866 = ~(l1 ? tmp35914 : tmp35723);
  assign tmp36864 = s1 ? tmp36865 : tmp36866;
  assign tmp36868 = l1 ? tmp35904 : tmp35806;
  assign tmp36870 = l1 ? tmp35926 : tmp36858;
  assign tmp36869 = s0 ? tmp36870 : tmp35775;
  assign tmp36867 = ~(s1 ? tmp36868 : tmp36869);
  assign tmp36863 = s2 ? tmp36864 : tmp36867;
  assign tmp36873 = l1 ? tmp35777 : tmp36835;
  assign tmp36872 = s1 ? tmp35994 : tmp36873;
  assign tmp36875 = s0 ? tmp36853 : tmp35850;
  assign tmp36878 = l2 ? 1 : tmp35727;
  assign tmp36877 = l1 ? tmp35966 : tmp36878;
  assign tmp36876 = s0 ? tmp36838 : tmp36877;
  assign tmp36874 = s1 ? tmp36875 : tmp36876;
  assign tmp36871 = s2 ? tmp36872 : tmp36874;
  assign tmp36862 = s3 ? tmp36863 : tmp36871;
  assign tmp36883 = l1 ? tmp35821 : tmp36854;
  assign tmp36882 = s0 ? tmp36883 : tmp36838;
  assign tmp36884 = ~(s0 ? tmp35827 : tmp35824);
  assign tmp36881 = s1 ? tmp36882 : tmp36884;
  assign tmp36886 = l1 ? tmp35914 : tmp35806;
  assign tmp36885 = ~(s1 ? tmp35827 : tmp36886);
  assign tmp36880 = s2 ? tmp36881 : tmp36885;
  assign tmp36890 = l1 ? 1 : tmp35731;
  assign tmp36891 = l1 ? tmp35821 : tmp36878;
  assign tmp36889 = s0 ? tmp36890 : tmp36891;
  assign tmp36894 = l2 ? tmp35716 : 1;
  assign tmp36893 = l1 ? tmp35926 : tmp36894;
  assign tmp36892 = ~(s0 ? tmp35827 : tmp36893);
  assign tmp36888 = s1 ? tmp36889 : tmp36892;
  assign tmp36895 = s1 ? tmp35986 : tmp36853;
  assign tmp36887 = s2 ? tmp36888 : tmp36895;
  assign tmp36879 = s3 ? tmp36880 : tmp36887;
  assign tmp36861 = s4 ? tmp36862 : tmp36879;
  assign tmp36900 = s0 ? tmp36873 : tmp35850;
  assign tmp36901 = ~(l1 ? tmp35857 : tmp35806);
  assign tmp36899 = s1 ? tmp36900 : tmp36901;
  assign tmp36903 = l1 ? 1 : tmp36713;
  assign tmp36902 = s1 ? tmp36903 : tmp35995;
  assign tmp36898 = s2 ? tmp36899 : tmp36902;
  assign tmp36906 = l1 ? tmp35812 : tmp35833;
  assign tmp36907 = ~(l1 ? 1 : tmp35740);
  assign tmp36905 = s1 ? tmp36906 : tmp36907;
  assign tmp36904 = ~(s2 ? tmp35997 : tmp36905);
  assign tmp36897 = s3 ? tmp36898 : tmp36904;
  assign tmp36911 = ~(l1 ? tmp35777 : tmp36854);
  assign tmp36910 = s1 ? tmp35856 : tmp36911;
  assign tmp36912 = l1 ? tmp35926 : tmp35806;
  assign tmp36909 = s2 ? tmp36910 : tmp36912;
  assign tmp36914 = l1 ? tmp35926 : tmp35833;
  assign tmp36913 = s1 ? tmp36008 : tmp36914;
  assign tmp36908 = ~(s3 ? tmp36909 : tmp36913);
  assign tmp36896 = s4 ? tmp36897 : tmp36908;
  assign tmp36860 = ~(s5 ? tmp36861 : tmp36896);
  assign tmp36822 = s6 ? tmp36823 : tmp36860;
  assign tmp36821 = s7 ? tmp35709 : tmp36822;
  assign tmp36921 = ~(l2 ? tmp35715 : tmp35727);
  assign tmp36920 = l1 ? tmp35904 : tmp36921;
  assign tmp36924 = l2 ? tmp35724 : tmp35719;
  assign tmp36923 = l1 ? tmp35908 : tmp36924;
  assign tmp36922 = ~(s0 ? tmp36103 : tmp36923);
  assign tmp36919 = s1 ? tmp36920 : tmp36922;
  assign tmp36929 = ~(l2 ? tmp35716 : tmp35725);
  assign tmp36928 = ~(l1 ? tmp36098 : tmp36929);
  assign tmp36927 = s0 ? tmp36574 : tmp36928;
  assign tmp36931 = l1 ? tmp35768 : tmp35724;
  assign tmp36932 = l1 ? tmp36098 : tmp36929;
  assign tmp36930 = ~(s0 ? tmp36931 : tmp36932);
  assign tmp36926 = s1 ? tmp36927 : tmp36930;
  assign tmp36934 = s0 ? tmp36931 : tmp36582;
  assign tmp36936 = ~(l1 ? tmp35904 : tmp36921);
  assign tmp36935 = s0 ? tmp36932 : tmp36936;
  assign tmp36933 = ~(s1 ? tmp36934 : tmp36935);
  assign tmp36925 = s2 ? tmp36926 : tmp36933;
  assign tmp36918 = s3 ? tmp36919 : tmp36925;
  assign tmp36941 = l1 ? tmp35768 : tmp36924;
  assign tmp36940 = s0 ? tmp36941 : tmp36456;
  assign tmp36942 = ~(s0 ? tmp36920 : tmp36928);
  assign tmp36939 = s1 ? tmp36940 : tmp36942;
  assign tmp36944 = s0 ? tmp36920 : tmp36115;
  assign tmp36945 = l1 ? tmp35724 : tmp35833;
  assign tmp36943 = ~(s1 ? tmp36944 : tmp36945);
  assign tmp36938 = s2 ? tmp36939 : tmp36943;
  assign tmp36947 = s1 ? tmp36103 : tmp36853;
  assign tmp36951 = l2 ? tmp35716 : tmp35725;
  assign tmp36950 = ~(l1 ? tmp35904 : tmp36951);
  assign tmp36949 = s0 ? tmp36932 : tmp36950;
  assign tmp36954 = l2 ? tmp35724 : tmp35716;
  assign tmp36953 = l1 ? tmp35777 : tmp36954;
  assign tmp36952 = s0 ? tmp36953 : tmp36932;
  assign tmp36948 = s1 ? tmp36949 : tmp36952;
  assign tmp36946 = s2 ? tmp36947 : tmp36948;
  assign tmp36937 = ~(s3 ? tmp36938 : tmp36946);
  assign tmp36917 = s4 ? tmp36918 : tmp36937;
  assign tmp36960 = s0 ? tmp36923 : tmp36474;
  assign tmp36959 = s1 ? tmp36960 : tmp36603;
  assign tmp36962 = l1 ? tmp35904 : tmp35833;
  assign tmp36964 = l1 ? tmp35904 : tmp36951;
  assign tmp36963 = s0 ? tmp36964 : tmp35775;
  assign tmp36961 = ~(s1 ? tmp36962 : tmp36963);
  assign tmp36958 = s2 ? tmp36959 : tmp36961;
  assign tmp36967 = l1 ? tmp35777 : tmp36929;
  assign tmp36966 = s1 ? tmp36077 : tmp36967;
  assign tmp36969 = s0 ? tmp36953 : tmp35850;
  assign tmp36972 = l2 ? tmp35724 : tmp35727;
  assign tmp36971 = l1 ? tmp35777 : tmp36972;
  assign tmp36970 = s0 ? tmp36932 : tmp36971;
  assign tmp36968 = s1 ? tmp36969 : tmp36970;
  assign tmp36965 = s2 ? tmp36966 : tmp36968;
  assign tmp36957 = s3 ? tmp36958 : tmp36965;
  assign tmp36976 = s0 ? tmp36883 : tmp36932;
  assign tmp36977 = ~(s0 ? tmp36147 : tmp36945);
  assign tmp36975 = s1 ? tmp36976 : tmp36977;
  assign tmp36978 = ~(l1 ? tmp35914 : tmp35833);
  assign tmp36974 = s2 ? tmp36975 : tmp36978;
  assign tmp36983 = ~(l2 ? tmp35716 : tmp35720);
  assign tmp36982 = l1 ? 1 : tmp36983;
  assign tmp36984 = l1 ? tmp35821 : tmp36972;
  assign tmp36981 = s0 ? tmp36982 : tmp36984;
  assign tmp36985 = ~(l1 ? tmp35926 : tmp36894);
  assign tmp36980 = s1 ? tmp36981 : tmp36985;
  assign tmp36979 = s2 ? tmp36980 : tmp36895;
  assign tmp36973 = s3 ? tmp36974 : tmp36979;
  assign tmp36956 = s4 ? tmp36957 : tmp36973;
  assign tmp36990 = s0 ? tmp36967 : tmp35850;
  assign tmp36991 = ~(l1 ? tmp35857 : tmp35833);
  assign tmp36989 = s1 ? tmp36990 : tmp36991;
  assign tmp36988 = s2 ? tmp36989 : tmp36902;
  assign tmp36987 = s3 ? tmp36988 : tmp36904;
  assign tmp36995 = ~(l1 ? tmp35777 : tmp36954);
  assign tmp36994 = s1 ? tmp35856 : tmp36995;
  assign tmp36993 = s2 ? tmp36994 : tmp36914;
  assign tmp36992 = ~(s3 ? tmp36993 : tmp36913);
  assign tmp36986 = s4 ? tmp36987 : tmp36992;
  assign tmp36955 = ~(s5 ? tmp36956 : tmp36986);
  assign tmp36916 = s6 ? tmp36917 : tmp36955;
  assign tmp36915 = s7 ? tmp35709 : tmp36916;
  assign tmp36820 = s8 ? tmp36821 : tmp36915;
  assign tmp36819 = s9 ? tmp36820 : tmp36915;
  assign tmp36997 = s8 ? tmp36915 : tmp35709;
  assign tmp37005 = s1 ? tmp36889 : tmp36985;
  assign tmp37004 = s2 ? tmp37005 : tmp36895;
  assign tmp37003 = s3 ? tmp36880 : tmp37004;
  assign tmp37002 = s4 ? tmp36862 : tmp37003;
  assign tmp37001 = ~(s5 ? tmp37002 : tmp36896);
  assign tmp37000 = s6 ? tmp36823 : tmp37001;
  assign tmp37011 = ~(l2 ? tmp35715 : tmp35716);
  assign tmp37010 = l1 ? tmp35904 : tmp37011;
  assign tmp37014 = l2 ? tmp35724 : tmp35778;
  assign tmp37013 = l1 ? tmp35908 : tmp37014;
  assign tmp37012 = ~(s0 ? tmp36103 : tmp37013);
  assign tmp37009 = s1 ? tmp37010 : tmp37012;
  assign tmp37019 = ~(l2 ? tmp35716 : tmp35717);
  assign tmp37018 = ~(l1 ? tmp36098 : tmp37019);
  assign tmp37017 = s0 ? tmp36441 : tmp37018;
  assign tmp37021 = l1 ? tmp36098 : tmp37019;
  assign tmp37020 = ~(s0 ? tmp36103 : tmp37021);
  assign tmp37016 = s1 ? tmp37017 : tmp37020;
  assign tmp37023 = s0 ? tmp36103 : tmp36582;
  assign tmp37025 = ~(l1 ? tmp35904 : tmp37011);
  assign tmp37024 = s0 ? tmp37021 : tmp37025;
  assign tmp37022 = ~(s1 ? tmp37023 : tmp37024);
  assign tmp37015 = s2 ? tmp37016 : tmp37022;
  assign tmp37008 = s3 ? tmp37009 : tmp37015;
  assign tmp37030 = l1 ? tmp35768 : tmp37014;
  assign tmp37029 = s0 ? tmp37030 : tmp36456;
  assign tmp37031 = ~(s0 ? tmp37010 : tmp37018);
  assign tmp37028 = s1 ? tmp37029 : tmp37031;
  assign tmp37033 = s0 ? tmp37010 : tmp36115;
  assign tmp37032 = ~(s1 ? tmp37033 : tmp36945);
  assign tmp37027 = s2 ? tmp37028 : tmp37032;
  assign tmp37038 = l2 ? tmp35716 : tmp35717;
  assign tmp37037 = ~(l1 ? tmp35904 : tmp37038);
  assign tmp37036 = s0 ? tmp37021 : tmp37037;
  assign tmp37039 = s0 ? tmp36953 : tmp37021;
  assign tmp37035 = s1 ? tmp37036 : tmp37039;
  assign tmp37034 = s2 ? tmp36947 : tmp37035;
  assign tmp37026 = ~(s3 ? tmp37027 : tmp37034);
  assign tmp37007 = s4 ? tmp37008 : tmp37026;
  assign tmp37045 = s0 ? tmp37013 : tmp36474;
  assign tmp37044 = s1 ? tmp37045 : tmp36475;
  assign tmp37047 = l1 ? tmp35904 : tmp35865;
  assign tmp37049 = l1 ? tmp35904 : tmp37038;
  assign tmp37048 = s0 ? tmp37049 : tmp35775;
  assign tmp37046 = ~(s1 ? tmp37047 : tmp37048);
  assign tmp37043 = s2 ? tmp37044 : tmp37046;
  assign tmp37052 = l1 ? tmp35777 : tmp37019;
  assign tmp37051 = s1 ? tmp35887 : tmp37052;
  assign tmp37054 = s0 ? tmp37021 : tmp36953;
  assign tmp37053 = s1 ? tmp36969 : tmp37054;
  assign tmp37050 = s2 ? tmp37051 : tmp37053;
  assign tmp37042 = s3 ? tmp37043 : tmp37050;
  assign tmp37058 = s0 ? tmp36883 : tmp37021;
  assign tmp37057 = s1 ? tmp37058 : tmp36977;
  assign tmp37059 = ~(l1 ? tmp35914 : tmp35865);
  assign tmp37056 = s2 ? tmp37057 : tmp37059;
  assign tmp37064 = ~(l2 ? tmp35716 : tmp36091);
  assign tmp37063 = l1 ? 1 : tmp37064;
  assign tmp37065 = l1 ? tmp35821 : tmp36954;
  assign tmp37062 = s0 ? tmp37063 : tmp37065;
  assign tmp37067 = l2 ? tmp35716 : tmp35724;
  assign tmp37066 = ~(l1 ? tmp35926 : tmp37067);
  assign tmp37061 = s1 ? tmp37062 : tmp37066;
  assign tmp37060 = s2 ? tmp37061 : tmp36895;
  assign tmp37055 = s3 ? tmp37056 : tmp37060;
  assign tmp37041 = s4 ? tmp37042 : tmp37055;
  assign tmp37072 = s0 ? tmp37052 : tmp35850;
  assign tmp37071 = s1 ? tmp37072 : tmp36991;
  assign tmp37073 = s1 ? tmp36502 : tmp35995;
  assign tmp37070 = s2 ? tmp37071 : tmp37073;
  assign tmp37076 = ~(l1 ? 1 : tmp35779);
  assign tmp37075 = s1 ? tmp36906 : tmp37076;
  assign tmp37074 = ~(s2 ? tmp35997 : tmp37075);
  assign tmp37069 = s3 ? tmp37070 : tmp37074;
  assign tmp37079 = l1 ? tmp35926 : tmp35865;
  assign tmp37078 = s2 ? tmp36994 : tmp37079;
  assign tmp37080 = s1 ? tmp36008 : tmp37079;
  assign tmp37077 = ~(s3 ? tmp37078 : tmp37080);
  assign tmp37068 = s4 ? tmp37069 : tmp37077;
  assign tmp37040 = ~(s5 ? tmp37041 : tmp37068);
  assign tmp37006 = s6 ? tmp37007 : tmp37040;
  assign tmp36999 = s7 ? tmp37000 : tmp37006;
  assign tmp36998 = s8 ? tmp36999 : tmp36916;
  assign tmp36996 = s9 ? tmp36997 : tmp36998;
  assign tmp36818 = s10 ? tmp36819 : tmp36996;
  assign tmp37084 = s7 ? tmp36822 : tmp37006;
  assign tmp37083 = s8 ? tmp37084 : tmp36916;
  assign tmp37082 = s9 ? tmp36997 : tmp37083;
  assign tmp37081 = s10 ? tmp36819 : tmp37082;
  assign tmp36817 = s11 ? tmp36818 : tmp37081;
  assign tmp36635 = s12 ? tmp36636 : tmp36817;
  assign tmp37095 = l1 ? tmp35714 : tmp35768;
  assign tmp37097 = l1 ? tmp35729 : tmp35909;
  assign tmp37096 = ~(s0 ? tmp35906 : tmp37097);
  assign tmp37094 = s1 ? tmp37095 : tmp37096;
  assign tmp37101 = ~(l1 ? tmp35739 : tmp35917);
  assign tmp37100 = s0 ? tmp35735 : tmp37101;
  assign tmp37103 = l1 ? tmp35743 : tmp35920;
  assign tmp37104 = l1 ? tmp35739 : tmp35917;
  assign tmp37102 = ~(s0 ? tmp37103 : tmp37104);
  assign tmp37099 = s1 ? tmp37100 : tmp37102;
  assign tmp37106 = s0 ? tmp37103 : tmp35749;
  assign tmp37108 = ~(l1 ? tmp35714 : tmp35768);
  assign tmp37107 = s0 ? tmp37104 : tmp37108;
  assign tmp37105 = ~(s1 ? tmp37106 : tmp37107);
  assign tmp37098 = s2 ? tmp37099 : tmp37105;
  assign tmp37093 = s3 ? tmp37094 : tmp37098;
  assign tmp37113 = l1 ? tmp35743 : tmp35909;
  assign tmp37112 = s0 ? tmp37113 : tmp35757;
  assign tmp37114 = ~(s0 ? tmp37095 : tmp37101);
  assign tmp37111 = s1 ? tmp37112 : tmp37114;
  assign tmp37116 = s0 ? tmp37095 : tmp36115;
  assign tmp37115 = ~(s1 ? tmp37116 : tmp35823);
  assign tmp37110 = s2 ? tmp37111 : tmp37115;
  assign tmp37120 = ~(l1 ? tmp35714 : tmp35942);
  assign tmp37119 = s0 ? tmp37104 : tmp37120;
  assign tmp37122 = l1 ? tmp35786 : tmp35945;
  assign tmp37121 = s0 ? tmp37122 : tmp37104;
  assign tmp37118 = s1 ? tmp37119 : tmp37121;
  assign tmp37117 = s2 ? tmp35937 : tmp37118;
  assign tmp37109 = ~(s3 ? tmp37110 : tmp37117);
  assign tmp37092 = s4 ? tmp37093 : tmp37109;
  assign tmp37128 = s0 ? tmp37097 : tmp35793;
  assign tmp37129 = ~(l1 ? tmp35736 : tmp35737);
  assign tmp37127 = s1 ? tmp37128 : tmp37129;
  assign tmp37131 = l1 ? tmp35714 : tmp35955;
  assign tmp37133 = l1 ? tmp35714 : tmp35942;
  assign tmp37132 = s0 ? tmp37133 : tmp35801;
  assign tmp37130 = ~(s1 ? tmp37131 : tmp37132);
  assign tmp37126 = s2 ? tmp37127 : tmp37130;
  assign tmp37136 = l1 ? tmp35806 : tmp35920;
  assign tmp37137 = l1 ? tmp35786 : tmp35917;
  assign tmp37135 = s1 ? tmp37136 : tmp37137;
  assign tmp37139 = s0 ? tmp37122 : tmp35850;
  assign tmp37141 = l1 ? tmp35815 : tmp35917;
  assign tmp37140 = s0 ? tmp37104 : tmp37141;
  assign tmp37138 = s1 ? tmp37139 : tmp37140;
  assign tmp37134 = s2 ? tmp37135 : tmp37138;
  assign tmp37125 = s3 ? tmp37126 : tmp37134;
  assign tmp37146 = l1 ? tmp35739 : tmp35973;
  assign tmp37145 = s0 ? tmp35971 : tmp37146;
  assign tmp37144 = s1 ? tmp37145 : tmp35974;
  assign tmp37147 = ~(l1 ? tmp35736 : tmp35955);
  assign tmp37143 = s2 ? tmp37144 : tmp37147;
  assign tmp37151 = l1 ? tmp35833 : tmp35982;
  assign tmp37152 = l1 ? tmp35835 : tmp35973;
  assign tmp37150 = s0 ? tmp37151 : tmp37152;
  assign tmp37153 = ~(l1 ? tmp35714 : tmp35821);
  assign tmp37149 = s1 ? tmp37150 : tmp37153;
  assign tmp37148 = s2 ? tmp37149 : tmp35985;
  assign tmp37142 = s3 ? tmp37143 : tmp37148;
  assign tmp37124 = s4 ? tmp37125 : tmp37142;
  assign tmp37158 = s0 ? tmp37137 : tmp35850;
  assign tmp37157 = s1 ? tmp37158 : tmp35879;
  assign tmp37160 = l1 ? tmp35833 : tmp35736;
  assign tmp37161 = ~(s0 ? tmp35827 : tmp35860);
  assign tmp37159 = s1 ? tmp37160 : tmp37161;
  assign tmp37156 = s2 ? tmp37157 : tmp37159;
  assign tmp37164 = s0 ? tmp35864 : 1;
  assign tmp37163 = s1 ? tmp37164 : tmp35998;
  assign tmp37166 = ~(l1 ? tmp35833 : tmp35982);
  assign tmp37165 = s1 ? tmp36000 : tmp37166;
  assign tmp37162 = ~(s2 ? tmp37163 : tmp37165);
  assign tmp37155 = s3 ? tmp37156 : tmp37162;
  assign tmp37170 = ~(l1 ? tmp35786 : tmp35945);
  assign tmp37169 = s1 ? tmp36000 : tmp37170;
  assign tmp37171 = s1 ? tmp37131 : tmp35886;
  assign tmp37168 = s2 ? tmp37169 : tmp37171;
  assign tmp37173 = l1 ? tmp35812 : tmp35821;
  assign tmp37174 = l1 ? tmp35714 : 1;
  assign tmp37172 = s1 ? tmp37173 : tmp37174;
  assign tmp37167 = ~(s3 ? tmp37168 : tmp37172);
  assign tmp37154 = s4 ? tmp37155 : tmp37167;
  assign tmp37123 = ~(s5 ? tmp37124 : tmp37154);
  assign tmp37091 = s6 ? tmp37092 : tmp37123;
  assign tmp37090 = s7 ? tmp35709 : tmp37091;
  assign tmp37181 = l2 ? tmp35724 : tmp35715;
  assign tmp37180 = l1 ? tmp37181 : tmp35723;
  assign tmp37184 = l2 ? tmp35778 : tmp35730;
  assign tmp37183 = l1 ? tmp37184 : tmp36751;
  assign tmp37182 = ~(s0 ? tmp36679 : tmp37183);
  assign tmp37179 = s1 ? tmp37180 : tmp37182;
  assign tmp37188 = l1 ? tmp35724 : tmp35737;
  assign tmp37190 = l2 ? tmp35716 : tmp35730;
  assign tmp37189 = ~(l1 ? tmp37190 : tmp35917);
  assign tmp37187 = s0 ? tmp37188 : tmp37189;
  assign tmp37193 = l2 ? tmp35778 : tmp35725;
  assign tmp37192 = l1 ? tmp37193 : tmp36758;
  assign tmp37194 = l1 ? tmp37190 : tmp35917;
  assign tmp37191 = ~(s0 ? tmp37192 : tmp37194);
  assign tmp37186 = s1 ? tmp37187 : tmp37191;
  assign tmp37196 = s0 ? tmp37192 : tmp36652;
  assign tmp37198 = ~(l1 ? tmp37181 : tmp35723);
  assign tmp37197 = s0 ? tmp37194 : tmp37198;
  assign tmp37195 = ~(s1 ? tmp37196 : tmp37197);
  assign tmp37185 = s2 ? tmp37186 : tmp37195;
  assign tmp37178 = s3 ? tmp37179 : tmp37185;
  assign tmp37203 = l1 ? tmp37193 : tmp36751;
  assign tmp37202 = s0 ? tmp37203 : tmp36111;
  assign tmp37204 = ~(s0 ? tmp37180 : tmp37189);
  assign tmp37201 = s1 ? tmp37202 : tmp37204;
  assign tmp37206 = s0 ? tmp37180 : tmp36115;
  assign tmp37205 = ~(s1 ? tmp37206 : tmp36698);
  assign tmp37200 = s2 ? tmp37201 : tmp37205;
  assign tmp37210 = ~(l1 ? tmp37181 : tmp35942);
  assign tmp37209 = s0 ? tmp37194 : tmp37210;
  assign tmp37212 = l1 ? tmp35786 : tmp35882;
  assign tmp37211 = s0 ? tmp37212 : tmp37194;
  assign tmp37208 = s1 ? tmp37209 : tmp37211;
  assign tmp37207 = s2 ? tmp36700 : tmp37208;
  assign tmp37199 = ~(s3 ? tmp37200 : tmp37207);
  assign tmp37177 = s4 ? tmp37178 : tmp37199;
  assign tmp37218 = s0 ? tmp37183 : tmp35793;
  assign tmp37219 = ~(l1 ? tmp35724 : tmp35737);
  assign tmp37217 = s1 ? tmp37218 : tmp37219;
  assign tmp37221 = l1 ? tmp37181 : tmp35955;
  assign tmp37223 = l1 ? tmp37181 : tmp35942;
  assign tmp37222 = s0 ? tmp37223 : tmp36716;
  assign tmp37220 = ~(s1 ? tmp37221 : tmp37222);
  assign tmp37216 = s2 ? tmp37217 : tmp37220;
  assign tmp37226 = l1 ? tmp35833 : tmp36758;
  assign tmp37225 = s1 ? tmp37226 : tmp37137;
  assign tmp37228 = s0 ? tmp37212 : tmp35850;
  assign tmp37229 = s0 ? tmp37194 : tmp37137;
  assign tmp37227 = s1 ? tmp37228 : tmp37229;
  assign tmp37224 = s2 ? tmp37225 : tmp37227;
  assign tmp37215 = s3 ? tmp37216 : tmp37224;
  assign tmp37233 = s0 ? tmp35971 : tmp37194;
  assign tmp37232 = s1 ? tmp37233 : tmp36726;
  assign tmp37234 = ~(l1 ? tmp35724 : tmp35955);
  assign tmp37231 = s2 ? tmp37232 : tmp37234;
  assign tmp37238 = l1 ? tmp36894 : tmp35917;
  assign tmp37237 = s0 ? tmp37151 : tmp37238;
  assign tmp37236 = s1 ? tmp37237 : tmp37153;
  assign tmp37235 = s2 ? tmp37236 : tmp35985;
  assign tmp37230 = s3 ? tmp37231 : tmp37235;
  assign tmp37214 = s4 ? tmp37215 : tmp37230;
  assign tmp37243 = ~(l1 ? tmp35812 : tmp35767);
  assign tmp37242 = s1 ? tmp37158 : tmp37243;
  assign tmp37244 = s1 ? tmp37160 : tmp36560;
  assign tmp37241 = s2 ? tmp37242 : tmp37244;
  assign tmp37240 = s3 ? tmp37241 : tmp37162;
  assign tmp37248 = ~(l1 ? tmp35786 : tmp35882);
  assign tmp37247 = s1 ? tmp36000 : tmp37248;
  assign tmp37249 = s1 ? tmp37131 : tmp35864;
  assign tmp37246 = s2 ? tmp37247 : tmp37249;
  assign tmp37245 = ~(s3 ? tmp37246 : tmp37172);
  assign tmp37239 = s4 ? tmp37240 : tmp37245;
  assign tmp37213 = ~(s5 ? tmp37214 : tmp37239);
  assign tmp37176 = s6 ? tmp37177 : tmp37213;
  assign tmp37175 = s7 ? tmp35709 : tmp37176;
  assign tmp37089 = s8 ? tmp37090 : tmp37175;
  assign tmp37256 = l1 ? tmp37181 : tmp35773;
  assign tmp37258 = l1 ? tmp37184 : tmp36090;
  assign tmp37257 = ~(s0 ? tmp36088 : tmp37258);
  assign tmp37255 = s1 ? tmp37256 : tmp37257;
  assign tmp37262 = l1 ? tmp35724 : tmp35725;
  assign tmp37263 = ~(l1 ? tmp37190 : tmp35945);
  assign tmp37261 = s0 ? tmp37262 : tmp37263;
  assign tmp37265 = l1 ? tmp37193 : tmp35764;
  assign tmp37266 = l1 ? tmp37190 : tmp35945;
  assign tmp37264 = ~(s0 ? tmp37265 : tmp37266);
  assign tmp37260 = s1 ? tmp37261 : tmp37264;
  assign tmp37268 = s0 ? tmp37265 : tmp36103;
  assign tmp37270 = ~(l1 ? tmp37181 : tmp35773);
  assign tmp37269 = s0 ? tmp37266 : tmp37270;
  assign tmp37267 = ~(s1 ? tmp37268 : tmp37269);
  assign tmp37259 = s2 ? tmp37260 : tmp37267;
  assign tmp37254 = s3 ? tmp37255 : tmp37259;
  assign tmp37275 = l1 ? tmp37193 : tmp36090;
  assign tmp37274 = s0 ? tmp37275 : tmp36111;
  assign tmp37276 = ~(s0 ? tmp37256 : tmp37263);
  assign tmp37273 = s1 ? tmp37274 : tmp37276;
  assign tmp37278 = s0 ? tmp37256 : tmp36115;
  assign tmp37277 = ~(s1 ? tmp37278 : tmp36116);
  assign tmp37272 = s2 ? tmp37273 : tmp37277;
  assign tmp37282 = ~(l1 ? tmp37181 : tmp36122);
  assign tmp37281 = s0 ? tmp37266 : tmp37282;
  assign tmp37283 = s0 ? tmp37122 : tmp37266;
  assign tmp37280 = s1 ? tmp37281 : tmp37283;
  assign tmp37279 = s2 ? tmp36118 : tmp37280;
  assign tmp37271 = ~(s3 ? tmp37272 : tmp37279);
  assign tmp37253 = s4 ? tmp37254 : tmp37271;
  assign tmp37289 = s0 ? tmp37258 : tmp35793;
  assign tmp37288 = s1 ? tmp37289 : tmp36111;
  assign tmp37291 = l1 ? tmp37181 : tmp35744;
  assign tmp37293 = l1 ? tmp37181 : tmp36122;
  assign tmp37292 = s0 ? tmp37293 : tmp36135;
  assign tmp37290 = ~(s1 ? tmp37291 : tmp37292);
  assign tmp37287 = s2 ? tmp37288 : tmp37290;
  assign tmp37296 = l1 ? tmp35833 : tmp35764;
  assign tmp37295 = s1 ? tmp37296 : tmp37122;
  assign tmp37298 = s0 ? tmp37266 : tmp37122;
  assign tmp37297 = s1 ? tmp37139 : tmp37298;
  assign tmp37294 = s2 ? tmp37295 : tmp37297;
  assign tmp37286 = s3 ? tmp37287 : tmp37294;
  assign tmp37302 = s0 ? tmp35971 : tmp37266;
  assign tmp37301 = s1 ? tmp37302 : tmp36146;
  assign tmp37303 = ~(l1 ? tmp35724 : tmp35744);
  assign tmp37300 = s2 ? tmp37301 : tmp37303;
  assign tmp37307 = l1 ? tmp35833 : tmp36153;
  assign tmp37308 = l1 ? tmp36894 : tmp35945;
  assign tmp37306 = s0 ? tmp37307 : tmp37308;
  assign tmp37309 = ~(l1 ? tmp35714 : tmp36288);
  assign tmp37305 = s1 ? tmp37306 : tmp37309;
  assign tmp37304 = s2 ? tmp37305 : tmp35985;
  assign tmp37299 = s3 ? tmp37300 : tmp37304;
  assign tmp37285 = s4 ? tmp37286 : tmp37299;
  assign tmp37313 = s1 ? tmp37139 : tmp35879;
  assign tmp37315 = l1 ? tmp35833 : tmp35767;
  assign tmp37314 = s1 ? tmp37315 : tmp36560;
  assign tmp37312 = s2 ? tmp37313 : tmp37314;
  assign tmp37318 = ~(l1 ? tmp35833 : tmp35778);
  assign tmp37317 = s1 ? tmp36000 : tmp37318;
  assign tmp37316 = ~(s2 ? tmp37163 : tmp37317);
  assign tmp37311 = s3 ? tmp37312 : tmp37316;
  assign tmp37322 = l1 ? tmp35714 : tmp35744;
  assign tmp37321 = s1 ? tmp37322 : tmp35864;
  assign tmp37320 = s2 ? tmp37169 : tmp37321;
  assign tmp37324 = l1 ? tmp35714 : tmp35736;
  assign tmp37323 = s1 ? tmp37173 : tmp37324;
  assign tmp37319 = ~(s3 ? tmp37320 : tmp37323);
  assign tmp37310 = s4 ? tmp37311 : tmp37319;
  assign tmp37284 = ~(s5 ? tmp37285 : tmp37310);
  assign tmp37252 = s6 ? tmp37253 : tmp37284;
  assign tmp37251 = s7 ? tmp35709 : tmp37252;
  assign tmp37250 = s8 ? tmp37175 : tmp37251;
  assign tmp37088 = s9 ? tmp37089 : tmp37250;
  assign tmp37332 = l1 ? tmp37181 : tmp35768;
  assign tmp37334 = l1 ? tmp37184 : tmp35909;
  assign tmp37333 = ~(s0 ? tmp36088 : tmp37334);
  assign tmp37331 = s1 ? tmp37332 : tmp37333;
  assign tmp37338 = ~(l1 ? tmp37190 : tmp35973);
  assign tmp37337 = s0 ? tmp37262 : tmp37338;
  assign tmp37340 = l1 ? tmp37193 : tmp35920;
  assign tmp37341 = l1 ? tmp37190 : tmp35973;
  assign tmp37339 = ~(s0 ? tmp37340 : tmp37341);
  assign tmp37336 = s1 ? tmp37337 : tmp37339;
  assign tmp37343 = s0 ? tmp37340 : tmp36103;
  assign tmp37345 = ~(l1 ? tmp37181 : tmp35768);
  assign tmp37344 = s0 ? tmp37341 : tmp37345;
  assign tmp37342 = ~(s1 ? tmp37343 : tmp37344);
  assign tmp37335 = s2 ? tmp37336 : tmp37342;
  assign tmp37330 = s3 ? tmp37331 : tmp37335;
  assign tmp37350 = l1 ? tmp37193 : tmp35909;
  assign tmp37349 = s0 ? tmp37350 : tmp36111;
  assign tmp37351 = ~(s0 ? tmp37332 : tmp37338);
  assign tmp37348 = s1 ? tmp37349 : tmp37351;
  assign tmp37353 = s0 ? tmp37332 : tmp36115;
  assign tmp37352 = ~(s1 ? tmp37353 : tmp36116);
  assign tmp37347 = s2 ? tmp37348 : tmp37352;
  assign tmp37357 = ~(l1 ? tmp37181 : tmp36041);
  assign tmp37356 = s0 ? tmp37341 : tmp37357;
  assign tmp37358 = s0 ? tmp37122 : tmp37341;
  assign tmp37355 = s1 ? tmp37356 : tmp37358;
  assign tmp37354 = s2 ? tmp36118 : tmp37355;
  assign tmp37346 = ~(s3 ? tmp37347 : tmp37354);
  assign tmp37329 = s4 ? tmp37330 : tmp37346;
  assign tmp37364 = s0 ? tmp37334 : tmp35793;
  assign tmp37363 = s1 ? tmp37364 : tmp36111;
  assign tmp37366 = l1 ? tmp37181 : tmp35726;
  assign tmp37368 = l1 ? tmp37181 : tmp36041;
  assign tmp37367 = s0 ? tmp37368 : tmp36135;
  assign tmp37365 = ~(s1 ? tmp37366 : tmp37367);
  assign tmp37362 = s2 ? tmp37363 : tmp37365;
  assign tmp37371 = l1 ? tmp35833 : tmp35920;
  assign tmp37372 = l1 ? tmp35786 : tmp35973;
  assign tmp37370 = s1 ? tmp37371 : tmp37372;
  assign tmp37374 = s0 ? tmp37341 : tmp37372;
  assign tmp37373 = s1 ? tmp37139 : tmp37374;
  assign tmp37369 = s2 ? tmp37370 : tmp37373;
  assign tmp37361 = s3 ? tmp37362 : tmp37369;
  assign tmp37378 = s0 ? tmp35971 : tmp37341;
  assign tmp37377 = s1 ? tmp37378 : tmp36146;
  assign tmp37379 = ~(l1 ? tmp35724 : tmp35726);
  assign tmp37376 = s2 ? tmp37377 : tmp37379;
  assign tmp37383 = l1 ? tmp35833 : tmp35719;
  assign tmp37384 = l1 ? tmp36894 : tmp35973;
  assign tmp37382 = s0 ? tmp37383 : tmp37384;
  assign tmp37381 = s1 ? tmp37382 : tmp37153;
  assign tmp37380 = s2 ? tmp37381 : tmp35985;
  assign tmp37375 = s3 ? tmp37376 : tmp37380;
  assign tmp37360 = s4 ? tmp37361 : tmp37375;
  assign tmp37389 = s0 ? tmp37372 : tmp35850;
  assign tmp37388 = s1 ? tmp37389 : tmp35879;
  assign tmp37391 = l1 ? tmp35833 : tmp35724;
  assign tmp37390 = s1 ? tmp37391 : tmp36560;
  assign tmp37387 = s2 ? tmp37388 : tmp37390;
  assign tmp37386 = s3 ? tmp37387 : tmp37162;
  assign tmp37395 = l1 ? tmp35714 : tmp35726;
  assign tmp37394 = s1 ? tmp37395 : tmp35864;
  assign tmp37393 = s2 ? tmp37169 : tmp37394;
  assign tmp37392 = ~(s3 ? tmp37393 : tmp37172);
  assign tmp37385 = s4 ? tmp37386 : tmp37392;
  assign tmp37359 = ~(s5 ? tmp37360 : tmp37385);
  assign tmp37328 = s6 ? tmp37329 : tmp37359;
  assign tmp37327 = s7 ? tmp35709 : tmp37328;
  assign tmp37326 = s8 ? tmp37327 : tmp35709;
  assign tmp37402 = s2 ? tmp37169 : tmp37131;
  assign tmp37401 = ~(s3 ? tmp37402 : tmp37172);
  assign tmp37400 = s4 ? tmp37155 : tmp37401;
  assign tmp37399 = ~(s5 ? tmp37124 : tmp37400);
  assign tmp37398 = s6 ? tmp37092 : tmp37399;
  assign tmp37407 = s2 ? tmp37169 : tmp37322;
  assign tmp37406 = ~(s3 ? tmp37407 : tmp37323);
  assign tmp37405 = s4 ? tmp37311 : tmp37406;
  assign tmp37404 = ~(s5 ? tmp37285 : tmp37405);
  assign tmp37403 = s6 ? tmp37253 : tmp37404;
  assign tmp37397 = s7 ? tmp37398 : tmp37403;
  assign tmp37413 = s2 ? tmp37247 : tmp37131;
  assign tmp37412 = ~(s3 ? tmp37413 : tmp37172);
  assign tmp37411 = s4 ? tmp37240 : tmp37412;
  assign tmp37410 = ~(s5 ? tmp37214 : tmp37411);
  assign tmp37409 = s6 ? tmp37177 : tmp37410;
  assign tmp37418 = s2 ? tmp37169 : tmp37395;
  assign tmp37417 = ~(s3 ? tmp37418 : tmp37172);
  assign tmp37416 = s4 ? tmp37386 : tmp37417;
  assign tmp37415 = ~(s5 ? tmp37360 : tmp37416);
  assign tmp37414 = s6 ? tmp37329 : tmp37415;
  assign tmp37408 = s7 ? tmp37409 : tmp37414;
  assign tmp37396 = s8 ? tmp37397 : tmp37408;
  assign tmp37325 = s9 ? tmp37326 : tmp37396;
  assign tmp37087 = s10 ? tmp37088 : tmp37325;
  assign tmp37422 = s7 ? tmp37091 : tmp37252;
  assign tmp37423 = s7 ? tmp37176 : tmp37328;
  assign tmp37421 = s8 ? tmp37422 : tmp37423;
  assign tmp37420 = s9 ? tmp37326 : tmp37421;
  assign tmp37419 = s10 ? tmp37088 : tmp37420;
  assign tmp37086 = s11 ? tmp37087 : tmp37419;
  assign tmp37433 = l1 ? tmp35714 : tmp35725;
  assign tmp37435 = l1 ? tmp35729 : tmp35982;
  assign tmp37434 = ~(s0 ? tmp36512 : tmp37435);
  assign tmp37432 = s1 ? tmp37433 : tmp37434;
  assign tmp37439 = l1 ? tmp35736 : tmp35723;
  assign tmp37441 = ~(l2 ? tmp35715 : tmp35725);
  assign tmp37440 = ~(l1 ? tmp35739 : tmp37441);
  assign tmp37438 = s0 ? tmp37439 : tmp37440;
  assign tmp37443 = l1 ? tmp35743 : tmp35914;
  assign tmp37444 = l1 ? tmp35739 : tmp37441;
  assign tmp37442 = ~(s0 ? tmp37443 : tmp37444);
  assign tmp37437 = s1 ? tmp37438 : tmp37442;
  assign tmp37446 = s0 ? tmp37443 : tmp36582;
  assign tmp37448 = ~(l1 ? tmp35714 : tmp35725);
  assign tmp37447 = s0 ? tmp37444 : tmp37448;
  assign tmp37445 = ~(s1 ? tmp37446 : tmp37447);
  assign tmp37436 = s2 ? tmp37437 : tmp37445;
  assign tmp37431 = s3 ? tmp37432 : tmp37436;
  assign tmp37453 = l1 ? tmp35743 : tmp35982;
  assign tmp37452 = s0 ? tmp37453 : tmp36530;
  assign tmp37454 = ~(s0 ? tmp37433 : tmp37440);
  assign tmp37451 = s1 ? tmp37452 : tmp37454;
  assign tmp37456 = s0 ? tmp37433 : tmp36115;
  assign tmp37455 = ~(s1 ? tmp37456 : tmp35827);
  assign tmp37450 = s2 ? tmp37451 : tmp37455;
  assign tmp37461 = l2 ? tmp35715 : tmp35725;
  assign tmp37460 = ~(l1 ? tmp35714 : tmp37461);
  assign tmp37459 = s0 ? tmp37444 : tmp37460;
  assign tmp37462 = s0 ? tmp37122 : tmp37444;
  assign tmp37458 = s1 ? tmp37459 : tmp37462;
  assign tmp37457 = s2 ? tmp36535 : tmp37458;
  assign tmp37449 = ~(s3 ? tmp37450 : tmp37457);
  assign tmp37430 = s4 ? tmp37431 : tmp37449;
  assign tmp37468 = s0 ? tmp37435 : tmp36474;
  assign tmp37469 = ~(l1 ? tmp35736 : tmp35723);
  assign tmp37467 = s1 ? tmp37468 : tmp37469;
  assign tmp37472 = l1 ? tmp35714 : tmp37461;
  assign tmp37471 = s0 ? tmp37472 : tmp35775;
  assign tmp37470 = ~(s1 ? tmp37174 : tmp37471);
  assign tmp37466 = s2 ? tmp37467 : tmp37470;
  assign tmp37475 = l1 ? tmp35806 : tmp35914;
  assign tmp37476 = l1 ? tmp35786 : tmp36576;
  assign tmp37474 = s1 ? tmp37475 : tmp37476;
  assign tmp37479 = l1 ? tmp35739 : tmp36576;
  assign tmp37478 = s0 ? tmp37479 : tmp37141;
  assign tmp37477 = s1 ? tmp37139 : tmp37478;
  assign tmp37473 = s2 ? tmp37474 : tmp37477;
  assign tmp37465 = s3 ? tmp37466 : tmp37473;
  assign tmp37483 = s0 ? tmp35971 : tmp37479;
  assign tmp37482 = s1 ? tmp37483 : tmp36560;
  assign tmp37481 = s2 ? tmp37482 : tmp36560;
  assign tmp37487 = l1 ? tmp35833 : tmp35909;
  assign tmp37486 = s0 ? tmp37487 : tmp37152;
  assign tmp37485 = s1 ? tmp37486 : tmp37153;
  assign tmp37484 = s2 ? tmp37485 : tmp35985;
  assign tmp37480 = s3 ? tmp37481 : tmp37484;
  assign tmp37464 = s4 ? tmp37465 : tmp37480;
  assign tmp37492 = s0 ? tmp37476 : tmp35850;
  assign tmp37491 = s1 ? tmp37492 : tmp35879;
  assign tmp37494 = l1 ? tmp35833 : tmp36713;
  assign tmp37493 = s1 ? tmp37494 : tmp36560;
  assign tmp37490 = s2 ? tmp37491 : tmp37493;
  assign tmp37489 = s3 ? tmp37490 : tmp37162;
  assign tmp37497 = s1 ? tmp37174 : tmp35864;
  assign tmp37496 = s2 ? tmp37169 : tmp37497;
  assign tmp37495 = ~(s3 ? tmp37496 : tmp37172);
  assign tmp37488 = s4 ? tmp37489 : tmp37495;
  assign tmp37463 = ~(s5 ? tmp37464 : tmp37488);
  assign tmp37429 = s6 ? tmp37430 : tmp37463;
  assign tmp37428 = s7 ? tmp35709 : tmp37429;
  assign tmp37503 = l1 ? tmp37181 : tmp35737;
  assign tmp37505 = l1 ? tmp35768 : tmp35833;
  assign tmp37506 = l1 ? tmp37184 : tmp35982;
  assign tmp37504 = ~(s0 ? tmp37505 : tmp37506);
  assign tmp37502 = s1 ? tmp37503 : tmp37504;
  assign tmp37510 = l1 ? tmp35724 : tmp35723;
  assign tmp37511 = ~(l1 ? tmp37190 : tmp37441);
  assign tmp37509 = s0 ? tmp37510 : tmp37511;
  assign tmp37513 = l1 ? tmp37193 : tmp35865;
  assign tmp37514 = l1 ? tmp37190 : tmp37441;
  assign tmp37512 = ~(s0 ? tmp37513 : tmp37514);
  assign tmp37508 = s1 ? tmp37509 : tmp37512;
  assign tmp37516 = s0 ? tmp37513 : tmp35795;
  assign tmp37518 = ~(l1 ? tmp37181 : tmp35737);
  assign tmp37517 = s0 ? tmp37514 : tmp37518;
  assign tmp37515 = ~(s1 ? tmp37516 : tmp37517);
  assign tmp37507 = s2 ? tmp37508 : tmp37515;
  assign tmp37501 = s3 ? tmp37502 : tmp37507;
  assign tmp37523 = l1 ? tmp37193 : tmp35982;
  assign tmp37522 = s0 ? tmp37523 : tmp36456;
  assign tmp37524 = ~(s0 ? tmp37503 : tmp37511);
  assign tmp37521 = s1 ? tmp37522 : tmp37524;
  assign tmp37526 = s0 ? tmp37503 : tmp36115;
  assign tmp37525 = ~(s1 ? tmp37526 : tmp36727);
  assign tmp37520 = s2 ? tmp37521 : tmp37525;
  assign tmp37528 = s1 ? tmp37505 : tmp35938;
  assign tmp37531 = ~(l1 ? tmp37181 : tmp37461);
  assign tmp37530 = s0 ? tmp37514 : tmp37531;
  assign tmp37532 = s0 ? tmp37212 : tmp37514;
  assign tmp37529 = s1 ? tmp37530 : tmp37532;
  assign tmp37527 = s2 ? tmp37528 : tmp37529;
  assign tmp37519 = ~(s3 ? tmp37520 : tmp37527);
  assign tmp37500 = s4 ? tmp37501 : tmp37519;
  assign tmp37538 = s0 ? tmp37506 : tmp36474;
  assign tmp37539 = ~(l1 ? tmp35724 : tmp35723);
  assign tmp37537 = s1 ? tmp37538 : tmp37539;
  assign tmp37541 = l1 ? tmp37181 : tmp35767;
  assign tmp37543 = l1 ? tmp37181 : tmp37461;
  assign tmp37544 = l1 ? tmp35767 : tmp35723;
  assign tmp37542 = s0 ? tmp37543 : tmp37544;
  assign tmp37540 = ~(s1 ? tmp37541 : tmp37542);
  assign tmp37536 = s2 ? tmp37537 : tmp37540;
  assign tmp37547 = l1 ? tmp35833 : tmp35865;
  assign tmp37548 = l1 ? tmp35786 : tmp37441;
  assign tmp37546 = s1 ? tmp37547 : tmp37548;
  assign tmp37550 = s0 ? tmp37514 : tmp37137;
  assign tmp37549 = s1 ? tmp37228 : tmp37550;
  assign tmp37545 = s2 ? tmp37546 : tmp37549;
  assign tmp37535 = s3 ? tmp37536 : tmp37545;
  assign tmp37554 = s0 ? tmp35971 : tmp37514;
  assign tmp37555 = ~(s0 ? tmp36147 : tmp36727);
  assign tmp37553 = s1 ? tmp37554 : tmp37555;
  assign tmp37556 = ~(l1 ? tmp35724 : tmp35767);
  assign tmp37552 = s2 ? tmp37553 : tmp37556;
  assign tmp37560 = l1 ? tmp35833 : tmp36751;
  assign tmp37559 = s0 ? tmp37560 : tmp37238;
  assign tmp37558 = s1 ? tmp37559 : tmp37153;
  assign tmp37557 = s2 ? tmp37558 : tmp35985;
  assign tmp37551 = s3 ? tmp37552 : tmp37557;
  assign tmp37534 = s4 ? tmp37535 : tmp37551;
  assign tmp37565 = s0 ? tmp37548 : tmp35850;
  assign tmp37564 = s1 ? tmp37565 : tmp37243;
  assign tmp37567 = l1 ? tmp35833 : tmp35744;
  assign tmp37566 = s1 ? tmp37567 : tmp36560;
  assign tmp37563 = s2 ? tmp37564 : tmp37566;
  assign tmp37562 = s3 ? tmp37563 : tmp37162;
  assign tmp37571 = l1 ? tmp35714 : tmp35767;
  assign tmp37570 = s1 ? tmp37571 : tmp35864;
  assign tmp37569 = s2 ? tmp37247 : tmp37570;
  assign tmp37568 = ~(s3 ? tmp37569 : tmp37172);
  assign tmp37561 = s4 ? tmp37562 : tmp37568;
  assign tmp37533 = ~(s5 ? tmp37534 : tmp37561);
  assign tmp37499 = s6 ? tmp37500 : tmp37533;
  assign tmp37498 = s7 ? tmp35709 : tmp37499;
  assign tmp37427 = s8 ? tmp37428 : tmp37498;
  assign tmp37578 = l1 ? tmp37181 : tmp36096;
  assign tmp37580 = l1 ? tmp37184 : tmp36153;
  assign tmp37579 = ~(s0 ? tmp36436 : tmp37580);
  assign tmp37577 = s1 ? tmp37578 : tmp37579;
  assign tmp37584 = l1 ? tmp35724 : tmp35773;
  assign tmp37585 = ~(l1 ? tmp37190 : tmp36443);
  assign tmp37583 = s0 ? tmp37584 : tmp37585;
  assign tmp37587 = l1 ? tmp37193 : tmp35806;
  assign tmp37588 = l1 ? tmp37190 : tmp36443;
  assign tmp37586 = ~(s0 ? tmp37587 : tmp37588);
  assign tmp37582 = s1 ? tmp37583 : tmp37586;
  assign tmp37590 = s0 ? tmp37587 : tmp36582;
  assign tmp37592 = ~(l1 ? tmp37181 : tmp36096);
  assign tmp37591 = s0 ? tmp37588 : tmp37592;
  assign tmp37589 = ~(s1 ? tmp37590 : tmp37591);
  assign tmp37581 = s2 ? tmp37582 : tmp37589;
  assign tmp37576 = s3 ? tmp37577 : tmp37581;
  assign tmp37597 = l1 ? tmp37193 : tmp36153;
  assign tmp37596 = s0 ? tmp37597 : tmp36456;
  assign tmp37598 = ~(s0 ? tmp37578 : tmp37585);
  assign tmp37595 = s1 ? tmp37596 : tmp37598;
  assign tmp37600 = s0 ? tmp37578 : tmp36115;
  assign tmp37599 = ~(s1 ? tmp37600 : tmp36147);
  assign tmp37594 = s2 ? tmp37595 : tmp37599;
  assign tmp37604 = ~(l1 ? tmp37181 : tmp36466);
  assign tmp37603 = s0 ? tmp37588 : tmp37604;
  assign tmp37605 = s0 ? tmp37122 : tmp37588;
  assign tmp37602 = s1 ? tmp37603 : tmp37605;
  assign tmp37601 = s2 ? tmp36592 : tmp37602;
  assign tmp37593 = ~(s3 ? tmp37594 : tmp37601);
  assign tmp37575 = s4 ? tmp37576 : tmp37593;
  assign tmp37611 = s0 ? tmp37580 : tmp36474;
  assign tmp37612 = ~(l1 ? tmp35724 : tmp35773);
  assign tmp37610 = s1 ? tmp37611 : tmp37612;
  assign tmp37614 = l1 ? tmp37181 : tmp35736;
  assign tmp37616 = l1 ? tmp37181 : tmp36466;
  assign tmp37615 = s0 ? tmp37616 : tmp35775;
  assign tmp37613 = ~(s1 ? tmp37614 : tmp37615);
  assign tmp37609 = s2 ? tmp37610 : tmp37613;
  assign tmp37619 = l1 ? tmp35833 : tmp35806;
  assign tmp37620 = l1 ? tmp35786 : tmp36443;
  assign tmp37618 = s1 ? tmp37619 : tmp37620;
  assign tmp37622 = s0 ? tmp37588 : tmp37122;
  assign tmp37621 = s1 ? tmp37139 : tmp37622;
  assign tmp37617 = s2 ? tmp37618 : tmp37621;
  assign tmp37608 = s3 ? tmp37609 : tmp37617;
  assign tmp37626 = s0 ? tmp35971 : tmp37588;
  assign tmp37625 = s1 ? tmp37626 : tmp36490;
  assign tmp37627 = ~(l1 ? tmp35724 : tmp35736);
  assign tmp37624 = s2 ? tmp37625 : tmp37627;
  assign tmp37631 = l1 ? tmp35833 : tmp36090;
  assign tmp37630 = s0 ? tmp37631 : tmp37308;
  assign tmp37629 = s1 ? tmp37630 : tmp37309;
  assign tmp37628 = s2 ? tmp37629 : tmp35985;
  assign tmp37623 = s3 ? tmp37624 : tmp37628;
  assign tmp37607 = s4 ? tmp37608 : tmp37623;
  assign tmp37636 = s0 ? tmp37620 : tmp35850;
  assign tmp37635 = s1 ? tmp37636 : tmp35879;
  assign tmp37638 = l1 ? tmp35833 : tmp35955;
  assign tmp37637 = s1 ? tmp37638 : tmp36560;
  assign tmp37634 = s2 ? tmp37635 : tmp37637;
  assign tmp37633 = s3 ? tmp37634 : tmp37316;
  assign tmp37641 = s1 ? tmp37324 : tmp35864;
  assign tmp37640 = s2 ? tmp37169 : tmp37641;
  assign tmp37639 = ~(s3 ? tmp37640 : tmp37323);
  assign tmp37632 = s4 ? tmp37633 : tmp37639;
  assign tmp37606 = ~(s5 ? tmp37607 : tmp37632);
  assign tmp37574 = s6 ? tmp37575 : tmp37606;
  assign tmp37573 = s7 ? tmp35709 : tmp37574;
  assign tmp37572 = s8 ? tmp37498 : tmp37573;
  assign tmp37426 = s9 ? tmp37427 : tmp37572;
  assign tmp37649 = l1 ? tmp37181 : tmp35725;
  assign tmp37651 = l1 ? tmp37184 : tmp35719;
  assign tmp37650 = ~(s0 ? tmp36436 : tmp37651);
  assign tmp37648 = s1 ? tmp37649 : tmp37650;
  assign tmp37655 = l1 ? tmp35724 : tmp35768;
  assign tmp37656 = ~(l1 ? tmp37190 : tmp36576);
  assign tmp37654 = s0 ? tmp37655 : tmp37656;
  assign tmp37658 = l1 ? tmp37193 : tmp35914;
  assign tmp37659 = l1 ? tmp37190 : tmp36576;
  assign tmp37657 = ~(s0 ? tmp37658 : tmp37659);
  assign tmp37653 = s1 ? tmp37654 : tmp37657;
  assign tmp37661 = s0 ? tmp37658 : tmp36582;
  assign tmp37663 = ~(l1 ? tmp37181 : tmp35725);
  assign tmp37662 = s0 ? tmp37659 : tmp37663;
  assign tmp37660 = ~(s1 ? tmp37661 : tmp37662);
  assign tmp37652 = s2 ? tmp37653 : tmp37660;
  assign tmp37647 = s3 ? tmp37648 : tmp37652;
  assign tmp37668 = l1 ? tmp37193 : tmp35719;
  assign tmp37667 = s0 ? tmp37668 : tmp36456;
  assign tmp37669 = ~(s0 ? tmp37649 : tmp37656);
  assign tmp37666 = s1 ? tmp37667 : tmp37669;
  assign tmp37671 = s0 ? tmp37649 : tmp36115;
  assign tmp37670 = ~(s1 ? tmp37671 : tmp36147);
  assign tmp37665 = s2 ? tmp37666 : tmp37670;
  assign tmp37675 = ~(l1 ? tmp37181 : tmp36596);
  assign tmp37674 = s0 ? tmp37659 : tmp37675;
  assign tmp37676 = s0 ? tmp37122 : tmp37659;
  assign tmp37673 = s1 ? tmp37674 : tmp37676;
  assign tmp37672 = s2 ? tmp36592 : tmp37673;
  assign tmp37664 = ~(s3 ? tmp37665 : tmp37672);
  assign tmp37646 = s4 ? tmp37647 : tmp37664;
  assign tmp37682 = s0 ? tmp37651 : tmp36474;
  assign tmp37681 = s1 ? tmp37682 : tmp36456;
  assign tmp37684 = l1 ? tmp37181 : 1;
  assign tmp37686 = l1 ? tmp37181 : tmp36596;
  assign tmp37685 = s0 ? tmp37686 : tmp35775;
  assign tmp37683 = ~(s1 ? tmp37684 : tmp37685);
  assign tmp37680 = s2 ? tmp37681 : tmp37683;
  assign tmp37689 = l1 ? tmp35833 : tmp35914;
  assign tmp37688 = s1 ? tmp37689 : tmp37476;
  assign tmp37691 = s0 ? tmp37659 : tmp37372;
  assign tmp37690 = s1 ? tmp37139 : tmp37691;
  assign tmp37687 = s2 ? tmp37688 : tmp37690;
  assign tmp37679 = s3 ? tmp37680 : tmp37687;
  assign tmp37695 = s0 ? tmp35971 : tmp37659;
  assign tmp37694 = s1 ? tmp37695 : tmp36490;
  assign tmp37693 = s2 ? tmp37694 : tmp36490;
  assign tmp37698 = s0 ? tmp37487 : tmp37384;
  assign tmp37697 = s1 ? tmp37698 : tmp37153;
  assign tmp37696 = s2 ? tmp37697 : tmp35985;
  assign tmp37692 = s3 ? tmp37693 : tmp37696;
  assign tmp37678 = s4 ? tmp37679 : tmp37692;
  assign tmp37677 = ~(s5 ? tmp37678 : tmp37488);
  assign tmp37645 = s6 ? tmp37646 : tmp37677;
  assign tmp37644 = s7 ? tmp35709 : tmp37645;
  assign tmp37643 = s8 ? tmp37644 : tmp35709;
  assign tmp37705 = s2 ? tmp37169 : tmp37174;
  assign tmp37704 = ~(s3 ? tmp37705 : tmp37172);
  assign tmp37703 = s4 ? tmp37489 : tmp37704;
  assign tmp37702 = ~(s5 ? tmp37464 : tmp37703);
  assign tmp37701 = s6 ? tmp37430 : tmp37702;
  assign tmp37710 = s2 ? tmp37169 : tmp37324;
  assign tmp37709 = ~(s3 ? tmp37710 : tmp37323);
  assign tmp37708 = s4 ? tmp37633 : tmp37709;
  assign tmp37707 = ~(s5 ? tmp37607 : tmp37708);
  assign tmp37706 = s6 ? tmp37575 : tmp37707;
  assign tmp37700 = s7 ? tmp37701 : tmp37706;
  assign tmp37716 = s2 ? tmp37247 : tmp37571;
  assign tmp37715 = ~(s3 ? tmp37716 : tmp37172);
  assign tmp37714 = s4 ? tmp37562 : tmp37715;
  assign tmp37713 = ~(s5 ? tmp37534 : tmp37714);
  assign tmp37712 = s6 ? tmp37500 : tmp37713;
  assign tmp37718 = ~(s5 ? tmp37678 : tmp37703);
  assign tmp37717 = s6 ? tmp37646 : tmp37718;
  assign tmp37711 = s7 ? tmp37712 : tmp37717;
  assign tmp37699 = s8 ? tmp37700 : tmp37711;
  assign tmp37642 = s9 ? tmp37643 : tmp37699;
  assign tmp37425 = s10 ? tmp37426 : tmp37642;
  assign tmp37722 = s7 ? tmp37429 : tmp37574;
  assign tmp37723 = s7 ? tmp37499 : tmp37645;
  assign tmp37721 = s8 ? tmp37722 : tmp37723;
  assign tmp37720 = s9 ? tmp37643 : tmp37721;
  assign tmp37719 = s10 ? tmp37426 : tmp37720;
  assign tmp37424 = s11 ? tmp37425 : tmp37719;
  assign tmp37085 = s12 ? tmp37086 : tmp37424;
  assign tmp36634 = s13 ? tmp36635 : tmp37085;
  assign tmp35702 = s14 ? tmp35703 : tmp36634;
  assign tmp37736 = ~(s0 ? tmp35852 : tmp35856);
  assign tmp37735 = s1 ? tmp36500 : tmp37736;
  assign tmp37734 = s2 ? tmp37735 : tmp36501;
  assign tmp37733 = s3 ? tmp37734 : tmp36160;
  assign tmp37739 = s0 ? tmp35852 : tmp36167;
  assign tmp37738 = s2 ? tmp36004 : tmp37739;
  assign tmp37737 = ~(s3 ? tmp37738 : tmp36166);
  assign tmp37732 = s4 ? tmp37733 : tmp37737;
  assign tmp37731 = ~(s5 ? tmp36469 : tmp37732);
  assign tmp37730 = s6 ? tmp36614 : tmp37731;
  assign tmp37729 = s7 ? tmp35709 : tmp37730;
  assign tmp37741 = s8 ? tmp37729 : tmp35709;
  assign tmp37744 = s4 ? tmp37733 : tmp36503;
  assign tmp37743 = ~(s5 ? tmp36469 : tmp37744);
  assign tmp37742 = s6 ? tmp36614 : tmp37743;
  assign tmp37740 = s9 ? tmp37741 : tmp37742;
  assign tmp37728 = s10 ? tmp37729 : tmp37740;
  assign tmp37746 = s9 ? tmp37741 : tmp37730;
  assign tmp37745 = s10 ? tmp37729 : tmp37746;
  assign tmp37727 = s11 ? tmp37728 : tmp37745;
  assign tmp37755 = ~(l2 ? tmp35727 : tmp35778);
  assign tmp37754 = l1 ? tmp35904 : tmp37755;
  assign tmp37753 = s1 ? tmp37754 : tmp36435;
  assign tmp37759 = ~(l1 ? tmp36098 : tmp36090);
  assign tmp37758 = s0 ? tmp36441 : tmp37759;
  assign tmp37761 = l1 ? tmp36098 : tmp36090;
  assign tmp37760 = ~(s0 ? tmp36436 : tmp37761);
  assign tmp37757 = s1 ? tmp37758 : tmp37760;
  assign tmp37764 = ~(l1 ? tmp35904 : tmp37755);
  assign tmp37763 = s0 ? tmp37761 : tmp37764;
  assign tmp37762 = ~(s1 ? tmp36618 : tmp37763);
  assign tmp37756 = s2 ? tmp37757 : tmp37762;
  assign tmp37752 = s3 ? tmp37753 : tmp37756;
  assign tmp37768 = ~(s0 ? tmp37754 : tmp37759);
  assign tmp37767 = s1 ? tmp36454 : tmp37768;
  assign tmp37770 = s0 ? tmp37754 : tmp36115;
  assign tmp37769 = ~(s1 ? tmp37770 : tmp36147);
  assign tmp37766 = s2 ? tmp37767 : tmp37769;
  assign tmp37773 = l1 ? tmp35777 : tmp35778;
  assign tmp37772 = s1 ? tmp36436 : tmp37773;
  assign tmp37777 = l2 ? tmp35765 : tmp36091;
  assign tmp37776 = ~(l1 ? tmp35904 : tmp37777);
  assign tmp37775 = s0 ? tmp37761 : tmp37776;
  assign tmp37779 = l1 ? tmp35777 : tmp36153;
  assign tmp37778 = s0 ? tmp37779 : tmp37761;
  assign tmp37774 = s1 ? tmp37775 : tmp37778;
  assign tmp37771 = s2 ? tmp37772 : tmp37774;
  assign tmp37765 = ~(s3 ? tmp37766 : tmp37771);
  assign tmp37751 = s4 ? tmp37752 : tmp37765;
  assign tmp37786 = l1 ? tmp35904 : tmp37777;
  assign tmp37785 = s0 ? tmp37786 : tmp35775;
  assign tmp37784 = ~(s1 ? tmp36477 : tmp37785);
  assign tmp37783 = s2 ? tmp36472 : tmp37784;
  assign tmp37789 = l1 ? tmp35777 : tmp36090;
  assign tmp37788 = s1 ? tmp36482 : tmp37789;
  assign tmp37791 = s0 ? tmp37779 : tmp35811;
  assign tmp37792 = s0 ? tmp37761 : tmp37779;
  assign tmp37790 = s1 ? tmp37791 : tmp37792;
  assign tmp37787 = s2 ? tmp37788 : tmp37790;
  assign tmp37782 = s3 ? tmp37783 : tmp37787;
  assign tmp37797 = l1 ? tmp35821 : tmp35778;
  assign tmp37796 = s0 ? tmp37797 : tmp37761;
  assign tmp37795 = s1 ? tmp37796 : tmp36490;
  assign tmp37794 = s2 ? tmp37795 : tmp36491;
  assign tmp37801 = l1 ? tmp35821 : tmp36153;
  assign tmp37800 = s0 ? tmp36495 : tmp37801;
  assign tmp37803 = l2 ? tmp35765 : tmp35715;
  assign tmp37802 = ~(l1 ? tmp35926 : tmp37803);
  assign tmp37799 = s1 ? tmp37800 : tmp37802;
  assign tmp37805 = s0 ? tmp37773 : tmp35842;
  assign tmp37804 = s1 ? tmp35840 : tmp37805;
  assign tmp37798 = s2 ? tmp37799 : tmp37804;
  assign tmp37793 = s3 ? tmp37794 : tmp37798;
  assign tmp37781 = s4 ? tmp37782 : tmp37793;
  assign tmp37810 = s0 ? tmp37789 : tmp35850;
  assign tmp37809 = s1 ? tmp37810 : tmp35992;
  assign tmp37808 = s2 ? tmp37809 : tmp36501;
  assign tmp37812 = s1 ? tmp35842 : tmp35867;
  assign tmp37813 = s1 ? tmp35812 : tmp36162;
  assign tmp37811 = ~(s2 ? tmp37812 : tmp37813);
  assign tmp37807 = s3 ? tmp37808 : tmp37811;
  assign tmp37817 = ~(l1 ? tmp35777 : tmp36153);
  assign tmp37816 = s1 ? tmp35856 : tmp37817;
  assign tmp37815 = s2 ? tmp37816 : tmp36167;
  assign tmp37819 = l1 ? tmp35857 : tmp35765;
  assign tmp37820 = l1 ? tmp35926 : tmp35714;
  assign tmp37818 = s1 ? tmp37819 : tmp37820;
  assign tmp37814 = ~(s3 ? tmp37815 : tmp37818);
  assign tmp37806 = s4 ? tmp37807 : tmp37814;
  assign tmp37780 = ~(s5 ? tmp37781 : tmp37806);
  assign tmp37750 = s6 ? tmp37751 : tmp37780;
  assign tmp37749 = s7 ? tmp35709 : tmp37750;
  assign tmp37822 = s8 ? tmp37749 : tmp35709;
  assign tmp37828 = s1 ? tmp35840 : tmp37773;
  assign tmp37827 = s2 ? tmp37799 : tmp37828;
  assign tmp37826 = s3 ? tmp37794 : tmp37827;
  assign tmp37825 = s4 ? tmp37782 : tmp37826;
  assign tmp37824 = ~(s5 ? tmp37825 : tmp37806);
  assign tmp37823 = s6 ? tmp37751 : tmp37824;
  assign tmp37821 = s9 ? tmp37822 : tmp37823;
  assign tmp37748 = s10 ? tmp37749 : tmp37821;
  assign tmp37830 = s9 ? tmp37822 : tmp37750;
  assign tmp37829 = s10 ? tmp37749 : tmp37830;
  assign tmp37747 = s11 ? tmp37748 : tmp37829;
  assign tmp37726 = s12 ? tmp37727 : tmp37747;
  assign tmp37842 = ~(l2 ? tmp35765 : tmp35778);
  assign tmp37841 = l1 ? tmp35904 : tmp37842;
  assign tmp37844 = l1 ? tmp35908 : tmp35779;
  assign tmp37843 = ~(s0 ? tmp36652 : tmp37844);
  assign tmp37840 = s1 ? tmp37841 : tmp37843;
  assign tmp37848 = l1 ? tmp35914 : tmp36677;
  assign tmp37850 = ~(l2 ? tmp35727 : tmp36091);
  assign tmp37849 = ~(l1 ? tmp36098 : tmp37850);
  assign tmp37847 = s0 ? tmp37848 : tmp37849;
  assign tmp37852 = l1 ? tmp36098 : tmp37850;
  assign tmp37851 = ~(s0 ? tmp36652 : tmp37852);
  assign tmp37846 = s1 ? tmp37847 : tmp37851;
  assign tmp37854 = s0 ? tmp36652 : tmp36582;
  assign tmp37856 = ~(l1 ? tmp35904 : tmp37842);
  assign tmp37855 = s0 ? tmp37852 : tmp37856;
  assign tmp37853 = ~(s1 ? tmp37854 : tmp37855);
  assign tmp37845 = s2 ? tmp37846 : tmp37853;
  assign tmp37839 = s3 ? tmp37840 : tmp37845;
  assign tmp37861 = l1 ? tmp35768 : tmp35779;
  assign tmp37860 = s0 ? tmp37861 : tmp36456;
  assign tmp37862 = ~(s0 ? tmp37841 : tmp37849);
  assign tmp37859 = s1 ? tmp37860 : tmp37862;
  assign tmp37864 = s0 ? tmp37841 : tmp36115;
  assign tmp37865 = l1 ? tmp35724 : tmp35806;
  assign tmp37863 = ~(s1 ? tmp37864 : tmp37865);
  assign tmp37858 = s2 ? tmp37859 : tmp37863;
  assign tmp37867 = s1 ? tmp36652 : tmp35776;
  assign tmp37871 = l2 ? tmp35727 : tmp36091;
  assign tmp37870 = ~(l1 ? tmp35904 : tmp37871);
  assign tmp37869 = s0 ? tmp37852 : tmp37870;
  assign tmp37872 = s0 ? tmp35776 : tmp37852;
  assign tmp37868 = s1 ? tmp37869 : tmp37872;
  assign tmp37866 = s2 ? tmp37867 : tmp37868;
  assign tmp37857 = ~(s3 ? tmp37858 : tmp37866);
  assign tmp37838 = s4 ? tmp37839 : tmp37857;
  assign tmp37878 = s0 ? tmp37844 : tmp36474;
  assign tmp37877 = s1 ? tmp37878 : tmp36475;
  assign tmp37880 = l1 ? tmp35904 : tmp35914;
  assign tmp37882 = l1 ? tmp35904 : tmp37871;
  assign tmp37881 = s0 ? tmp37882 : tmp35775;
  assign tmp37879 = ~(s1 ? tmp37880 : tmp37881);
  assign tmp37876 = s2 ? tmp37877 : tmp37879;
  assign tmp37885 = l1 ? tmp35777 : tmp37850;
  assign tmp37884 = s1 ? 1 : tmp37885;
  assign tmp37887 = s0 ? tmp35776 : tmp35811;
  assign tmp37888 = s0 ? tmp37852 : tmp35776;
  assign tmp37886 = s1 ? tmp37887 : tmp37888;
  assign tmp37883 = s2 ? tmp37884 : tmp37886;
  assign tmp37875 = s3 ? tmp37876 : tmp37883;
  assign tmp37892 = s0 ? tmp35820 : tmp37852;
  assign tmp37893 = ~(s0 ? tmp36147 : tmp37865);
  assign tmp37891 = s1 ? tmp37892 : tmp37893;
  assign tmp37894 = ~(l2 ? tmp35719 : tmp35724);
  assign tmp37890 = s2 ? tmp37891 : tmp37894;
  assign tmp37898 = l1 ? 1 : tmp37850;
  assign tmp37897 = s0 ? tmp37898 : tmp35820;
  assign tmp37900 = l2 ? tmp35716 : tmp35715;
  assign tmp37899 = ~(l1 ? tmp35926 : tmp37900);
  assign tmp37896 = s1 ? tmp37897 : tmp37899;
  assign tmp37901 = s1 ? tmp35841 : tmp35776;
  assign tmp37895 = s2 ? tmp37896 : tmp37901;
  assign tmp37889 = s3 ? tmp37890 : tmp37895;
  assign tmp37874 = s4 ? tmp37875 : tmp37889;
  assign tmp37906 = s0 ? tmp37885 : tmp35850;
  assign tmp37905 = s1 ? tmp37906 : tmp36901;
  assign tmp37904 = s2 ? tmp37905 : tmp36501;
  assign tmp37909 = l1 ? tmp35812 : tmp35857;
  assign tmp37910 = s0 ? tmp35872 : tmp37076;
  assign tmp37908 = s1 ? tmp37909 : tmp37910;
  assign tmp37907 = ~(s2 ? tmp37812 : tmp37908);
  assign tmp37903 = s3 ? tmp37904 : tmp37907;
  assign tmp37914 = ~(l1 ? tmp35777 : tmp35779);
  assign tmp37913 = s1 ? tmp35856 : tmp37914;
  assign tmp37915 = l1 ? tmp35926 : tmp35914;
  assign tmp37912 = s2 ? tmp37913 : tmp37915;
  assign tmp37917 = s1 ? tmp37819 : tmp35926;
  assign tmp37916 = s2 ? tmp37917 : tmp35872;
  assign tmp37911 = ~(s3 ? tmp37912 : tmp37916);
  assign tmp37902 = s4 ? tmp37903 : tmp37911;
  assign tmp37873 = ~(s5 ? tmp37874 : tmp37902);
  assign tmp37837 = s6 ? tmp37838 : tmp37873;
  assign tmp37836 = s7 ? tmp35709 : tmp37837;
  assign tmp37924 = ~(l2 ? tmp35715 : tmp35778);
  assign tmp37923 = l1 ? tmp35904 : tmp37924;
  assign tmp37922 = s1 ? tmp37923 : tmp37012;
  assign tmp37928 = ~(l1 ? tmp36098 : tmp37064);
  assign tmp37927 = s0 ? tmp36441 : tmp37928;
  assign tmp37930 = l1 ? tmp36098 : tmp37064;
  assign tmp37929 = ~(s0 ? tmp36103 : tmp37930);
  assign tmp37926 = s1 ? tmp37927 : tmp37929;
  assign tmp37933 = ~(l1 ? tmp35904 : tmp37924);
  assign tmp37932 = s0 ? tmp37930 : tmp37933;
  assign tmp37931 = ~(s1 ? tmp37023 : tmp37932);
  assign tmp37925 = s2 ? tmp37926 : tmp37931;
  assign tmp37921 = s3 ? tmp37922 : tmp37925;
  assign tmp37937 = ~(s0 ? tmp37923 : tmp37928);
  assign tmp37936 = s1 ? tmp37029 : tmp37937;
  assign tmp37939 = s0 ? tmp37923 : tmp36115;
  assign tmp37938 = ~(s1 ? tmp37939 : tmp36945);
  assign tmp37935 = s2 ? tmp37936 : tmp37938;
  assign tmp37941 = s1 ? tmp36103 : tmp35776;
  assign tmp37945 = l2 ? tmp35716 : tmp36091;
  assign tmp37944 = ~(l1 ? tmp35904 : tmp37945);
  assign tmp37943 = s0 ? tmp37930 : tmp37944;
  assign tmp37947 = l1 ? tmp35777 : tmp37014;
  assign tmp37946 = s0 ? tmp37947 : tmp37930;
  assign tmp37942 = s1 ? tmp37943 : tmp37946;
  assign tmp37940 = s2 ? tmp37941 : tmp37942;
  assign tmp37934 = ~(s3 ? tmp37935 : tmp37940);
  assign tmp37920 = s4 ? tmp37921 : tmp37934;
  assign tmp37954 = l1 ? tmp35904 : tmp37945;
  assign tmp37953 = s0 ? tmp37954 : tmp35775;
  assign tmp37952 = ~(s1 ? tmp37047 : tmp37953);
  assign tmp37951 = s2 ? tmp37044 : tmp37952;
  assign tmp37957 = l1 ? tmp35777 : tmp37064;
  assign tmp37956 = s1 ? tmp35887 : tmp37957;
  assign tmp37959 = s0 ? tmp37947 : tmp35811;
  assign tmp37960 = s0 ? tmp37930 : tmp37947;
  assign tmp37958 = s1 ? tmp37959 : tmp37960;
  assign tmp37955 = s2 ? tmp37956 : tmp37958;
  assign tmp37950 = s3 ? tmp37951 : tmp37955;
  assign tmp37964 = s0 ? tmp35820 : tmp37930;
  assign tmp37963 = s1 ? tmp37964 : tmp36977;
  assign tmp37962 = s2 ? tmp37963 : tmp37059;
  assign tmp37968 = l1 ? tmp35821 : tmp37014;
  assign tmp37967 = s0 ? tmp37063 : tmp37968;
  assign tmp37966 = s1 ? tmp37967 : tmp37899;
  assign tmp37965 = s2 ? tmp37966 : tmp37901;
  assign tmp37961 = s3 ? tmp37962 : tmp37965;
  assign tmp37949 = s4 ? tmp37950 : tmp37961;
  assign tmp37973 = s0 ? tmp37957 : tmp35850;
  assign tmp37972 = s1 ? tmp37973 : tmp36991;
  assign tmp37971 = s2 ? tmp37972 : tmp36501;
  assign tmp37970 = s3 ? tmp37971 : tmp37907;
  assign tmp37977 = ~(l1 ? tmp35777 : tmp37014);
  assign tmp37976 = s1 ? tmp35856 : tmp37977;
  assign tmp37975 = s2 ? tmp37976 : tmp37079;
  assign tmp37974 = ~(s3 ? tmp37975 : tmp37916);
  assign tmp37969 = s4 ? tmp37970 : tmp37974;
  assign tmp37948 = ~(s5 ? tmp37949 : tmp37969);
  assign tmp37919 = s6 ? tmp37920 : tmp37948;
  assign tmp37918 = s7 ? tmp35709 : tmp37919;
  assign tmp37835 = s8 ? tmp37836 : tmp37918;
  assign tmp37985 = ~(l2 ? tmp35715 : tmp35719);
  assign tmp37984 = l1 ? tmp35904 : tmp37985;
  assign tmp37983 = s1 ? tmp37984 : tmp36922;
  assign tmp37989 = ~(l1 ? tmp36098 : tmp36983);
  assign tmp37988 = s0 ? tmp36441 : tmp37989;
  assign tmp37991 = l1 ? tmp36098 : tmp36983;
  assign tmp37990 = ~(s0 ? tmp36103 : tmp37991);
  assign tmp37987 = s1 ? tmp37988 : tmp37990;
  assign tmp37994 = ~(l1 ? tmp35904 : tmp37985);
  assign tmp37993 = s0 ? tmp37991 : tmp37994;
  assign tmp37992 = ~(s1 ? tmp37023 : tmp37993);
  assign tmp37986 = s2 ? tmp37987 : tmp37992;
  assign tmp37982 = s3 ? tmp37983 : tmp37986;
  assign tmp37998 = ~(s0 ? tmp37984 : tmp37989);
  assign tmp37997 = s1 ? tmp36940 : tmp37998;
  assign tmp38000 = s0 ? tmp37984 : tmp36115;
  assign tmp37999 = ~(s1 ? tmp38000 : tmp36945);
  assign tmp37996 = s2 ? tmp37997 : tmp37999;
  assign tmp38005 = l2 ? tmp35716 : tmp35720;
  assign tmp38004 = ~(l1 ? tmp35904 : tmp38005);
  assign tmp38003 = s0 ? tmp37991 : tmp38004;
  assign tmp38006 = s0 ? tmp37947 : tmp37991;
  assign tmp38002 = s1 ? tmp38003 : tmp38006;
  assign tmp38001 = s2 ? tmp37941 : tmp38002;
  assign tmp37995 = ~(s3 ? tmp37996 : tmp38001);
  assign tmp37981 = s4 ? tmp37982 : tmp37995;
  assign tmp38011 = s1 ? tmp36960 : tmp36475;
  assign tmp38014 = l1 ? tmp35904 : tmp38005;
  assign tmp38013 = s0 ? tmp38014 : tmp35775;
  assign tmp38012 = ~(s1 ? tmp36962 : tmp38013);
  assign tmp38010 = s2 ? tmp38011 : tmp38012;
  assign tmp38017 = l1 ? tmp35777 : tmp36983;
  assign tmp38016 = s1 ? tmp35887 : tmp38017;
  assign tmp38020 = l1 ? tmp35777 : tmp36924;
  assign tmp38019 = s0 ? tmp37991 : tmp38020;
  assign tmp38018 = s1 ? tmp37959 : tmp38019;
  assign tmp38015 = s2 ? tmp38016 : tmp38018;
  assign tmp38009 = s3 ? tmp38010 : tmp38015;
  assign tmp38024 = s0 ? tmp35820 : tmp37991;
  assign tmp38023 = s1 ? tmp38024 : tmp36977;
  assign tmp38022 = s2 ? tmp38023 : tmp36978;
  assign tmp38028 = l1 ? tmp35821 : tmp36924;
  assign tmp38027 = s0 ? tmp36982 : tmp38028;
  assign tmp38029 = ~(l1 ? tmp35926 : tmp35838);
  assign tmp38026 = s1 ? tmp38027 : tmp38029;
  assign tmp38025 = s2 ? tmp38026 : tmp37901;
  assign tmp38021 = s3 ? tmp38022 : tmp38025;
  assign tmp38008 = s4 ? tmp38009 : tmp38021;
  assign tmp38034 = s0 ? tmp38017 : tmp35850;
  assign tmp38033 = s1 ? tmp38034 : tmp36991;
  assign tmp38032 = s2 ? tmp38033 : tmp36501;
  assign tmp38037 = s0 ? tmp35872 : tmp36907;
  assign tmp38036 = s1 ? tmp37909 : tmp38037;
  assign tmp38035 = ~(s2 ? tmp37812 : tmp38036);
  assign tmp38031 = s3 ? tmp38032 : tmp38035;
  assign tmp38039 = s2 ? tmp37976 : tmp36914;
  assign tmp38042 = l1 ? tmp35926 : tmp35857;
  assign tmp38041 = s1 ? tmp37819 : tmp38042;
  assign tmp38040 = s2 ? tmp38041 : tmp35872;
  assign tmp38038 = ~(s3 ? tmp38039 : tmp38040);
  assign tmp38030 = s4 ? tmp38031 : tmp38038;
  assign tmp38007 = ~(s5 ? tmp38008 : tmp38030);
  assign tmp37980 = s6 ? tmp37981 : tmp38007;
  assign tmp37979 = s7 ? tmp35709 : tmp37980;
  assign tmp37978 = s8 ? tmp37918 : tmp37979;
  assign tmp37834 = s9 ? tmp37835 : tmp37978;
  assign tmp38044 = s8 ? tmp37918 : tmp35709;
  assign tmp38050 = ~(s3 ? tmp37912 : tmp37917);
  assign tmp38049 = s4 ? tmp37903 : tmp38050;
  assign tmp38048 = ~(s5 ? tmp37874 : tmp38049);
  assign tmp38047 = s6 ? tmp37838 : tmp38048;
  assign tmp38054 = ~(s3 ? tmp38039 : tmp38041);
  assign tmp38053 = s4 ? tmp38031 : tmp38054;
  assign tmp38052 = ~(s5 ? tmp38008 : tmp38053);
  assign tmp38051 = s6 ? tmp37981 : tmp38052;
  assign tmp38046 = s7 ? tmp38047 : tmp38051;
  assign tmp38058 = ~(s3 ? tmp37975 : tmp37917);
  assign tmp38057 = s4 ? tmp37970 : tmp38058;
  assign tmp38056 = ~(s5 ? tmp37949 : tmp38057);
  assign tmp38055 = s6 ? tmp37920 : tmp38056;
  assign tmp38045 = s8 ? tmp38046 : tmp38055;
  assign tmp38043 = s9 ? tmp38044 : tmp38045;
  assign tmp37833 = s10 ? tmp37834 : tmp38043;
  assign tmp38062 = s7 ? tmp37837 : tmp37980;
  assign tmp38061 = s8 ? tmp38062 : tmp37919;
  assign tmp38060 = s9 ? tmp38044 : tmp38061;
  assign tmp38059 = s10 ? tmp37834 : tmp38060;
  assign tmp37832 = s11 ? tmp37833 : tmp38059;
  assign tmp38071 = s1 ? tmp35841 : tmp37773;
  assign tmp38070 = s2 ? tmp37799 : tmp38071;
  assign tmp38069 = s3 ? tmp37794 : tmp38070;
  assign tmp38068 = s4 ? tmp37782 : tmp38069;
  assign tmp38077 = ~(l2 ? 1 : tmp35765);
  assign tmp38076 = s0 ? tmp35842 : tmp38077;
  assign tmp38075 = ~(s1 ? tmp38076 : tmp36732);
  assign tmp38074 = ~(s2 ? tmp37812 : tmp38075);
  assign tmp38073 = s3 ? tmp37808 : tmp38074;
  assign tmp38081 = ~(l1 ? tmp35926 : tmp35714);
  assign tmp38080 = ~(s0 ? tmp35842 : tmp38081);
  assign tmp38079 = s1 ? tmp37819 : tmp38080;
  assign tmp38078 = ~(s3 ? tmp37815 : tmp38079);
  assign tmp38072 = s4 ? tmp38073 : tmp38078;
  assign tmp38067 = ~(s5 ? tmp38068 : tmp38072);
  assign tmp38066 = s6 ? tmp37751 : tmp38067;
  assign tmp38065 = s7 ? tmp35709 : tmp38066;
  assign tmp38083 = s8 ? tmp38065 : tmp35709;
  assign tmp38086 = s4 ? tmp38073 : tmp37814;
  assign tmp38085 = ~(s5 ? tmp38068 : tmp38086);
  assign tmp38084 = s6 ? tmp37751 : tmp38085;
  assign tmp38082 = s9 ? tmp38083 : tmp38084;
  assign tmp38064 = s10 ? tmp38065 : tmp38082;
  assign tmp38088 = s9 ? tmp38083 : tmp38066;
  assign tmp38087 = s10 ? tmp38065 : tmp38088;
  assign tmp38063 = s11 ? tmp38064 : tmp38087;
  assign tmp37831 = s12 ? tmp37832 : tmp38063;
  assign tmp37725 = s13 ? tmp37726 : tmp37831;
  assign tmp38100 = l1 ? tmp35714 : tmp36827;
  assign tmp38102 = l1 ? tmp35729 : tmp35740;
  assign tmp38101 = ~(s0 ? tmp35749 : tmp38102);
  assign tmp38099 = s1 ? tmp38100 : tmp38101;
  assign tmp38106 = ~(l1 ? tmp35739 : tmp36835);
  assign tmp38105 = s0 ? tmp37439 : tmp38106;
  assign tmp38108 = l1 ? tmp35743 : tmp35736;
  assign tmp38109 = l1 ? tmp35739 : tmp36835;
  assign tmp38107 = ~(s0 ? tmp38108 : tmp38109);
  assign tmp38104 = s1 ? tmp38105 : tmp38107;
  assign tmp38111 = s0 ? tmp38108 : tmp36582;
  assign tmp38113 = ~(l1 ? tmp35714 : tmp36827);
  assign tmp38112 = s0 ? tmp38109 : tmp38113;
  assign tmp38110 = ~(s1 ? tmp38111 : tmp38112);
  assign tmp38103 = s2 ? tmp38104 : tmp38110;
  assign tmp38098 = s3 ? tmp38099 : tmp38103;
  assign tmp38118 = l1 ? tmp35743 : tmp35740;
  assign tmp38117 = s0 ? tmp38118 : tmp36530;
  assign tmp38119 = ~(s0 ? tmp38100 : tmp38106);
  assign tmp38116 = s1 ? tmp38117 : tmp38119;
  assign tmp38121 = s0 ? tmp38100 : tmp36115;
  assign tmp38120 = ~(s1 ? tmp38121 : tmp35824);
  assign tmp38115 = s2 ? tmp38116 : tmp38120;
  assign tmp38125 = ~(l1 ? tmp35714 : tmp36858);
  assign tmp38124 = s0 ? tmp38109 : tmp38125;
  assign tmp38127 = l1 ? tmp35786 : tmp36854;
  assign tmp38126 = s0 ? tmp38127 : tmp38109;
  assign tmp38123 = s1 ? tmp38124 : tmp38126;
  assign tmp38122 = s2 ? tmp36852 : tmp38123;
  assign tmp38114 = ~(s3 ? tmp38115 : tmp38122);
  assign tmp38097 = s4 ? tmp38098 : tmp38114;
  assign tmp38133 = s0 ? tmp38102 : tmp36474;
  assign tmp38132 = s1 ? tmp38133 : tmp37469;
  assign tmp38135 = l1 ? tmp35714 : tmp35806;
  assign tmp38137 = l1 ? tmp35714 : tmp36858;
  assign tmp38136 = s0 ? tmp38137 : tmp35775;
  assign tmp38134 = ~(s1 ? tmp38135 : tmp38136);
  assign tmp38131 = s2 ? tmp38132 : tmp38134;
  assign tmp38140 = l1 ? tmp35806 : tmp35736;
  assign tmp38141 = l1 ? tmp35786 : tmp36835;
  assign tmp38139 = s1 ? tmp38140 : tmp38141;
  assign tmp38143 = s0 ? tmp38127 : tmp35850;
  assign tmp38145 = l1 ? tmp35815 : tmp36878;
  assign tmp38144 = s0 ? tmp38109 : tmp38145;
  assign tmp38142 = s1 ? tmp38143 : tmp38144;
  assign tmp38138 = s2 ? tmp38139 : tmp38142;
  assign tmp38130 = s3 ? tmp38131 : tmp38138;
  assign tmp38149 = s0 ? tmp36883 : tmp38109;
  assign tmp38148 = s1 ? tmp38149 : tmp36884;
  assign tmp38150 = ~(s1 ? tmp35827 : tmp35824);
  assign tmp38147 = s2 ? tmp38148 : tmp38150;
  assign tmp38154 = l1 ? tmp35833 : tmp35731;
  assign tmp38155 = l1 ? tmp35835 : tmp36878;
  assign tmp38153 = s0 ? tmp38154 : tmp38155;
  assign tmp38157 = l1 ? tmp35714 : tmp36894;
  assign tmp38156 = ~(s0 ? tmp35827 : tmp38157);
  assign tmp38152 = s1 ? tmp38153 : tmp38156;
  assign tmp38151 = s2 ? tmp38152 : tmp36895;
  assign tmp38146 = s3 ? tmp38147 : tmp38151;
  assign tmp38129 = s4 ? tmp38130 : tmp38146;
  assign tmp38162 = s0 ? tmp38141 : tmp35850;
  assign tmp38163 = ~(l1 ? tmp35812 : tmp35806);
  assign tmp38161 = s1 ? tmp38162 : tmp38163;
  assign tmp38160 = s2 ? tmp38161 : tmp37493;
  assign tmp38165 = s1 ? tmp36906 : tmp35873;
  assign tmp38164 = ~(s2 ? tmp37163 : tmp38165);
  assign tmp38159 = s3 ? tmp38160 : tmp38164;
  assign tmp38168 = s1 ? tmp35877 : tmp38127;
  assign tmp38169 = ~(s1 ? tmp38135 : tmp35864);
  assign tmp38167 = s2 ? tmp38168 : tmp38169;
  assign tmp38172 = l1 ? tmp35714 : tmp35833;
  assign tmp38171 = s1 ? tmp37173 : tmp38172;
  assign tmp38170 = ~(s2 ? tmp38171 : tmp35897);
  assign tmp38166 = s3 ? tmp38167 : tmp38170;
  assign tmp38158 = s4 ? tmp38159 : tmp38166;
  assign tmp38128 = ~(s5 ? tmp38129 : tmp38158);
  assign tmp38096 = s6 ? tmp38097 : tmp38128;
  assign tmp38095 = s7 ? tmp35709 : tmp38096;
  assign tmp38178 = l1 ? tmp37181 : tmp36827;
  assign tmp38180 = l1 ? tmp37184 : tmp35740;
  assign tmp38179 = ~(s0 ? tmp36652 : tmp38180);
  assign tmp38177 = s1 ? tmp38178 : tmp38179;
  assign tmp38184 = ~(l1 ? tmp37190 : tmp36835);
  assign tmp38183 = s0 ? tmp37510 : tmp38184;
  assign tmp38186 = l1 ? tmp37193 : tmp35736;
  assign tmp38187 = l1 ? tmp37190 : tmp36835;
  assign tmp38185 = ~(s0 ? tmp38186 : tmp38187);
  assign tmp38182 = s1 ? tmp38183 : tmp38185;
  assign tmp38189 = s0 ? tmp38186 : tmp35795;
  assign tmp38191 = ~(l1 ? tmp37181 : tmp36827);
  assign tmp38190 = s0 ? tmp38187 : tmp38191;
  assign tmp38188 = ~(s1 ? tmp38189 : tmp38190);
  assign tmp38181 = s2 ? tmp38182 : tmp38188;
  assign tmp38176 = s3 ? tmp38177 : tmp38181;
  assign tmp38196 = l1 ? tmp37193 : tmp35740;
  assign tmp38195 = s0 ? tmp38196 : tmp36456;
  assign tmp38197 = ~(s0 ? tmp38178 : tmp38184);
  assign tmp38194 = s1 ? tmp38195 : tmp38197;
  assign tmp38199 = s0 ? tmp38178 : tmp36115;
  assign tmp38198 = ~(s1 ? tmp38199 : tmp37865);
  assign tmp38193 = s2 ? tmp38194 : tmp38198;
  assign tmp38201 = s1 ? tmp36652 : tmp36853;
  assign tmp38204 = ~(l1 ? tmp37181 : tmp36858);
  assign tmp38203 = s0 ? tmp38187 : tmp38204;
  assign tmp38205 = s0 ? tmp38127 : tmp38187;
  assign tmp38202 = s1 ? tmp38203 : tmp38205;
  assign tmp38200 = s2 ? tmp38201 : tmp38202;
  assign tmp38192 = ~(s3 ? tmp38193 : tmp38200);
  assign tmp38175 = s4 ? tmp38176 : tmp38192;
  assign tmp38211 = s0 ? tmp38180 : tmp36474;
  assign tmp38210 = s1 ? tmp38211 : tmp37539;
  assign tmp38213 = l1 ? tmp37181 : tmp35806;
  assign tmp38215 = l1 ? tmp37181 : tmp36858;
  assign tmp38214 = s0 ? tmp38215 : tmp37544;
  assign tmp38212 = ~(s1 ? tmp38213 : tmp38214);
  assign tmp38209 = s2 ? tmp38210 : tmp38212;
  assign tmp38217 = s1 ? tmp37160 : tmp38141;
  assign tmp38220 = l1 ? tmp35786 : tmp36878;
  assign tmp38219 = s0 ? tmp38187 : tmp38220;
  assign tmp38218 = s1 ? tmp38143 : tmp38219;
  assign tmp38216 = s2 ? tmp38217 : tmp38218;
  assign tmp38208 = s3 ? tmp38209 : tmp38216;
  assign tmp38224 = s0 ? tmp36883 : tmp38187;
  assign tmp38223 = s1 ? tmp38224 : tmp37893;
  assign tmp38225 = ~(l1 ? tmp35724 : tmp35806);
  assign tmp38222 = s2 ? tmp38223 : tmp38225;
  assign tmp38229 = l1 ? tmp36894 : tmp36878;
  assign tmp38228 = s0 ? tmp38154 : tmp38229;
  assign tmp38230 = ~(l1 ? tmp35714 : tmp36894);
  assign tmp38227 = s1 ? tmp38228 : tmp38230;
  assign tmp38226 = s2 ? tmp38227 : tmp36895;
  assign tmp38221 = s3 ? tmp38222 : tmp38226;
  assign tmp38207 = s4 ? tmp38208 : tmp38221;
  assign tmp38233 = s2 ? tmp38161 : tmp37566;
  assign tmp38232 = s3 ? tmp38233 : tmp38164;
  assign tmp38231 = s4 ? tmp38232 : tmp38166;
  assign tmp38206 = ~(s5 ? tmp38207 : tmp38231);
  assign tmp38174 = s6 ? tmp38175 : tmp38206;
  assign tmp38173 = s7 ? tmp35709 : tmp38174;
  assign tmp38094 = s8 ? tmp38095 : tmp38173;
  assign tmp38240 = l1 ? tmp37181 : tmp36921;
  assign tmp38242 = l1 ? tmp37184 : tmp36924;
  assign tmp38241 = ~(s0 ? tmp36103 : tmp38242);
  assign tmp38239 = s1 ? tmp38240 : tmp38241;
  assign tmp38246 = ~(l1 ? tmp37190 : tmp36929);
  assign tmp38245 = s0 ? tmp37584 : tmp38246;
  assign tmp38248 = l1 ? tmp37193 : tmp35767;
  assign tmp38249 = l1 ? tmp37190 : tmp36929;
  assign tmp38247 = ~(s0 ? tmp38248 : tmp38249);
  assign tmp38244 = s1 ? tmp38245 : tmp38247;
  assign tmp38251 = s0 ? tmp38248 : tmp36582;
  assign tmp38253 = ~(l1 ? tmp37181 : tmp36921);
  assign tmp38252 = s0 ? tmp38249 : tmp38253;
  assign tmp38250 = ~(s1 ? tmp38251 : tmp38252);
  assign tmp38243 = s2 ? tmp38244 : tmp38250;
  assign tmp38238 = s3 ? tmp38239 : tmp38243;
  assign tmp38258 = l1 ? tmp37193 : tmp36924;
  assign tmp38257 = s0 ? tmp38258 : tmp36456;
  assign tmp38259 = ~(s0 ? tmp38240 : tmp38246);
  assign tmp38256 = s1 ? tmp38257 : tmp38259;
  assign tmp38261 = s0 ? tmp38240 : tmp36115;
  assign tmp38260 = ~(s1 ? tmp38261 : tmp36945);
  assign tmp38255 = s2 ? tmp38256 : tmp38260;
  assign tmp38265 = ~(l1 ? tmp37181 : tmp36951);
  assign tmp38264 = s0 ? tmp38249 : tmp38265;
  assign tmp38267 = l1 ? tmp35786 : tmp36954;
  assign tmp38266 = s0 ? tmp38267 : tmp38249;
  assign tmp38263 = s1 ? tmp38264 : tmp38266;
  assign tmp38262 = s2 ? tmp36947 : tmp38263;
  assign tmp38254 = ~(s3 ? tmp38255 : tmp38262);
  assign tmp38237 = s4 ? tmp38238 : tmp38254;
  assign tmp38273 = s0 ? tmp38242 : tmp36474;
  assign tmp38272 = s1 ? tmp38273 : tmp37612;
  assign tmp38275 = l1 ? tmp37181 : tmp35833;
  assign tmp38277 = l1 ? tmp37181 : tmp36951;
  assign tmp38276 = s0 ? tmp38277 : tmp35775;
  assign tmp38274 = ~(s1 ? tmp38275 : tmp38276);
  assign tmp38271 = s2 ? tmp38272 : tmp38274;
  assign tmp38280 = l1 ? tmp35786 : tmp36929;
  assign tmp38279 = s1 ? tmp37315 : tmp38280;
  assign tmp38282 = s0 ? tmp38267 : tmp35850;
  assign tmp38284 = l1 ? tmp35786 : tmp36972;
  assign tmp38283 = s0 ? tmp38249 : tmp38284;
  assign tmp38281 = s1 ? tmp38282 : tmp38283;
  assign tmp38278 = s2 ? tmp38279 : tmp38281;
  assign tmp38270 = s3 ? tmp38271 : tmp38278;
  assign tmp38288 = s0 ? tmp36883 : tmp38249;
  assign tmp38287 = s1 ? tmp38288 : tmp36977;
  assign tmp38289 = ~(l1 ? tmp35724 : tmp35833);
  assign tmp38286 = s2 ? tmp38287 : tmp38289;
  assign tmp38293 = l1 ? tmp35833 : tmp36983;
  assign tmp38294 = l1 ? tmp36894 : tmp36972;
  assign tmp38292 = s0 ? tmp38293 : tmp38294;
  assign tmp38291 = s1 ? tmp38292 : tmp38230;
  assign tmp38290 = s2 ? tmp38291 : tmp36895;
  assign tmp38285 = s3 ? tmp38286 : tmp38290;
  assign tmp38269 = s4 ? tmp38270 : tmp38285;
  assign tmp38299 = s0 ? tmp38280 : tmp35850;
  assign tmp38300 = ~(l1 ? tmp35812 : tmp35833);
  assign tmp38298 = s1 ? tmp38299 : tmp38300;
  assign tmp38297 = s2 ? tmp38298 : tmp37637;
  assign tmp38296 = s3 ? tmp38297 : tmp38164;
  assign tmp38303 = s1 ? tmp35877 : tmp38267;
  assign tmp38304 = ~(s1 ? tmp38172 : tmp35864);
  assign tmp38302 = s2 ? tmp38303 : tmp38304;
  assign tmp38301 = s3 ? tmp38302 : tmp38170;
  assign tmp38295 = s4 ? tmp38296 : tmp38301;
  assign tmp38268 = ~(s5 ? tmp38269 : tmp38295);
  assign tmp38236 = s6 ? tmp38237 : tmp38268;
  assign tmp38235 = s7 ? tmp35709 : tmp38236;
  assign tmp38234 = s8 ? tmp38173 : tmp38235;
  assign tmp38093 = s9 ? tmp38094 : tmp38234;
  assign tmp38313 = s0 ? tmp37655 : tmp38246;
  assign tmp38315 = l1 ? tmp37193 : tmp35724;
  assign tmp38314 = ~(s0 ? tmp38315 : tmp38249);
  assign tmp38312 = s1 ? tmp38313 : tmp38314;
  assign tmp38317 = s0 ? tmp38315 : tmp36582;
  assign tmp38316 = ~(s1 ? tmp38317 : tmp38252);
  assign tmp38311 = s2 ? tmp38312 : tmp38316;
  assign tmp38310 = s3 ? tmp38239 : tmp38311;
  assign tmp38309 = s4 ? tmp38310 : tmp38254;
  assign tmp38322 = s1 ? tmp38273 : tmp36456;
  assign tmp38321 = s2 ? tmp38322 : tmp38274;
  assign tmp38324 = s1 ? tmp37391 : tmp38280;
  assign tmp38323 = s2 ? tmp38324 : tmp38281;
  assign tmp38320 = s3 ? tmp38321 : tmp38323;
  assign tmp38319 = s4 ? tmp38320 : tmp38285;
  assign tmp38327 = s2 ? tmp38298 : tmp37493;
  assign tmp38326 = s3 ? tmp38327 : tmp38164;
  assign tmp38325 = s4 ? tmp38326 : tmp38301;
  assign tmp38318 = ~(s5 ? tmp38319 : tmp38325);
  assign tmp38308 = s6 ? tmp38309 : tmp38318;
  assign tmp38307 = s7 ? tmp35709 : tmp38308;
  assign tmp38306 = s8 ? tmp38307 : tmp35709;
  assign tmp38335 = s1 ? tmp38153 : tmp38230;
  assign tmp38334 = s2 ? tmp38335 : tmp36895;
  assign tmp38333 = s3 ? tmp38147 : tmp38334;
  assign tmp38332 = s4 ? tmp38130 : tmp38333;
  assign tmp38339 = ~(l1 ? tmp35714 : tmp35806);
  assign tmp38338 = s2 ? tmp38168 : tmp38339;
  assign tmp38340 = ~(s1 ? tmp37173 : tmp38172);
  assign tmp38337 = s3 ? tmp38338 : tmp38340;
  assign tmp38336 = s4 ? tmp38159 : tmp38337;
  assign tmp38331 = ~(s5 ? tmp38332 : tmp38336);
  assign tmp38330 = s6 ? tmp38097 : tmp38331;
  assign tmp38346 = ~(l1 ? tmp35714 : tmp35833);
  assign tmp38345 = s2 ? tmp38303 : tmp38346;
  assign tmp38344 = s3 ? tmp38345 : tmp38340;
  assign tmp38343 = s4 ? tmp38296 : tmp38344;
  assign tmp38342 = ~(s5 ? tmp38269 : tmp38343);
  assign tmp38341 = s6 ? tmp38237 : tmp38342;
  assign tmp38329 = s7 ? tmp38330 : tmp38341;
  assign tmp38350 = s4 ? tmp38232 : tmp38337;
  assign tmp38349 = ~(s5 ? tmp38207 : tmp38350);
  assign tmp38348 = s6 ? tmp38175 : tmp38349;
  assign tmp38353 = s4 ? tmp38326 : tmp38344;
  assign tmp38352 = ~(s5 ? tmp38319 : tmp38353);
  assign tmp38351 = s6 ? tmp38309 : tmp38352;
  assign tmp38347 = s7 ? tmp38348 : tmp38351;
  assign tmp38328 = s8 ? tmp38329 : tmp38347;
  assign tmp38305 = s9 ? tmp38306 : tmp38328;
  assign tmp38092 = s10 ? tmp38093 : tmp38305;
  assign tmp38357 = s7 ? tmp38096 : tmp38236;
  assign tmp38358 = s7 ? tmp38174 : tmp38308;
  assign tmp38356 = s8 ? tmp38357 : tmp38358;
  assign tmp38355 = s9 ? tmp38306 : tmp38356;
  assign tmp38354 = s10 ? tmp38093 : tmp38355;
  assign tmp38091 = s11 ? tmp38092 : tmp38354;
  assign tmp38368 = ~(s0 ? tmp36652 : tmp38102);
  assign tmp38367 = s1 ? tmp38100 : tmp38368;
  assign tmp38366 = s3 ? tmp38367 : tmp38103;
  assign tmp38372 = s0 ? tmp38118 : tmp36456;
  assign tmp38371 = s1 ? tmp38372 : tmp38119;
  assign tmp38373 = ~(s1 ? tmp38121 : tmp37865);
  assign tmp38370 = s2 ? tmp38371 : tmp38373;
  assign tmp38374 = s2 ? tmp38201 : tmp38123;
  assign tmp38369 = ~(s3 ? tmp38370 : tmp38374);
  assign tmp38365 = s4 ? tmp38366 : tmp38369;
  assign tmp38379 = s1 ? tmp38149 : tmp37893;
  assign tmp38380 = ~(l1 ? tmp35736 : tmp35806);
  assign tmp38378 = s2 ? tmp38379 : tmp38380;
  assign tmp38377 = s3 ? tmp38378 : tmp38334;
  assign tmp38376 = s4 ? tmp38130 : tmp38377;
  assign tmp38386 = ~(l1 ? tmp35833 : tmp36713);
  assign tmp38385 = s0 ? tmp35856 : tmp38386;
  assign tmp38384 = ~(s1 ? tmp38385 : tmp35827);
  assign tmp38383 = s2 ? tmp38161 : tmp38384;
  assign tmp38387 = ~(s2 ? tmp35997 : tmp38165);
  assign tmp38382 = s3 ? tmp38383 : tmp38387;
  assign tmp38391 = ~(l1 ? tmp35786 : tmp36854);
  assign tmp38390 = s1 ? tmp36000 : tmp38391;
  assign tmp38389 = s2 ? tmp38390 : tmp38135;
  assign tmp38393 = s0 ? tmp35856 : tmp37173;
  assign tmp38392 = s1 ? tmp38393 : tmp38172;
  assign tmp38388 = ~(s3 ? tmp38389 : tmp38392);
  assign tmp38381 = s4 ? tmp38382 : tmp38388;
  assign tmp38375 = ~(s5 ? tmp38376 : tmp38381);
  assign tmp38364 = s6 ? tmp38365 : tmp38375;
  assign tmp38363 = s7 ? tmp35709 : tmp38364;
  assign tmp38398 = s3 ? tmp38233 : tmp38387;
  assign tmp38399 = ~(s3 ? tmp38389 : tmp38171);
  assign tmp38397 = s4 ? tmp38398 : tmp38399;
  assign tmp38396 = ~(s5 ? tmp38207 : tmp38397);
  assign tmp38395 = s6 ? tmp38175 : tmp38396;
  assign tmp38394 = s7 ? tmp35709 : tmp38395;
  assign tmp38362 = s8 ? tmp38363 : tmp38394;
  assign tmp38406 = l1 ? tmp37181 : tmp37011;
  assign tmp38408 = l1 ? tmp37184 : tmp37014;
  assign tmp38407 = ~(s0 ? tmp36103 : tmp38408);
  assign tmp38405 = s1 ? tmp38406 : tmp38407;
  assign tmp38412 = ~(l1 ? tmp37190 : tmp37019);
  assign tmp38411 = s0 ? tmp37584 : tmp38412;
  assign tmp38414 = l1 ? tmp37190 : tmp37019;
  assign tmp38413 = ~(s0 ? tmp38248 : tmp38414);
  assign tmp38410 = s1 ? tmp38411 : tmp38413;
  assign tmp38417 = ~(l1 ? tmp37181 : tmp37011);
  assign tmp38416 = s0 ? tmp38414 : tmp38417;
  assign tmp38415 = ~(s1 ? tmp38251 : tmp38416);
  assign tmp38409 = s2 ? tmp38410 : tmp38415;
  assign tmp38404 = s3 ? tmp38405 : tmp38409;
  assign tmp38422 = l1 ? tmp37193 : tmp37014;
  assign tmp38421 = s0 ? tmp38422 : tmp36456;
  assign tmp38423 = ~(s0 ? tmp38406 : tmp38412);
  assign tmp38420 = s1 ? tmp38421 : tmp38423;
  assign tmp38425 = s0 ? tmp38406 : tmp36115;
  assign tmp38424 = ~(s1 ? tmp38425 : tmp36945);
  assign tmp38419 = s2 ? tmp38420 : tmp38424;
  assign tmp38429 = ~(l1 ? tmp37181 : tmp37038);
  assign tmp38428 = s0 ? tmp38414 : tmp38429;
  assign tmp38430 = s0 ? tmp38267 : tmp38414;
  assign tmp38427 = s1 ? tmp38428 : tmp38430;
  assign tmp38426 = s2 ? tmp36947 : tmp38427;
  assign tmp38418 = ~(s3 ? tmp38419 : tmp38426);
  assign tmp38403 = s4 ? tmp38404 : tmp38418;
  assign tmp38436 = s0 ? tmp38408 : tmp36474;
  assign tmp38435 = s1 ? tmp38436 : tmp37612;
  assign tmp38438 = l1 ? tmp37181 : tmp35865;
  assign tmp38440 = l1 ? tmp37181 : tmp37038;
  assign tmp38439 = s0 ? tmp38440 : tmp35775;
  assign tmp38437 = ~(s1 ? tmp38438 : tmp38439);
  assign tmp38434 = s2 ? tmp38435 : tmp38437;
  assign tmp38443 = l1 ? tmp35786 : tmp37019;
  assign tmp38442 = s1 ? tmp37315 : tmp38443;
  assign tmp38445 = s0 ? tmp38414 : tmp38267;
  assign tmp38444 = s1 ? tmp38282 : tmp38445;
  assign tmp38441 = s2 ? tmp38442 : tmp38444;
  assign tmp38433 = s3 ? tmp38434 : tmp38441;
  assign tmp38449 = s0 ? tmp36883 : tmp38414;
  assign tmp38448 = s1 ? tmp38449 : tmp36977;
  assign tmp38450 = ~(l1 ? tmp35724 : tmp35865);
  assign tmp38447 = s2 ? tmp38448 : tmp38450;
  assign tmp38454 = l1 ? tmp35833 : tmp37064;
  assign tmp38455 = l1 ? tmp36894 : tmp36954;
  assign tmp38453 = s0 ? tmp38454 : tmp38455;
  assign tmp38456 = ~(l1 ? tmp35714 : tmp37067);
  assign tmp38452 = s1 ? tmp38453 : tmp38456;
  assign tmp38451 = s2 ? tmp38452 : tmp36895;
  assign tmp38446 = s3 ? tmp38447 : tmp38451;
  assign tmp38432 = s4 ? tmp38433 : tmp38446;
  assign tmp38461 = s0 ? tmp38443 : tmp35850;
  assign tmp38460 = s1 ? tmp38461 : tmp38300;
  assign tmp38463 = ~(l2 ? 1 : tmp35724);
  assign tmp38462 = s1 ? tmp37638 : tmp38463;
  assign tmp38459 = s2 ? tmp38460 : tmp38462;
  assign tmp38466 = ~(l1 ? tmp35833 : tmp35779);
  assign tmp38465 = s1 ? tmp36906 : tmp38466;
  assign tmp38464 = ~(s2 ? tmp35997 : tmp38465);
  assign tmp38458 = s3 ? tmp38459 : tmp38464;
  assign tmp38470 = ~(l1 ? tmp35786 : tmp36954);
  assign tmp38469 = s1 ? tmp36000 : tmp38470;
  assign tmp38471 = l1 ? tmp35714 : tmp35865;
  assign tmp38468 = s2 ? tmp38469 : tmp38471;
  assign tmp38472 = s1 ? tmp37173 : tmp38471;
  assign tmp38467 = ~(s3 ? tmp38468 : tmp38472);
  assign tmp38457 = s4 ? tmp38458 : tmp38467;
  assign tmp38431 = ~(s5 ? tmp38432 : tmp38457);
  assign tmp38402 = s6 ? tmp38403 : tmp38431;
  assign tmp38401 = s7 ? tmp35709 : tmp38402;
  assign tmp38400 = s8 ? tmp38394 : tmp38401;
  assign tmp38361 = s9 ? tmp38362 : tmp38400;
  assign tmp38479 = s3 ? tmp38327 : tmp38387;
  assign tmp38481 = s2 ? tmp38469 : tmp38172;
  assign tmp38480 = ~(s3 ? tmp38481 : tmp38171);
  assign tmp38478 = s4 ? tmp38479 : tmp38480;
  assign tmp38477 = ~(s5 ? tmp38319 : tmp38478);
  assign tmp38476 = s6 ? tmp38309 : tmp38477;
  assign tmp38475 = s7 ? tmp35709 : tmp38476;
  assign tmp38474 = s8 ? tmp38475 : tmp35709;
  assign tmp38486 = s4 ? tmp38382 : tmp38399;
  assign tmp38485 = ~(s5 ? tmp38376 : tmp38486);
  assign tmp38484 = s6 ? tmp38365 : tmp38485;
  assign tmp38483 = s7 ? tmp38484 : tmp38402;
  assign tmp38487 = s7 ? tmp38395 : tmp38476;
  assign tmp38482 = s8 ? tmp38483 : tmp38487;
  assign tmp38473 = s9 ? tmp38474 : tmp38482;
  assign tmp38360 = s10 ? tmp38361 : tmp38473;
  assign tmp38491 = s7 ? tmp38364 : tmp38402;
  assign tmp38490 = s8 ? tmp38491 : tmp38487;
  assign tmp38489 = s9 ? tmp38474 : tmp38490;
  assign tmp38488 = s10 ? tmp38361 : tmp38489;
  assign tmp38359 = s11 ? tmp38360 : tmp38488;
  assign tmp38090 = s12 ? tmp38091 : tmp38359;
  assign tmp38502 = s1 ? tmp35842 : tmp35866;
  assign tmp38501 = ~(s2 ? tmp38502 : tmp37813);
  assign tmp38500 = s3 ? tmp37808 : tmp38501;
  assign tmp38504 = s2 ? tmp37818 : tmp35779;
  assign tmp38503 = ~(s3 ? tmp37815 : tmp38504);
  assign tmp38499 = s4 ? tmp38500 : tmp38503;
  assign tmp38498 = ~(s5 ? tmp38068 : tmp38499);
  assign tmp38497 = s6 ? tmp37751 : tmp38498;
  assign tmp38496 = s7 ? tmp35709 : tmp38497;
  assign tmp38512 = ~(l2 ? tmp35727 : tmp35719);
  assign tmp38511 = l1 ? tmp35904 : tmp38512;
  assign tmp38514 = l1 ? tmp35908 : tmp35719;
  assign tmp38513 = ~(s0 ? tmp36436 : tmp38514);
  assign tmp38510 = s1 ? tmp38511 : tmp38513;
  assign tmp38518 = ~(l1 ? tmp36098 : tmp35909);
  assign tmp38517 = s0 ? tmp36441 : tmp38518;
  assign tmp38520 = l1 ? tmp36098 : tmp35909;
  assign tmp38519 = ~(s0 ? tmp36436 : tmp38520);
  assign tmp38516 = s1 ? tmp38517 : tmp38519;
  assign tmp38523 = ~(l1 ? tmp35904 : tmp38512);
  assign tmp38522 = s0 ? tmp38520 : tmp38523;
  assign tmp38521 = ~(s1 ? tmp36618 : tmp38522);
  assign tmp38515 = s2 ? tmp38516 : tmp38521;
  assign tmp38509 = s3 ? tmp38510 : tmp38515;
  assign tmp38528 = l1 ? tmp35768 : tmp35719;
  assign tmp38527 = s0 ? tmp38528 : tmp36456;
  assign tmp38529 = ~(s0 ? tmp38511 : tmp38518);
  assign tmp38526 = s1 ? tmp38527 : tmp38529;
  assign tmp38531 = s0 ? tmp38511 : tmp36115;
  assign tmp38530 = ~(s1 ? tmp38531 : tmp36147);
  assign tmp38525 = s2 ? tmp38526 : tmp38530;
  assign tmp38536 = l2 ? tmp35765 : tmp35720;
  assign tmp38535 = ~(l1 ? tmp35904 : tmp38536);
  assign tmp38534 = s0 ? tmp38520 : tmp38535;
  assign tmp38537 = s0 ? tmp37779 : tmp38520;
  assign tmp38533 = s1 ? tmp38534 : tmp38537;
  assign tmp38532 = s2 ? tmp37772 : tmp38533;
  assign tmp38524 = ~(s3 ? tmp38525 : tmp38532);
  assign tmp38508 = s4 ? tmp38509 : tmp38524;
  assign tmp38543 = s0 ? tmp38514 : tmp36474;
  assign tmp38542 = s1 ? tmp38543 : tmp36475;
  assign tmp38545 = l1 ? tmp35904 : 1;
  assign tmp38547 = l1 ? tmp35904 : tmp38536;
  assign tmp38546 = s0 ? tmp38547 : tmp35775;
  assign tmp38544 = ~(s1 ? tmp38545 : tmp38546);
  assign tmp38541 = s2 ? tmp38542 : tmp38544;
  assign tmp38550 = l1 ? tmp35777 : tmp35909;
  assign tmp38549 = s1 ? tmp36482 : tmp38550;
  assign tmp38553 = l1 ? tmp35777 : tmp35719;
  assign tmp38552 = s0 ? tmp38520 : tmp38553;
  assign tmp38551 = s1 ? tmp37791 : tmp38552;
  assign tmp38548 = s2 ? tmp38549 : tmp38551;
  assign tmp38540 = s3 ? tmp38541 : tmp38548;
  assign tmp38557 = s0 ? tmp37797 : tmp38520;
  assign tmp38556 = s1 ? tmp38557 : tmp36490;
  assign tmp38558 = ~(l1 ? tmp35914 : 1);
  assign tmp38555 = s2 ? tmp38556 : tmp38558;
  assign tmp38562 = l1 ? 1 : tmp35909;
  assign tmp38563 = l1 ? tmp35821 : tmp35719;
  assign tmp38561 = s0 ? tmp38562 : tmp38563;
  assign tmp38564 = ~(l1 ? tmp35926 : tmp35765);
  assign tmp38560 = s1 ? tmp38561 : tmp38564;
  assign tmp38559 = s2 ? tmp38560 : tmp38071;
  assign tmp38554 = s3 ? tmp38555 : tmp38559;
  assign tmp38539 = s4 ? tmp38540 : tmp38554;
  assign tmp38569 = s0 ? tmp38550 : tmp35850;
  assign tmp38568 = s1 ? tmp38569 : tmp35992;
  assign tmp38567 = s2 ? tmp38568 : tmp36501;
  assign tmp38571 = s1 ? tmp35812 : tmp36001;
  assign tmp38570 = ~(s2 ? tmp38502 : tmp38571);
  assign tmp38566 = s3 ? tmp38567 : tmp38570;
  assign tmp38573 = s2 ? tmp37816 : tmp36009;
  assign tmp38576 = l1 ? tmp35926 : tmp35812;
  assign tmp38575 = s1 ? tmp37819 : tmp38576;
  assign tmp38574 = s2 ? tmp38575 : tmp35779;
  assign tmp38572 = ~(s3 ? tmp38573 : tmp38574);
  assign tmp38565 = s4 ? tmp38566 : tmp38572;
  assign tmp38538 = ~(s5 ? tmp38539 : tmp38565);
  assign tmp38507 = s6 ? tmp38508 : tmp38538;
  assign tmp38506 = s7 ? tmp35709 : tmp38507;
  assign tmp38505 = s8 ? tmp38496 : tmp38506;
  assign tmp38495 = s9 ? tmp38496 : tmp38505;
  assign tmp38578 = s8 ? tmp38496 : tmp35709;
  assign tmp38583 = s4 ? tmp38500 : tmp37814;
  assign tmp38582 = ~(s5 ? tmp38068 : tmp38583);
  assign tmp38581 = s6 ? tmp37751 : tmp38582;
  assign tmp38587 = ~(s3 ? tmp38573 : tmp38575);
  assign tmp38586 = s4 ? tmp38566 : tmp38587;
  assign tmp38585 = ~(s5 ? tmp38539 : tmp38586);
  assign tmp38584 = s6 ? tmp38508 : tmp38585;
  assign tmp38580 = s7 ? tmp38581 : tmp38584;
  assign tmp38579 = s8 ? tmp38580 : tmp38581;
  assign tmp38577 = s9 ? tmp38578 : tmp38579;
  assign tmp38494 = s10 ? tmp38495 : tmp38577;
  assign tmp38591 = s7 ? tmp38497 : tmp38507;
  assign tmp38590 = s8 ? tmp38591 : tmp38497;
  assign tmp38589 = s9 ? tmp38578 : tmp38590;
  assign tmp38588 = s10 ? tmp38495 : tmp38589;
  assign tmp38493 = s11 ? tmp38494 : tmp38588;
  assign tmp38602 = l1 ? tmp35729 : tmp35719;
  assign tmp38601 = ~(s0 ? tmp36512 : tmp38602);
  assign tmp38600 = s1 ? tmp37433 : tmp38601;
  assign tmp38606 = ~(l1 ? tmp35739 : tmp36576);
  assign tmp38605 = s0 ? tmp37439 : tmp38606;
  assign tmp38607 = ~(s0 ? tmp37443 : tmp37479);
  assign tmp38604 = s1 ? tmp38605 : tmp38607;
  assign tmp38609 = s0 ? tmp37479 : tmp37448;
  assign tmp38608 = ~(s1 ? tmp37446 : tmp38609);
  assign tmp38603 = s2 ? tmp38604 : tmp38608;
  assign tmp38599 = s3 ? tmp38600 : tmp38603;
  assign tmp38614 = l1 ? tmp35743 : tmp35719;
  assign tmp38613 = s0 ? tmp38614 : tmp36456;
  assign tmp38615 = ~(s0 ? tmp37433 : tmp38606);
  assign tmp38612 = s1 ? tmp38613 : tmp38615;
  assign tmp38616 = ~(s1 ? tmp37456 : tmp36147);
  assign tmp38611 = s2 ? tmp38612 : tmp38616;
  assign tmp38620 = ~(l1 ? tmp35714 : tmp36596);
  assign tmp38619 = s0 ? tmp37479 : tmp38620;
  assign tmp38621 = s0 ? tmp37122 : tmp37479;
  assign tmp38618 = s1 ? tmp38619 : tmp38621;
  assign tmp38617 = s2 ? tmp36592 : tmp38618;
  assign tmp38610 = ~(s3 ? tmp38611 : tmp38617);
  assign tmp38598 = s4 ? tmp38599 : tmp38610;
  assign tmp38627 = s0 ? tmp38602 : tmp36474;
  assign tmp38626 = s1 ? tmp38627 : tmp37469;
  assign tmp38630 = l1 ? tmp35714 : tmp36596;
  assign tmp38629 = s0 ? tmp38630 : tmp35775;
  assign tmp38628 = ~(s1 ? tmp37174 : tmp38629);
  assign tmp38625 = s2 ? tmp38626 : tmp38628;
  assign tmp38634 = l1 ? tmp35815 : tmp35973;
  assign tmp38633 = s0 ? tmp37479 : tmp38634;
  assign tmp38632 = s1 ? tmp37139 : tmp38633;
  assign tmp38631 = s2 ? tmp37474 : tmp38632;
  assign tmp38624 = s3 ? tmp38625 : tmp38631;
  assign tmp38637 = s1 ? tmp37483 : tmp36490;
  assign tmp38636 = s2 ? tmp38637 : tmp36560;
  assign tmp38635 = s3 ? tmp38636 : tmp37484;
  assign tmp38623 = s4 ? tmp38624 : tmp38635;
  assign tmp38640 = ~(s2 ? tmp35997 : tmp37165);
  assign tmp38639 = s3 ? tmp37490 : tmp38640;
  assign tmp38644 = s0 ? tmp35881 : tmp37170;
  assign tmp38643 = s1 ? tmp36000 : tmp38644;
  assign tmp38642 = s2 ? tmp38643 : tmp37174;
  assign tmp38645 = s2 ? tmp37172 : tmp35881;
  assign tmp38641 = ~(s3 ? tmp38642 : tmp38645);
  assign tmp38638 = s4 ? tmp38639 : tmp38641;
  assign tmp38622 = ~(s5 ? tmp38623 : tmp38638);
  assign tmp38597 = s6 ? tmp38598 : tmp38622;
  assign tmp38596 = s7 ? tmp35709 : tmp38597;
  assign tmp38650 = s3 ? tmp37563 : tmp38640;
  assign tmp38654 = s0 ? tmp35881 : tmp37248;
  assign tmp38653 = s1 ? tmp36000 : tmp38654;
  assign tmp38652 = s2 ? tmp38653 : tmp37571;
  assign tmp38651 = ~(s3 ? tmp38652 : tmp38645);
  assign tmp38649 = s4 ? tmp38650 : tmp38651;
  assign tmp38648 = ~(s5 ? tmp37534 : tmp38649);
  assign tmp38647 = s6 ? tmp37500 : tmp38648;
  assign tmp38646 = s7 ? tmp35709 : tmp38647;
  assign tmp38595 = s8 ? tmp38596 : tmp38646;
  assign tmp38662 = s0 ? tmp37584 : tmp37656;
  assign tmp38663 = ~(s0 ? tmp37587 : tmp37659);
  assign tmp38661 = s1 ? tmp38662 : tmp38663;
  assign tmp38664 = ~(s1 ? tmp37590 : tmp37662);
  assign tmp38660 = s2 ? tmp38661 : tmp38664;
  assign tmp38659 = s3 ? tmp37648 : tmp38660;
  assign tmp38658 = s4 ? tmp38659 : tmp37664;
  assign tmp38669 = s1 ? tmp37682 : tmp37612;
  assign tmp38668 = s2 ? tmp38669 : tmp37683;
  assign tmp38671 = s1 ? tmp37619 : tmp37476;
  assign tmp38670 = s2 ? tmp38671 : tmp37690;
  assign tmp38667 = s3 ? tmp38668 : tmp38670;
  assign tmp38666 = s4 ? tmp38667 : tmp37692;
  assign tmp38674 = s2 ? tmp37491 : tmp38462;
  assign tmp38673 = s3 ? tmp38674 : tmp38640;
  assign tmp38672 = s4 ? tmp38673 : tmp38641;
  assign tmp38665 = ~(s5 ? tmp38666 : tmp38672);
  assign tmp38657 = s6 ? tmp38658 : tmp38665;
  assign tmp38656 = s7 ? tmp35709 : tmp38657;
  assign tmp38655 = s8 ? tmp38646 : tmp38656;
  assign tmp38594 = s9 ? tmp38595 : tmp38655;
  assign tmp38679 = ~(s5 ? tmp37678 : tmp38638);
  assign tmp38678 = s6 ? tmp37646 : tmp38679;
  assign tmp38677 = s7 ? tmp35709 : tmp38678;
  assign tmp38676 = s8 ? tmp38677 : tmp35709;
  assign tmp38685 = ~(s3 ? tmp38642 : tmp37172);
  assign tmp38684 = s4 ? tmp38639 : tmp38685;
  assign tmp38683 = ~(s5 ? tmp38623 : tmp38684);
  assign tmp38682 = s6 ? tmp38598 : tmp38683;
  assign tmp38688 = s4 ? tmp38673 : tmp38685;
  assign tmp38687 = ~(s5 ? tmp38666 : tmp38688);
  assign tmp38686 = s6 ? tmp38658 : tmp38687;
  assign tmp38681 = s7 ? tmp38682 : tmp38686;
  assign tmp38693 = ~(s3 ? tmp38652 : tmp37172);
  assign tmp38692 = s4 ? tmp38650 : tmp38693;
  assign tmp38691 = ~(s5 ? tmp37534 : tmp38692);
  assign tmp38690 = s6 ? tmp37500 : tmp38691;
  assign tmp38695 = ~(s5 ? tmp37678 : tmp38684);
  assign tmp38694 = s6 ? tmp37646 : tmp38695;
  assign tmp38689 = s7 ? tmp38690 : tmp38694;
  assign tmp38680 = s8 ? tmp38681 : tmp38689;
  assign tmp38675 = s9 ? tmp38676 : tmp38680;
  assign tmp38593 = s10 ? tmp38594 : tmp38675;
  assign tmp38699 = s7 ? tmp38597 : tmp38657;
  assign tmp38700 = s7 ? tmp38647 : tmp38678;
  assign tmp38698 = s8 ? tmp38699 : tmp38700;
  assign tmp38697 = s9 ? tmp38676 : tmp38698;
  assign tmp38696 = s10 ? tmp38594 : tmp38697;
  assign tmp38592 = s11 ? tmp38593 : tmp38696;
  assign tmp38492 = s12 ? tmp38493 : tmp38592;
  assign tmp38089 = s13 ? tmp38090 : tmp38492;
  assign tmp37724 = s14 ? tmp37725 : tmp38089;
  assign tmp35701 = s15 ? tmp35702 : tmp37724;
  assign tmp38716 = l1 ? tmp35865 : tmp35726;
  assign tmp38715 = s0 ? tmp38716 : tmp35772;
  assign tmp38714 = ~(s1 ? tmp35772 : tmp38715);
  assign tmp38713 = s2 ? tmp35969 : tmp38714;
  assign tmp38712 = s3 ? tmp38713 : tmp36065;
  assign tmp38711 = s4 ? tmp36045 : tmp38712;
  assign tmp38710 = ~(s5 ? tmp38711 : tmp36071);
  assign tmp38709 = s6 ? tmp36012 : tmp38710;
  assign tmp38708 = s7 ? tmp35709 : tmp38709;
  assign tmp38707 = s8 ? tmp35708 : tmp38708;
  assign tmp38706 = s9 ? tmp38707 : tmp38708;
  assign tmp38718 = s8 ? tmp38708 : tmp35709;
  assign tmp38727 = ~(l1 ? tmp35865 : tmp36096);
  assign tmp38726 = s1 ? tmp36332 : tmp38727;
  assign tmp38725 = s2 ? tmp38726 : tmp36414;
  assign tmp38724 = s3 ? tmp38725 : tmp36338;
  assign tmp38731 = l1 ? tmp35865 : tmp35744;
  assign tmp38730 = ~(s1 ? tmp35772 : tmp38731);
  assign tmp38729 = s2 ? tmp36346 : tmp38730;
  assign tmp38733 = s1 ? tmp36351 : tmp35984;
  assign tmp38732 = s2 ? tmp38733 : tmp35985;
  assign tmp38728 = s3 ? tmp38729 : tmp38732;
  assign tmp38723 = s4 ? tmp38724 : tmp38728;
  assign tmp38722 = ~(s5 ? tmp38723 : tmp36155);
  assign tmp38721 = s6 ? tmp36297 : tmp38722;
  assign tmp38720 = s7 ? tmp36220 : tmp38721;
  assign tmp38739 = ~(s1 ? tmp35772 : tmp38716);
  assign tmp38738 = s2 ? tmp35969 : tmp38739;
  assign tmp38737 = s3 ? tmp38738 : tmp36065;
  assign tmp38736 = s4 ? tmp36045 : tmp38737;
  assign tmp38735 = ~(s5 ? tmp38736 : tmp36071);
  assign tmp38734 = s6 ? tmp36012 : tmp38735;
  assign tmp38719 = s8 ? tmp38720 : tmp38734;
  assign tmp38717 = s9 ? tmp38718 : tmp38719;
  assign tmp38705 = s10 ? tmp38706 : tmp38717;
  assign tmp38750 = s0 ? tmp38731 : tmp35772;
  assign tmp38749 = ~(s1 ? tmp35772 : tmp38750);
  assign tmp38748 = s2 ? tmp36346 : tmp38749;
  assign tmp38747 = s3 ? tmp38748 : tmp38732;
  assign tmp38746 = s4 ? tmp38724 : tmp38747;
  assign tmp38745 = ~(s5 ? tmp38746 : tmp36155);
  assign tmp38744 = s6 ? tmp36297 : tmp38745;
  assign tmp38743 = s7 ? tmp35899 : tmp38744;
  assign tmp38742 = s8 ? tmp38743 : tmp38709;
  assign tmp38741 = s9 ? tmp38718 : tmp38742;
  assign tmp38740 = s10 ? tmp38706 : tmp38741;
  assign tmp38704 = s11 ? tmp38705 : tmp38740;
  assign tmp38762 = s0 ? tmp35827 : tmp35766;
  assign tmp38761 = ~(s1 ? tmp36533 : tmp38762);
  assign tmp38760 = s2 ? tmp36527 : tmp38761;
  assign tmp38764 = s1 ? tmp36512 : tmp36259;
  assign tmp38763 = s2 ? tmp38764 : tmp36536;
  assign tmp38759 = ~(s3 ? tmp38760 : tmp38763);
  assign tmp38758 = s4 ? tmp36508 : tmp38759;
  assign tmp38757 = s6 ? tmp38758 : tmp36540;
  assign tmp38756 = s7 ? tmp35709 : tmp38757;
  assign tmp38755 = s8 ? tmp36429 : tmp38756;
  assign tmp38771 = l1 ? tmp35926 : tmp35725;
  assign tmp38770 = s1 ? tmp38771 : tmp36511;
  assign tmp38775 = l1 ? tmp35865 : tmp35768;
  assign tmp38776 = ~(l1 ? tmp35916 : tmp36576);
  assign tmp38774 = s0 ? tmp38775 : tmp38776;
  assign tmp38778 = l1 ? tmp35723 : tmp35914;
  assign tmp38779 = l1 ? tmp35916 : tmp36576;
  assign tmp38777 = ~(s0 ? tmp38778 : tmp38779);
  assign tmp38773 = s1 ? tmp38774 : tmp38777;
  assign tmp38781 = s0 ? tmp38778 : tmp36448;
  assign tmp38783 = ~(l1 ? tmp35926 : tmp35725);
  assign tmp38782 = s0 ? tmp38779 : tmp38783;
  assign tmp38780 = ~(s1 ? tmp38781 : tmp38782);
  assign tmp38772 = s2 ? tmp38773 : tmp38780;
  assign tmp38769 = s3 ? tmp38770 : tmp38772;
  assign tmp38787 = ~(s0 ? tmp38771 : tmp38776);
  assign tmp38786 = s1 ? tmp36528 : tmp38787;
  assign tmp38789 = s0 ? tmp38771 : tmp35761;
  assign tmp38788 = ~(s1 ? tmp38789 : tmp38762);
  assign tmp38785 = s2 ? tmp38786 : tmp38788;
  assign tmp38793 = ~(l1 ? tmp35926 : tmp36596);
  assign tmp38792 = s0 ? tmp38779 : tmp38793;
  assign tmp38794 = s0 ? tmp35944 : tmp38779;
  assign tmp38791 = s1 ? tmp38792 : tmp38794;
  assign tmp38790 = s2 ? tmp38764 : tmp38791;
  assign tmp38784 = ~(s3 ? tmp38785 : tmp38790);
  assign tmp38768 = s4 ? tmp38769 : tmp38784;
  assign tmp38800 = ~(l1 ? tmp35865 : tmp35768);
  assign tmp38799 = s1 ? tmp36545 : tmp38800;
  assign tmp38803 = l1 ? tmp35926 : tmp36596;
  assign tmp38802 = s0 ? tmp38803 : tmp36550;
  assign tmp38801 = ~(s1 ? tmp36167 : tmp38802);
  assign tmp38798 = s2 ? tmp38799 : tmp38801;
  assign tmp38806 = l1 ? tmp35767 : tmp35914;
  assign tmp38805 = s1 ? tmp38806 : tmp36483;
  assign tmp38804 = s2 ? tmp38805 : tmp36554;
  assign tmp38797 = s3 ? tmp38798 : tmp38804;
  assign tmp38796 = s4 ? tmp38797 : tmp36556;
  assign tmp38795 = ~(s5 ? tmp38796 : tmp36496);
  assign tmp38767 = s6 ? tmp38768 : tmp38795;
  assign tmp38766 = s7 ? tmp35709 : tmp38767;
  assign tmp38765 = s8 ? tmp38756 : tmp38766;
  assign tmp38754 = s9 ? tmp38755 : tmp38765;
  assign tmp38808 = s8 ? tmp38756 : tmp35709;
  assign tmp38814 = s2 ? tmp36535 : tmp38791;
  assign tmp38813 = ~(s3 ? tmp38785 : tmp38814);
  assign tmp38812 = s4 ? tmp38769 : tmp38813;
  assign tmp38811 = s6 ? tmp38812 : tmp38795;
  assign tmp38810 = s7 ? tmp36626 : tmp38811;
  assign tmp38817 = ~(s3 ? tmp38760 : tmp36534);
  assign tmp38816 = s4 ? tmp36508 : tmp38817;
  assign tmp38815 = s6 ? tmp38816 : tmp36540;
  assign tmp38809 = s8 ? tmp38810 : tmp38815;
  assign tmp38807 = s9 ? tmp38808 : tmp38809;
  assign tmp38753 = s10 ? tmp38754 : tmp38807;
  assign tmp38821 = s7 ? tmp36430 : tmp38767;
  assign tmp38820 = s8 ? tmp38821 : tmp38757;
  assign tmp38819 = s9 ? tmp38808 : tmp38820;
  assign tmp38818 = s10 ? tmp38754 : tmp38819;
  assign tmp38752 = s11 ? tmp38753 : tmp38818;
  assign tmp38751 = s12 ? tmp36232 : tmp38752;
  assign tmp38703 = s13 ? tmp38704 : tmp38751;
  assign tmp38832 = l1 ? tmp35926 : tmp36677;
  assign tmp38834 = l1 ? tmp35723 : tmp36680;
  assign tmp38835 = l1 ? tmp36017 : tmp36682;
  assign tmp38833 = ~(s0 ? tmp38834 : tmp38835);
  assign tmp38831 = s1 ? tmp38832 : tmp38833;
  assign tmp38839 = l1 ? tmp35865 : tmp35717;
  assign tmp38838 = s0 ? tmp38839 : tmp36244;
  assign tmp38840 = ~(s0 ? tmp38834 : tmp36246);
  assign tmp38837 = s1 ? tmp38838 : tmp38840;
  assign tmp38842 = s0 ? tmp38834 : tmp35749;
  assign tmp38844 = ~(l1 ? tmp35926 : tmp36677);
  assign tmp38843 = s0 ? tmp36246 : tmp38844;
  assign tmp38841 = ~(s1 ? tmp38842 : tmp38843);
  assign tmp38836 = s2 ? tmp38837 : tmp38841;
  assign tmp38830 = s3 ? tmp38831 : tmp38836;
  assign tmp38849 = l1 ? tmp35723 : tmp36682;
  assign tmp38848 = s0 ? tmp38849 : tmp35757;
  assign tmp38850 = ~(s0 ? tmp38832 : tmp36244);
  assign tmp38847 = s1 ? tmp38848 : tmp38850;
  assign tmp38852 = s0 ? tmp38832 : tmp35761;
  assign tmp38853 = l1 ? tmp35736 : tmp35955;
  assign tmp38851 = ~(s1 ? tmp38852 : tmp38853);
  assign tmp38846 = s2 ? tmp38847 : tmp38851;
  assign tmp38855 = s1 ? tmp38834 : tmp35938;
  assign tmp38857 = s0 ? tmp35938 : tmp36246;
  assign tmp38856 = s1 ? tmp36261 : tmp38857;
  assign tmp38854 = s2 ? tmp38855 : tmp38856;
  assign tmp38845 = ~(s3 ? tmp38846 : tmp38854);
  assign tmp38829 = s4 ? tmp38830 : tmp38845;
  assign tmp38863 = s0 ? tmp38835 : tmp35793;
  assign tmp38864 = ~(l1 ? tmp35865 : tmp35717);
  assign tmp38862 = s1 ? tmp38863 : tmp38864;
  assign tmp38865 = ~(s1 ? tmp36741 : tmp36273);
  assign tmp38861 = s2 ? tmp38862 : tmp38865;
  assign tmp38869 = ~(l1 ? tmp35767 : tmp36680);
  assign tmp38868 = s0 ? 1 : tmp38869;
  assign tmp38867 = s1 ? tmp38868 : tmp36279;
  assign tmp38870 = ~(s1 ? tmp36293 : tmp36282);
  assign tmp38866 = ~(s2 ? tmp38867 : tmp38870);
  assign tmp38860 = s3 ? tmp38861 : tmp38866;
  assign tmp38874 = s0 ? tmp35971 : tmp36246;
  assign tmp38876 = l1 ? tmp35736 : tmp35767;
  assign tmp38875 = ~(s0 ? tmp35823 : tmp38876);
  assign tmp38873 = s1 ? tmp38874 : tmp38875;
  assign tmp38877 = ~(l1 ? tmp35865 : tmp36713);
  assign tmp38872 = s2 ? tmp38873 : tmp38877;
  assign tmp38881 = l1 ? tmp36070 : tmp35882;
  assign tmp38880 = s0 ? tmp36732 : tmp38881;
  assign tmp38879 = s1 ? tmp38880 : tmp36287;
  assign tmp38878 = s2 ? tmp38879 : tmp35985;
  assign tmp38871 = s3 ? tmp38872 : tmp38878;
  assign tmp38859 = s4 ? tmp38860 : tmp38871;
  assign tmp38858 = ~(s5 ? tmp38859 : tmp36733);
  assign tmp38828 = s6 ? tmp38829 : tmp38858;
  assign tmp38827 = s7 ? tmp35709 : tmp38828;
  assign tmp38888 = l1 ? tmp35926 : tmp35723;
  assign tmp38890 = l1 ? tmp36017 : tmp36751;
  assign tmp38889 = ~(s0 ? tmp38834 : tmp38890);
  assign tmp38887 = s1 ? tmp38888 : tmp38889;
  assign tmp38894 = l1 ? tmp35865 : tmp35737;
  assign tmp38893 = s0 ? tmp38894 : tmp35915;
  assign tmp38896 = l1 ? tmp35723 : tmp36758;
  assign tmp38895 = ~(s0 ? tmp38896 : tmp35921);
  assign tmp38892 = s1 ? tmp38893 : tmp38895;
  assign tmp38898 = s0 ? tmp38896 : tmp35749;
  assign tmp38900 = ~(l1 ? tmp35926 : tmp35723);
  assign tmp38899 = s0 ? tmp35921 : tmp38900;
  assign tmp38897 = ~(s1 ? tmp38898 : tmp38899);
  assign tmp38891 = s2 ? tmp38892 : tmp38897;
  assign tmp38886 = s3 ? tmp38887 : tmp38891;
  assign tmp38905 = l1 ? tmp35723 : tmp36751;
  assign tmp38904 = s0 ? tmp38905 : tmp35757;
  assign tmp38906 = ~(s0 ? tmp38888 : tmp35915);
  assign tmp38903 = s1 ? tmp38904 : tmp38906;
  assign tmp38908 = s0 ? tmp38888 : tmp35761;
  assign tmp38907 = ~(s1 ? tmp38908 : tmp38853);
  assign tmp38902 = s2 ? tmp38903 : tmp38907;
  assign tmp38911 = s0 ? tmp35938 : tmp35921;
  assign tmp38910 = s1 ? tmp35940 : tmp38911;
  assign tmp38909 = s2 ? tmp38855 : tmp38910;
  assign tmp38901 = ~(s3 ? tmp38902 : tmp38909);
  assign tmp38885 = s4 ? tmp38886 : tmp38901;
  assign tmp38917 = s0 ? tmp38890 : tmp35793;
  assign tmp38918 = ~(l1 ? tmp35865 : tmp35737);
  assign tmp38916 = s1 ? tmp38917 : tmp38918;
  assign tmp38919 = ~(s1 ? tmp36006 : tmp35956);
  assign tmp38915 = s2 ? tmp38916 : tmp38919;
  assign tmp38923 = ~(l1 ? tmp35767 : tmp36758);
  assign tmp38922 = s0 ? 1 : tmp38923;
  assign tmp38925 = ~(l1 ? tmp35777 : tmp35917);
  assign tmp38924 = s0 ? 1 : tmp38925;
  assign tmp38921 = s1 ? tmp38922 : tmp38924;
  assign tmp38926 = ~(s1 ? tmp36293 : tmp35964);
  assign tmp38920 = ~(s2 ? tmp38921 : tmp38926);
  assign tmp38914 = s3 ? tmp38915 : tmp38920;
  assign tmp38929 = ~(l1 ? tmp35865 : tmp35955);
  assign tmp38928 = s2 ? tmp38873 : tmp38929;
  assign tmp38932 = s0 ? tmp35981 : tmp38881;
  assign tmp38931 = s1 ? tmp38932 : tmp36287;
  assign tmp38930 = s2 ? tmp38931 : tmp35985;
  assign tmp38927 = s3 ? tmp38928 : tmp38930;
  assign tmp38913 = s4 ? tmp38914 : tmp38927;
  assign tmp38912 = ~(s5 ? tmp38913 : tmp36797);
  assign tmp38884 = s6 ? tmp38885 : tmp38912;
  assign tmp38883 = s7 ? tmp35709 : tmp38884;
  assign tmp38882 = s8 ? tmp38827 : tmp38883;
  assign tmp38826 = s9 ? tmp38827 : tmp38882;
  assign tmp38934 = s8 ? tmp38827 : tmp35709;
  assign tmp38942 = s1 ? tmp38922 : tmp38925;
  assign tmp38941 = ~(s2 ? tmp38942 : tmp38926);
  assign tmp38940 = s3 ? tmp38915 : tmp38941;
  assign tmp38939 = s4 ? tmp38940 : tmp38927;
  assign tmp38938 = ~(s5 ? tmp38939 : tmp36797);
  assign tmp38937 = s6 ? tmp38885 : tmp38938;
  assign tmp38936 = s7 ? tmp36808 : tmp38937;
  assign tmp38948 = s1 ? tmp38868 : tmp36280;
  assign tmp38947 = ~(s2 ? tmp38948 : tmp38870);
  assign tmp38946 = s3 ? tmp38861 : tmp38947;
  assign tmp38945 = s4 ? tmp38946 : tmp38871;
  assign tmp38944 = ~(s5 ? tmp38945 : tmp36733);
  assign tmp38943 = s6 ? tmp38829 : tmp38944;
  assign tmp38935 = s8 ? tmp38936 : tmp38943;
  assign tmp38933 = s9 ? tmp38934 : tmp38935;
  assign tmp38825 = s10 ? tmp38826 : tmp38933;
  assign tmp38952 = s7 ? tmp36641 : tmp38884;
  assign tmp38951 = s8 ? tmp38952 : tmp38828;
  assign tmp38950 = s9 ? tmp38934 : tmp38951;
  assign tmp38949 = s10 ? tmp38826 : tmp38950;
  assign tmp38824 = s11 ? tmp38825 : tmp38949;
  assign tmp38960 = l1 ? tmp35926 : tmp36827;
  assign tmp38962 = l1 ? tmp36017 : tmp35740;
  assign tmp38961 = ~(s0 ? tmp35749 : tmp38962);
  assign tmp38959 = s1 ? tmp38960 : tmp38961;
  assign tmp38966 = l1 ? tmp35865 : tmp35723;
  assign tmp38967 = ~(l1 ? tmp35916 : tmp36835);
  assign tmp38965 = s0 ? tmp38966 : tmp38967;
  assign tmp38969 = l1 ? tmp35723 : tmp35736;
  assign tmp38970 = l1 ? tmp35916 : tmp36835;
  assign tmp38968 = ~(s0 ? tmp38969 : tmp38970);
  assign tmp38964 = s1 ? tmp38965 : tmp38968;
  assign tmp38972 = s0 ? tmp38969 : tmp35722;
  assign tmp38974 = ~(l1 ? tmp35926 : tmp36827);
  assign tmp38973 = s0 ? tmp38970 : tmp38974;
  assign tmp38971 = ~(s1 ? tmp38972 : tmp38973);
  assign tmp38963 = s2 ? tmp38964 : tmp38971;
  assign tmp38958 = s3 ? tmp38959 : tmp38963;
  assign tmp38979 = l1 ? tmp35723 : tmp35740;
  assign tmp38978 = s0 ? tmp38979 : tmp36530;
  assign tmp38980 = ~(s0 ? tmp38960 : tmp38967);
  assign tmp38977 = s1 ? tmp38978 : tmp38980;
  assign tmp38982 = s0 ? tmp38960 : tmp35761;
  assign tmp38981 = ~(s1 ? tmp38982 : tmp35824);
  assign tmp38976 = s2 ? tmp38977 : tmp38981;
  assign tmp38985 = s0 ? tmp38970 : tmp36857;
  assign tmp38986 = s0 ? tmp36853 : tmp38970;
  assign tmp38984 = s1 ? tmp38985 : tmp38986;
  assign tmp38983 = s2 ? tmp36852 : tmp38984;
  assign tmp38975 = ~(s3 ? tmp38976 : tmp38983);
  assign tmp38957 = s4 ? tmp38958 : tmp38975;
  assign tmp38992 = s0 ? tmp38962 : tmp36474;
  assign tmp38993 = ~(l1 ? tmp35865 : tmp35723);
  assign tmp38991 = s1 ? tmp38992 : tmp38993;
  assign tmp38996 = l1 ? 1 : tmp35723;
  assign tmp38995 = s0 ? tmp36870 : tmp38996;
  assign tmp38994 = ~(s1 ? tmp36912 : tmp38995);
  assign tmp38990 = s2 ? tmp38991 : tmp38994;
  assign tmp38999 = l1 ? tmp35767 : tmp35736;
  assign tmp38998 = s1 ? tmp38999 : tmp36873;
  assign tmp39001 = s0 ? tmp38970 : tmp36877;
  assign tmp39000 = s1 ? tmp36875 : tmp39001;
  assign tmp38997 = s2 ? tmp38998 : tmp39000;
  assign tmp38989 = s3 ? tmp38990 : tmp38997;
  assign tmp39005 = s0 ? tmp36883 : tmp38970;
  assign tmp39004 = s1 ? tmp39005 : tmp36884;
  assign tmp39007 = l1 ? tmp35865 : tmp35806;
  assign tmp39006 = ~(s1 ? tmp35827 : tmp39007);
  assign tmp39003 = s2 ? tmp39004 : tmp39006;
  assign tmp39011 = l1 ? tmp36070 : tmp36878;
  assign tmp39010 = s0 ? tmp36890 : tmp39011;
  assign tmp39009 = s1 ? tmp39010 : tmp36892;
  assign tmp39008 = s2 ? tmp39009 : tmp36895;
  assign tmp39002 = s3 ? tmp39003 : tmp39008;
  assign tmp38988 = s4 ? tmp38989 : tmp39002;
  assign tmp39016 = l1 ? 1 : tmp35744;
  assign tmp39015 = s1 ? tmp39016 : tmp35995;
  assign tmp39014 = s2 ? tmp36899 : tmp39015;
  assign tmp39013 = s3 ? tmp39014 : tmp36904;
  assign tmp39012 = s4 ? tmp39013 : tmp36908;
  assign tmp38987 = ~(s5 ? tmp38988 : tmp39012);
  assign tmp38956 = s6 ? tmp38957 : tmp38987;
  assign tmp38955 = s7 ? tmp35709 : tmp38956;
  assign tmp39018 = s8 ? tmp38955 : tmp35709;
  assign tmp39024 = s1 ? tmp39010 : tmp36985;
  assign tmp39023 = s2 ? tmp39024 : tmp36895;
  assign tmp39022 = s3 ? tmp39003 : tmp39023;
  assign tmp39021 = s4 ? tmp38989 : tmp39022;
  assign tmp39020 = ~(s5 ? tmp39021 : tmp39012);
  assign tmp39019 = s6 ? tmp38957 : tmp39020;
  assign tmp39017 = s9 ? tmp39018 : tmp39019;
  assign tmp38954 = s10 ? tmp38955 : tmp39017;
  assign tmp39026 = s9 ? tmp39018 : tmp38956;
  assign tmp39025 = s10 ? tmp38955 : tmp39026;
  assign tmp38953 = s11 ? tmp38954 : tmp39025;
  assign tmp38823 = s12 ? tmp38824 : tmp38953;
  assign tmp39037 = s2 ? tmp37157 : tmp37244;
  assign tmp39036 = s3 ? tmp39037 : tmp38640;
  assign tmp39035 = s4 ? tmp39036 : tmp37401;
  assign tmp39034 = ~(s5 ? tmp37124 : tmp39035);
  assign tmp39033 = s6 ? tmp37092 : tmp39034;
  assign tmp39032 = s7 ? tmp35709 : tmp39033;
  assign tmp39042 = s3 ? tmp37241 : tmp38640;
  assign tmp39041 = s4 ? tmp39042 : tmp37412;
  assign tmp39040 = ~(s5 ? tmp37214 : tmp39041);
  assign tmp39039 = s6 ? tmp37177 : tmp39040;
  assign tmp39038 = s7 ? tmp35709 : tmp39039;
  assign tmp39031 = s8 ? tmp39032 : tmp39038;
  assign tmp39049 = s2 ? tmp37242 : tmp37159;
  assign tmp39048 = s3 ? tmp39049 : tmp37162;
  assign tmp39051 = s2 ? tmp37247 : tmp37171;
  assign tmp39050 = ~(s3 ? tmp39051 : tmp37172);
  assign tmp39047 = s4 ? tmp39048 : tmp39050;
  assign tmp39046 = ~(s5 ? tmp37214 : tmp39047);
  assign tmp39045 = s6 ? tmp37177 : tmp39046;
  assign tmp39044 = s7 ? tmp35709 : tmp39045;
  assign tmp39043 = s8 ? tmp39038 : tmp39044;
  assign tmp39030 = s9 ? tmp39031 : tmp39043;
  assign tmp39053 = s8 ? tmp39038 : tmp35709;
  assign tmp39060 = l1 ? tmp37181 : tmp36677;
  assign tmp39062 = l1 ? tmp37184 : tmp36682;
  assign tmp39061 = ~(s0 ? tmp36679 : tmp39062);
  assign tmp39059 = s1 ? tmp39060 : tmp39061;
  assign tmp39066 = l1 ? tmp35724 : tmp35717;
  assign tmp39067 = ~(l1 ? tmp37190 : tmp35882);
  assign tmp39065 = s0 ? tmp39066 : tmp39067;
  assign tmp39069 = l1 ? tmp37193 : tmp36680;
  assign tmp39070 = l1 ? tmp37190 : tmp35882;
  assign tmp39068 = ~(s0 ? tmp39069 : tmp39070);
  assign tmp39064 = s1 ? tmp39065 : tmp39068;
  assign tmp39072 = s0 ? tmp39069 : tmp36652;
  assign tmp39074 = ~(l1 ? tmp37181 : tmp36677);
  assign tmp39073 = s0 ? tmp39070 : tmp39074;
  assign tmp39071 = ~(s1 ? tmp39072 : tmp39073);
  assign tmp39063 = s2 ? tmp39064 : tmp39071;
  assign tmp39058 = s3 ? tmp39059 : tmp39063;
  assign tmp39079 = l1 ? tmp37193 : tmp36682;
  assign tmp39078 = s0 ? tmp39079 : tmp36111;
  assign tmp39080 = ~(s0 ? tmp39060 : tmp39067);
  assign tmp39077 = s1 ? tmp39078 : tmp39080;
  assign tmp39082 = s0 ? tmp39060 : tmp36115;
  assign tmp39081 = ~(s1 ? tmp39082 : tmp36698);
  assign tmp39076 = s2 ? tmp39077 : tmp39081;
  assign tmp39086 = ~(l1 ? tmp37181 : tmp36263);
  assign tmp39085 = s0 ? tmp39070 : tmp39086;
  assign tmp39087 = s0 ? tmp37212 : tmp39070;
  assign tmp39084 = s1 ? tmp39085 : tmp39087;
  assign tmp39083 = s2 ? tmp36700 : tmp39084;
  assign tmp39075 = ~(s3 ? tmp39076 : tmp39083);
  assign tmp39057 = s4 ? tmp39058 : tmp39075;
  assign tmp39093 = s0 ? tmp39062 : tmp35793;
  assign tmp39094 = ~(l1 ? tmp35724 : tmp35717);
  assign tmp39092 = s1 ? tmp39093 : tmp39094;
  assign tmp39097 = l1 ? tmp37181 : tmp36263;
  assign tmp39096 = s0 ? tmp39097 : tmp36716;
  assign tmp39095 = ~(s1 ? tmp37221 : tmp39096);
  assign tmp39091 = s2 ? tmp39092 : tmp39095;
  assign tmp39100 = l1 ? tmp35833 : tmp36680;
  assign tmp39099 = s1 ? tmp39100 : tmp37137;
  assign tmp39098 = s2 ? tmp39099 : tmp37227;
  assign tmp39090 = s3 ? tmp39091 : tmp39098;
  assign tmp39104 = s0 ? tmp35971 : tmp39070;
  assign tmp39103 = s1 ? tmp39104 : tmp36726;
  assign tmp39102 = s2 ? tmp39103 : tmp37234;
  assign tmp39108 = l1 ? tmp36894 : tmp35882;
  assign tmp39107 = s0 ? tmp37151 : tmp39108;
  assign tmp39106 = s1 ? tmp39107 : tmp37309;
  assign tmp39105 = s2 ? tmp39106 : tmp35985;
  assign tmp39101 = s3 ? tmp39102 : tmp39105;
  assign tmp39089 = s4 ? tmp39090 : tmp39101;
  assign tmp39110 = s3 ? tmp39049 : tmp37316;
  assign tmp39111 = ~(s3 ? tmp37413 : tmp37323);
  assign tmp39109 = s4 ? tmp39110 : tmp39111;
  assign tmp39088 = ~(s5 ? tmp39089 : tmp39109);
  assign tmp39056 = s6 ? tmp39057 : tmp39088;
  assign tmp39055 = s7 ? tmp39033 : tmp39056;
  assign tmp39054 = s8 ? tmp39055 : tmp39039;
  assign tmp39052 = s9 ? tmp39053 : tmp39054;
  assign tmp39029 = s10 ? tmp39030 : tmp39052;
  assign tmp39119 = ~(s3 ? tmp39051 : tmp37323);
  assign tmp39118 = s4 ? tmp39110 : tmp39119;
  assign tmp39117 = ~(s5 ? tmp39089 : tmp39118);
  assign tmp39116 = s6 ? tmp39057 : tmp39117;
  assign tmp39115 = s7 ? tmp39033 : tmp39116;
  assign tmp39114 = s8 ? tmp39115 : tmp39039;
  assign tmp39113 = s9 ? tmp39053 : tmp39114;
  assign tmp39112 = s10 ? tmp39030 : tmp39113;
  assign tmp39028 = s11 ? tmp39029 : tmp39112;
  assign tmp39127 = s4 ? tmp38639 : tmp37704;
  assign tmp39126 = ~(s5 ? tmp37464 : tmp39127);
  assign tmp39125 = s6 ? tmp37430 : tmp39126;
  assign tmp39124 = s7 ? tmp35709 : tmp39125;
  assign tmp39131 = s4 ? tmp38650 : tmp37715;
  assign tmp39130 = ~(s5 ? tmp37534 : tmp39131);
  assign tmp39129 = s6 ? tmp37500 : tmp39130;
  assign tmp39128 = s7 ? tmp35709 : tmp39129;
  assign tmp39123 = s8 ? tmp39124 : tmp39128;
  assign tmp39132 = s8 ? tmp39128 : tmp37573;
  assign tmp39122 = s9 ? tmp39123 : tmp39132;
  assign tmp39137 = ~(s5 ? tmp37678 : tmp39127);
  assign tmp39136 = s6 ? tmp37646 : tmp39137;
  assign tmp39135 = s7 ? tmp35709 : tmp39136;
  assign tmp39134 = s8 ? tmp39135 : tmp35709;
  assign tmp39139 = s7 ? tmp39125 : tmp37706;
  assign tmp39140 = s7 ? tmp39129 : tmp39136;
  assign tmp39138 = s8 ? tmp39139 : tmp39140;
  assign tmp39133 = s9 ? tmp39134 : tmp39138;
  assign tmp39121 = s10 ? tmp39122 : tmp39133;
  assign tmp39144 = s7 ? tmp39125 : tmp37574;
  assign tmp39143 = s8 ? tmp39144 : tmp39140;
  assign tmp39142 = s9 ? tmp39134 : tmp39143;
  assign tmp39141 = s10 ? tmp39122 : tmp39142;
  assign tmp39120 = s11 ? tmp39121 : tmp39141;
  assign tmp39027 = s12 ? tmp39028 : tmp39120;
  assign tmp38822 = s13 ? tmp38823 : tmp39027;
  assign tmp38702 = s14 ? tmp38703 : tmp38822;
  assign tmp39156 = s3 ? tmp38160 : tmp38387;
  assign tmp39155 = s4 ? tmp39156 : tmp38399;
  assign tmp39154 = ~(s5 ? tmp38129 : tmp39155);
  assign tmp39153 = s6 ? tmp38097 : tmp39154;
  assign tmp39152 = s7 ? tmp35709 : tmp39153;
  assign tmp39151 = s8 ? tmp39152 : tmp38394;
  assign tmp39157 = s8 ? tmp38394 : tmp38235;
  assign tmp39150 = s9 ? tmp39151 : tmp39157;
  assign tmp39162 = ~(s5 ? tmp38332 : tmp39155);
  assign tmp39161 = s6 ? tmp38097 : tmp39162;
  assign tmp39160 = s7 ? tmp39161 : tmp38341;
  assign tmp39159 = s8 ? tmp39160 : tmp38487;
  assign tmp39158 = s9 ? tmp38474 : tmp39159;
  assign tmp39149 = s10 ? tmp39150 : tmp39158;
  assign tmp39166 = s7 ? tmp39153 : tmp38236;
  assign tmp39165 = s8 ? tmp39166 : tmp38487;
  assign tmp39164 = s9 ? tmp38474 : tmp39165;
  assign tmp39163 = s10 ? tmp39150 : tmp39164;
  assign tmp39148 = s11 ? tmp39149 : tmp39163;
  assign tmp39179 = ~(l1 ? tmp35833 : tmp35744);
  assign tmp39178 = s0 ? tmp35856 : tmp39179;
  assign tmp39177 = ~(s1 ? tmp39178 : tmp35827);
  assign tmp39176 = s2 ? tmp38161 : tmp39177;
  assign tmp39175 = s3 ? tmp39176 : tmp38387;
  assign tmp39174 = s4 ? tmp39175 : tmp38388;
  assign tmp39173 = ~(s5 ? tmp38207 : tmp39174);
  assign tmp39172 = s6 ? tmp38175 : tmp39173;
  assign tmp39171 = s7 ? tmp35709 : tmp39172;
  assign tmp39170 = s8 ? tmp38363 : tmp39171;
  assign tmp39169 = s9 ? tmp39170 : tmp39171;
  assign tmp39181 = s8 ? tmp39171 : tmp35709;
  assign tmp39189 = ~(l2 ? tmp35765 : tmp35716);
  assign tmp39188 = l1 ? tmp37181 : tmp39189;
  assign tmp39191 = l1 ? tmp37184 : tmp35779;
  assign tmp39190 = ~(s0 ? tmp36652 : tmp39191);
  assign tmp39187 = s1 ? tmp39188 : tmp39190;
  assign tmp39196 = ~(l2 ? tmp35727 : tmp35717);
  assign tmp39195 = ~(l1 ? tmp37190 : tmp39196);
  assign tmp39194 = s0 ? tmp37510 : tmp39195;
  assign tmp39198 = l1 ? tmp37190 : tmp39196;
  assign tmp39197 = ~(s0 ? tmp38186 : tmp39198);
  assign tmp39193 = s1 ? tmp39194 : tmp39197;
  assign tmp39201 = ~(l1 ? tmp37181 : tmp39189);
  assign tmp39200 = s0 ? tmp39198 : tmp39201;
  assign tmp39199 = ~(s1 ? tmp38189 : tmp39200);
  assign tmp39192 = s2 ? tmp39193 : tmp39199;
  assign tmp39186 = s3 ? tmp39187 : tmp39192;
  assign tmp39206 = l1 ? tmp37193 : tmp35779;
  assign tmp39205 = s0 ? tmp39206 : tmp36456;
  assign tmp39207 = ~(s0 ? tmp39188 : tmp39195);
  assign tmp39204 = s1 ? tmp39205 : tmp39207;
  assign tmp39209 = s0 ? tmp39188 : tmp36115;
  assign tmp39208 = ~(s1 ? tmp39209 : tmp37865);
  assign tmp39203 = s2 ? tmp39204 : tmp39208;
  assign tmp39214 = l2 ? tmp35727 : tmp35717;
  assign tmp39213 = ~(l1 ? tmp37181 : tmp39214);
  assign tmp39212 = s0 ? tmp39198 : tmp39213;
  assign tmp39215 = s0 ? tmp38127 : tmp39198;
  assign tmp39211 = s1 ? tmp39212 : tmp39215;
  assign tmp39210 = s2 ? tmp38201 : tmp39211;
  assign tmp39202 = ~(s3 ? tmp39203 : tmp39210);
  assign tmp39185 = s4 ? tmp39186 : tmp39202;
  assign tmp39221 = s0 ? tmp39191 : tmp36474;
  assign tmp39220 = s1 ? tmp39221 : tmp37539;
  assign tmp39223 = l1 ? tmp37181 : tmp35914;
  assign tmp39225 = l1 ? tmp37181 : tmp39214;
  assign tmp39224 = s0 ? tmp39225 : tmp37544;
  assign tmp39222 = ~(s1 ? tmp39223 : tmp39224);
  assign tmp39219 = s2 ? tmp39220 : tmp39222;
  assign tmp39228 = l1 ? tmp35786 : tmp39196;
  assign tmp39227 = s1 ? tmp37160 : tmp39228;
  assign tmp39230 = s0 ? tmp39198 : tmp38127;
  assign tmp39229 = s1 ? tmp38143 : tmp39230;
  assign tmp39226 = s2 ? tmp39227 : tmp39229;
  assign tmp39218 = s3 ? tmp39219 : tmp39226;
  assign tmp39234 = s0 ? tmp36883 : tmp39198;
  assign tmp39233 = s1 ? tmp39234 : tmp37893;
  assign tmp39235 = ~(l1 ? tmp35724 : tmp35914);
  assign tmp39232 = s2 ? tmp39233 : tmp39235;
  assign tmp39239 = l1 ? tmp35833 : tmp37850;
  assign tmp39240 = l1 ? tmp36894 : tmp36854;
  assign tmp39238 = s0 ? tmp39239 : tmp39240;
  assign tmp39237 = s1 ? tmp39238 : tmp38456;
  assign tmp39236 = s2 ? tmp39237 : tmp36895;
  assign tmp39231 = s3 ? tmp39232 : tmp39236;
  assign tmp39217 = s4 ? tmp39218 : tmp39231;
  assign tmp39245 = s0 ? tmp39228 : tmp35850;
  assign tmp39244 = s1 ? tmp39245 : tmp38163;
  assign tmp39246 = ~(s1 ? tmp39178 : tmp35736);
  assign tmp39243 = s2 ? tmp39244 : tmp39246;
  assign tmp39242 = s3 ? tmp39243 : tmp38464;
  assign tmp39249 = l1 ? tmp35714 : tmp35914;
  assign tmp39248 = s2 ? tmp38390 : tmp39249;
  assign tmp39247 = ~(s3 ? tmp39248 : tmp38472);
  assign tmp39241 = s4 ? tmp39242 : tmp39247;
  assign tmp39216 = ~(s5 ? tmp39217 : tmp39241);
  assign tmp39184 = s6 ? tmp39185 : tmp39216;
  assign tmp39183 = s7 ? tmp38484 : tmp39184;
  assign tmp39252 = s4 ? tmp39175 : tmp38399;
  assign tmp39251 = ~(s5 ? tmp38207 : tmp39252);
  assign tmp39250 = s6 ? tmp38175 : tmp39251;
  assign tmp39182 = s8 ? tmp39183 : tmp39250;
  assign tmp39180 = s9 ? tmp39181 : tmp39182;
  assign tmp39168 = s10 ? tmp39169 : tmp39180;
  assign tmp39261 = s1 ? tmp38393 : tmp38471;
  assign tmp39260 = ~(s3 ? tmp39248 : tmp39261);
  assign tmp39259 = s4 ? tmp39242 : tmp39260;
  assign tmp39258 = ~(s5 ? tmp39217 : tmp39259);
  assign tmp39257 = s6 ? tmp39185 : tmp39258;
  assign tmp39256 = s7 ? tmp38364 : tmp39257;
  assign tmp39255 = s8 ? tmp39256 : tmp39172;
  assign tmp39254 = s9 ? tmp39181 : tmp39255;
  assign tmp39253 = s10 ? tmp39169 : tmp39254;
  assign tmp39167 = s11 ? tmp39168 : tmp39253;
  assign tmp39147 = s12 ? tmp39148 : tmp39167;
  assign tmp39146 = s13 ? tmp39147 : tmp38492;
  assign tmp39145 = s14 ? tmp37725 : tmp39146;
  assign tmp38701 = s15 ? tmp38702 : tmp39145;
  assign tmp35700 = s16 ? tmp35701 : tmp38701;
  assign tmp39269 = s8 ? tmp38708 : tmp36081;
  assign tmp39268 = s9 ? tmp38707 : tmp39269;
  assign tmp39272 = s7 ? tmp38734 : tmp36171;
  assign tmp39271 = s8 ? tmp36219 : tmp39272;
  assign tmp39270 = s9 ? tmp36169 : tmp39271;
  assign tmp39267 = s10 ? tmp39268 : tmp39270;
  assign tmp39276 = s7 ? tmp38709 : tmp36171;
  assign tmp39275 = s8 ? tmp36230 : tmp39276;
  assign tmp39274 = s9 ? tmp36169 : tmp39275;
  assign tmp39273 = s10 ? tmp39268 : tmp39274;
  assign tmp39266 = s11 ? tmp39267 : tmp39273;
  assign tmp39281 = s8 ? tmp38756 : tmp36565;
  assign tmp39280 = s9 ? tmp38755 : tmp39281;
  assign tmp39284 = s7 ? tmp38815 : tmp36613;
  assign tmp39283 = s8 ? tmp36625 : tmp39284;
  assign tmp39282 = s9 ? tmp36611 : tmp39283;
  assign tmp39279 = s10 ? tmp39280 : tmp39282;
  assign tmp39288 = s7 ? tmp38757 : tmp36613;
  assign tmp39287 = s8 ? tmp36633 : tmp39288;
  assign tmp39286 = s9 ? tmp36611 : tmp39287;
  assign tmp39285 = s10 ? tmp39280 : tmp39286;
  assign tmp39278 = s11 ? tmp39279 : tmp39285;
  assign tmp39277 = s12 ? tmp36232 : tmp39278;
  assign tmp39265 = s13 ? tmp39266 : tmp39277;
  assign tmp39294 = s8 ? tmp38827 : tmp36743;
  assign tmp39293 = s9 ? tmp38827 : tmp39294;
  assign tmp39297 = s7 ? tmp38943 : tmp36672;
  assign tmp39296 = s8 ? tmp36807 : tmp39297;
  assign tmp39295 = s9 ? tmp36805 : tmp39296;
  assign tmp39292 = s10 ? tmp39293 : tmp39295;
  assign tmp39301 = s7 ? tmp38828 : tmp36672;
  assign tmp39300 = s8 ? tmp36816 : tmp39301;
  assign tmp39299 = s9 ? tmp36805 : tmp39300;
  assign tmp39298 = s10 ? tmp39293 : tmp39299;
  assign tmp39291 = s11 ? tmp39292 : tmp39298;
  assign tmp39306 = s7 ? tmp35709 : tmp37006;
  assign tmp39305 = s8 ? tmp38955 : tmp39306;
  assign tmp39304 = s9 ? tmp38955 : tmp39305;
  assign tmp39308 = s7 ? tmp39019 : tmp36916;
  assign tmp39307 = s9 ? tmp36997 : tmp39308;
  assign tmp39303 = s10 ? tmp39304 : tmp39307;
  assign tmp39311 = s7 ? tmp38956 : tmp36916;
  assign tmp39310 = s9 ? tmp36997 : tmp39311;
  assign tmp39309 = s10 ? tmp39304 : tmp39310;
  assign tmp39302 = s11 ? tmp39303 : tmp39309;
  assign tmp39290 = s12 ? tmp39291 : tmp39302;
  assign tmp39316 = s8 ? tmp37090 : tmp39044;
  assign tmp39317 = s8 ? tmp39044 : tmp37251;
  assign tmp39315 = s9 ? tmp39316 : tmp39317;
  assign tmp39323 = s4 ? tmp39048 : tmp37412;
  assign tmp39322 = ~(s5 ? tmp37214 : tmp39323);
  assign tmp39321 = s6 ? tmp37177 : tmp39322;
  assign tmp39320 = s7 ? tmp39321 : tmp37414;
  assign tmp39319 = s8 ? tmp37397 : tmp39320;
  assign tmp39318 = s9 ? tmp37326 : tmp39319;
  assign tmp39314 = s10 ? tmp39315 : tmp39318;
  assign tmp39327 = s7 ? tmp39045 : tmp37328;
  assign tmp39326 = s8 ? tmp37422 : tmp39327;
  assign tmp39325 = s9 ? tmp37326 : tmp39326;
  assign tmp39324 = s10 ? tmp39315 : tmp39325;
  assign tmp39313 = s11 ? tmp39314 : tmp39324;
  assign tmp39312 = s12 ? tmp39313 : tmp37424;
  assign tmp39289 = s13 ? tmp39290 : tmp39312;
  assign tmp39264 = s14 ? tmp39265 : tmp39289;
  assign tmp39334 = s8 ? tmp39171 : tmp38401;
  assign tmp39333 = s9 ? tmp39170 : tmp39334;
  assign tmp39337 = s7 ? tmp39250 : tmp38476;
  assign tmp39336 = s8 ? tmp38483 : tmp39337;
  assign tmp39335 = s9 ? tmp38474 : tmp39336;
  assign tmp39332 = s10 ? tmp39333 : tmp39335;
  assign tmp39341 = s7 ? tmp39172 : tmp38476;
  assign tmp39340 = s8 ? tmp38491 : tmp39341;
  assign tmp39339 = s9 ? tmp38474 : tmp39340;
  assign tmp39338 = s10 ? tmp39333 : tmp39339;
  assign tmp39331 = s11 ? tmp39332 : tmp39338;
  assign tmp39330 = s12 ? tmp38091 : tmp39331;
  assign tmp39329 = s13 ? tmp39330 : tmp38492;
  assign tmp39328 = s14 ? tmp37725 : tmp39329;
  assign tmp39263 = s15 ? tmp39264 : tmp39328;
  assign tmp39348 = s9 ? tmp39316 : tmp39044;
  assign tmp39350 = s8 ? tmp39044 : tmp35709;
  assign tmp39352 = s7 ? tmp37398 : tmp39056;
  assign tmp39351 = s8 ? tmp39352 : tmp39321;
  assign tmp39349 = s9 ? tmp39350 : tmp39351;
  assign tmp39347 = s10 ? tmp39348 : tmp39349;
  assign tmp39356 = s7 ? tmp37091 : tmp39116;
  assign tmp39355 = s8 ? tmp39356 : tmp39045;
  assign tmp39354 = s9 ? tmp39350 : tmp39355;
  assign tmp39353 = s10 ? tmp39348 : tmp39354;
  assign tmp39346 = s11 ? tmp39347 : tmp39353;
  assign tmp39345 = s12 ? tmp39346 : tmp37424;
  assign tmp39344 = s13 ? tmp38823 : tmp39345;
  assign tmp39343 = s14 ? tmp38703 : tmp39344;
  assign tmp39359 = s12 ? tmp38091 : tmp39167;
  assign tmp39358 = s13 ? tmp39359 : tmp38492;
  assign tmp39357 = s14 ? tmp37725 : tmp39358;
  assign tmp39342 = s15 ? tmp39343 : tmp39357;
  assign tmp39262 = s16 ? tmp39263 : tmp39342;
  assign tmp35699 = s17 ? tmp35700 : tmp39262;
  assign s2n = tmp35699;

  assign tmp39376 = l3 ? 1 : 0;
  assign tmp39375 = l2 ? tmp39376 : 1;
  assign tmp39379 = l4 ? 1 : 0;
  assign tmp39378 = l3 ? tmp39379 : 1;
  assign tmp39381 = ~(l4 ? 1 : 0);
  assign tmp39380 = ~(l3 ? tmp39379 : tmp39381);
  assign tmp39377 = ~(l2 ? tmp39378 : tmp39380);
  assign tmp39374 = l1 ? tmp39375 : tmp39377;
  assign tmp39384 = l2 ? 1 : tmp39381;
  assign tmp39386 = ~(l3 ? tmp39379 : 0);
  assign tmp39385 = l2 ? 1 : tmp39386;
  assign tmp39383 = l1 ? tmp39384 : tmp39385;
  assign tmp39389 = ~(l3 ? 1 : tmp39381);
  assign tmp39388 = ~(l2 ? tmp39378 : tmp39389);
  assign tmp39387 = ~(l1 ? tmp39375 : tmp39388);
  assign tmp39382 = ~(s0 ? tmp39383 : tmp39387);
  assign tmp39373 = s1 ? tmp39374 : tmp39382;
  assign tmp39394 = ~(l2 ? 1 : tmp39380);
  assign tmp39393 = ~(l1 ? tmp39375 : tmp39394);
  assign tmp39392 = s0 ? tmp39383 : tmp39393;
  assign tmp39398 = ~(l3 ? 1 : tmp39379);
  assign tmp39397 = l2 ? 1 : tmp39398;
  assign tmp39396 = l1 ? tmp39397 : tmp39385;
  assign tmp39395 = s0 ? tmp39396 : tmp39393;
  assign tmp39391 = s1 ? tmp39392 : tmp39395;
  assign tmp39403 = l3 ? 1 : tmp39381;
  assign tmp39402 = l2 ? tmp39403 : 1;
  assign tmp39404 = ~(l2 ? tmp39379 : 0);
  assign tmp39401 = ~(l1 ? tmp39402 : tmp39404);
  assign tmp39400 = s0 ? tmp39396 : tmp39401;
  assign tmp39406 = l1 ? tmp39375 : tmp39394;
  assign tmp39408 = l2 ? tmp39378 : 0;
  assign tmp39409 = l2 ? 1 : tmp39380;
  assign tmp39407 = ~(l1 ? tmp39408 : tmp39409);
  assign tmp39405 = ~(s0 ? tmp39406 : tmp39407);
  assign tmp39399 = s1 ? tmp39400 : tmp39405;
  assign tmp39390 = ~(s2 ? tmp39391 : tmp39399);
  assign tmp39372 = s3 ? tmp39373 : tmp39390;
  assign tmp39414 = l1 ? tmp39375 : tmp39388;
  assign tmp39415 = ~(l1 ? tmp39384 : tmp39385);
  assign tmp39413 = s0 ? tmp39414 : tmp39415;
  assign tmp39417 = l1 ? tmp39408 : tmp39409;
  assign tmp39416 = ~(s0 ? tmp39417 : tmp39393);
  assign tmp39412 = s1 ? tmp39413 : tmp39416;
  assign tmp39420 = ~(l2 ? 1 : tmp39386);
  assign tmp39419 = s0 ? tmp39374 : tmp39420;
  assign tmp39423 = ~(l2 ? tmp39378 : 0);
  assign tmp39422 = l1 ? tmp39402 : tmp39423;
  assign tmp39424 = ~(l1 ? tmp39402 : tmp39385);
  assign tmp39421 = s0 ? tmp39422 : tmp39424;
  assign tmp39418 = s1 ? tmp39419 : tmp39421;
  assign tmp39411 = s2 ? tmp39412 : tmp39418;
  assign tmp39430 = l3 ? 1 : tmp39379;
  assign tmp39429 = l2 ? tmp39430 : 1;
  assign tmp39428 = l1 ? tmp39385 : tmp39429;
  assign tmp39427 = s0 ? tmp39428 : tmp39415;
  assign tmp39432 = l1 ? tmp39402 : tmp39385;
  assign tmp39434 = l2 ? tmp39378 : tmp39379;
  assign tmp39435 = l2 ? 1 : tmp39430;
  assign tmp39433 = l1 ? tmp39434 : tmp39435;
  assign tmp39431 = ~(s0 ? tmp39432 : tmp39433);
  assign tmp39426 = s1 ? tmp39427 : tmp39431;
  assign tmp39440 = l3 ? tmp39379 : 0;
  assign tmp39439 = l2 ? tmp39440 : tmp39378;
  assign tmp39438 = l1 ? tmp39429 : tmp39439;
  assign tmp39437 = s0 ? tmp39438 : tmp39406;
  assign tmp39436 = s1 ? tmp39406 : tmp39437;
  assign tmp39425 = s2 ? tmp39426 : tmp39436;
  assign tmp39410 = s3 ? tmp39411 : tmp39425;
  assign tmp39371 = s4 ? tmp39372 : tmp39410;
  assign tmp39446 = s0 ? tmp39414 : tmp39420;
  assign tmp39448 = l1 ? 1 : tmp39386;
  assign tmp39447 = ~(s0 ? tmp39448 : tmp39383);
  assign tmp39445 = s1 ? tmp39446 : tmp39447;
  assign tmp39450 = s0 ? tmp39448 : tmp39387;
  assign tmp39452 = ~(l1 ? 1 : tmp39385);
  assign tmp39451 = ~(s0 ? tmp39406 : tmp39452);
  assign tmp39449 = ~(s1 ? tmp39450 : tmp39451);
  assign tmp39444 = s2 ? tmp39445 : tmp39449;
  assign tmp39457 = ~(l2 ? tmp39379 : tmp39440);
  assign tmp39456 = l1 ? tmp39402 : tmp39457;
  assign tmp39460 = l3 ? tmp39379 : tmp39381;
  assign tmp39459 = l2 ? 1 : tmp39460;
  assign tmp39458 = l1 ? tmp39459 : tmp39385;
  assign tmp39455 = s0 ? tmp39456 : tmp39458;
  assign tmp39462 = ~(l1 ? tmp39429 : tmp39394);
  assign tmp39461 = s0 ? tmp39456 : tmp39462;
  assign tmp39454 = s1 ? tmp39455 : tmp39461;
  assign tmp39465 = l1 ? 1 : tmp39378;
  assign tmp39464 = s0 ? tmp39438 : tmp39465;
  assign tmp39467 = l1 ? tmp39408 : tmp39435;
  assign tmp39469 = l2 ? tmp39378 : tmp39440;
  assign tmp39468 = l1 ? tmp39469 : tmp39435;
  assign tmp39466 = ~(s0 ? tmp39467 : tmp39468);
  assign tmp39463 = ~(s1 ? tmp39464 : tmp39466);
  assign tmp39453 = ~(s2 ? tmp39454 : tmp39463);
  assign tmp39443 = s3 ? tmp39444 : tmp39453;
  assign tmp39475 = l2 ? tmp39379 : tmp39378;
  assign tmp39474 = l1 ? 1 : tmp39475;
  assign tmp39473 = s0 ? tmp39474 : tmp39374;
  assign tmp39478 = ~(l2 ? tmp39440 : 0);
  assign tmp39477 = l1 ? tmp39402 : tmp39478;
  assign tmp39480 = l2 ? 1 : tmp39403;
  assign tmp39479 = ~(l1 ? tmp39480 : 1);
  assign tmp39476 = s0 ? tmp39477 : tmp39479;
  assign tmp39472 = s1 ? tmp39473 : tmp39476;
  assign tmp39483 = l1 ? tmp39385 : 1;
  assign tmp39484 = ~(l1 ? tmp39403 : tmp39402);
  assign tmp39482 = s0 ? tmp39483 : tmp39484;
  assign tmp39486 = l1 ? tmp39384 : tmp39435;
  assign tmp39487 = ~(l1 ? tmp39385 : 1);
  assign tmp39485 = ~(s0 ? tmp39486 : tmp39487);
  assign tmp39481 = s1 ? tmp39482 : tmp39485;
  assign tmp39471 = s2 ? tmp39472 : tmp39481;
  assign tmp39491 = l1 ? tmp39480 : tmp39435;
  assign tmp39493 = l2 ? tmp39376 : tmp39460;
  assign tmp39492 = ~(l1 ? tmp39375 : tmp39493);
  assign tmp39490 = s0 ? tmp39491 : tmp39492;
  assign tmp39495 = l1 ? tmp39403 : tmp39402;
  assign tmp39497 = l2 ? tmp39379 : tmp39460;
  assign tmp39496 = ~(l1 ? tmp39429 : tmp39497);
  assign tmp39494 = s0 ? tmp39495 : tmp39496;
  assign tmp39489 = s1 ? tmp39490 : tmp39494;
  assign tmp39501 = l2 ? tmp39378 : 1;
  assign tmp39500 = l1 ? tmp39501 : 1;
  assign tmp39499 = s0 ? tmp39500 : tmp39465;
  assign tmp39502 = s0 ? tmp39433 : tmp39465;
  assign tmp39498 = s1 ? tmp39499 : tmp39502;
  assign tmp39488 = ~(s2 ? tmp39489 : tmp39498);
  assign tmp39470 = s3 ? tmp39471 : tmp39488;
  assign tmp39442 = s4 ? tmp39443 : tmp39470;
  assign tmp39508 = l1 ? tmp39429 : tmp39394;
  assign tmp39509 = ~(l1 ? tmp39378 : 1);
  assign tmp39507 = s0 ? tmp39508 : tmp39509;
  assign tmp39511 = l1 ? 1 : tmp39501;
  assign tmp39513 = l2 ? 1 : tmp39378;
  assign tmp39512 = l1 ? tmp39513 : 1;
  assign tmp39510 = ~(s0 ? tmp39511 : tmp39512);
  assign tmp39506 = s1 ? tmp39507 : tmp39510;
  assign tmp39516 = l1 ? 1 : tmp39402;
  assign tmp39518 = ~(l2 ? tmp39379 : tmp39389);
  assign tmp39517 = ~(l1 ? tmp39429 : tmp39518);
  assign tmp39515 = s0 ? tmp39516 : tmp39517;
  assign tmp39520 = l1 ? tmp39480 : 1;
  assign tmp39521 = ~(l1 ? tmp39429 : 1);
  assign tmp39519 = s0 ? tmp39520 : tmp39521;
  assign tmp39514 = ~(s1 ? tmp39515 : tmp39519);
  assign tmp39505 = s2 ? tmp39506 : tmp39514;
  assign tmp39524 = s0 ? tmp39480 : tmp39435;
  assign tmp39527 = l2 ? 1 : tmp39379;
  assign tmp39526 = l1 ? tmp39435 : tmp39527;
  assign tmp39528 = ~(l1 ? 1 : tmp39378);
  assign tmp39525 = s0 ? tmp39526 : tmp39528;
  assign tmp39523 = s1 ? tmp39524 : tmp39525;
  assign tmp39532 = l2 ? tmp39430 : tmp39378;
  assign tmp39531 = l1 ? 1 : tmp39532;
  assign tmp39530 = s0 ? tmp39512 : tmp39531;
  assign tmp39534 = l1 ? tmp39378 : tmp39429;
  assign tmp39535 = ~(l1 ? tmp39480 : tmp39435);
  assign tmp39533 = s0 ? tmp39534 : tmp39535;
  assign tmp39529 = ~(s1 ? tmp39530 : tmp39533);
  assign tmp39522 = ~(s2 ? tmp39523 : tmp39529);
  assign tmp39504 = s3 ? tmp39505 : tmp39522;
  assign tmp39541 = l2 ? 1 : tmp39376;
  assign tmp39540 = l1 ? tmp39480 : tmp39541;
  assign tmp39539 = s0 ? tmp39540 : tmp39521;
  assign tmp39543 = l1 ? tmp39532 : 1;
  assign tmp39542 = ~(s0 ? tmp39543 : tmp39438);
  assign tmp39538 = s1 ? tmp39539 : tmp39542;
  assign tmp39547 = l2 ? 1 : tmp39440;
  assign tmp39546 = l1 ? tmp39547 : tmp39435;
  assign tmp39545 = s0 ? tmp39511 : tmp39546;
  assign tmp39549 = l1 ? tmp39429 : 1;
  assign tmp39550 = ~(l2 ? 1 : tmp39403);
  assign tmp39548 = ~(s0 ? tmp39549 : tmp39550);
  assign tmp39544 = s1 ? tmp39545 : tmp39548;
  assign tmp39537 = s2 ? tmp39538 : tmp39544;
  assign tmp39554 = ~(l1 ? tmp39429 : tmp39378);
  assign tmp39553 = s0 ? tmp39516 : tmp39554;
  assign tmp39556 = ~(l1 ? tmp39469 : tmp39435);
  assign tmp39555 = ~(s0 ? tmp39512 : tmp39556);
  assign tmp39552 = s1 ? tmp39553 : tmp39555;
  assign tmp39559 = ~(l1 ? tmp39480 : tmp39541);
  assign tmp39558 = s0 ? tmp39534 : tmp39559;
  assign tmp39561 = ~(l1 ? tmp39532 : 1);
  assign tmp39560 = ~(s0 ? tmp39526 : tmp39561);
  assign tmp39557 = ~(s1 ? tmp39558 : tmp39560);
  assign tmp39551 = s2 ? tmp39552 : tmp39557;
  assign tmp39536 = ~(s3 ? tmp39537 : tmp39551);
  assign tmp39503 = s4 ? tmp39504 : tmp39536;
  assign tmp39441 = s5 ? tmp39442 : tmp39503;
  assign tmp39370 = s6 ? tmp39371 : tmp39441;
  assign tmp39567 = ~(l2 ? tmp39440 : tmp39378);
  assign tmp39566 = l1 ? tmp39378 : tmp39567;
  assign tmp39569 = l1 ? tmp39384 : tmp39375;
  assign tmp39570 = ~(l1 ? tmp39527 : tmp39567);
  assign tmp39568 = ~(s0 ? tmp39569 : tmp39570);
  assign tmp39565 = s1 ? tmp39566 : tmp39568;
  assign tmp39575 = l2 ? tmp39376 : tmp39381;
  assign tmp39574 = l1 ? tmp39575 : 1;
  assign tmp39577 = l2 ? tmp39460 : tmp39379;
  assign tmp39578 = ~(l2 ? tmp39430 : tmp39378);
  assign tmp39576 = ~(l1 ? tmp39577 : tmp39578);
  assign tmp39573 = s0 ? tmp39574 : tmp39576;
  assign tmp39580 = l1 ? tmp39575 : tmp39375;
  assign tmp39579 = s0 ? tmp39580 : tmp39576;
  assign tmp39572 = s1 ? tmp39573 : tmp39579;
  assign tmp39583 = ~(l1 ? tmp39402 : tmp39457);
  assign tmp39582 = s0 ? tmp39580 : tmp39583;
  assign tmp39585 = l1 ? tmp39577 : tmp39578;
  assign tmp39587 = l2 ? tmp39430 : tmp39381;
  assign tmp39588 = l2 ? tmp39376 : tmp39378;
  assign tmp39586 = ~(l1 ? tmp39587 : tmp39588);
  assign tmp39584 = ~(s0 ? tmp39585 : tmp39586);
  assign tmp39581 = s1 ? tmp39582 : tmp39584;
  assign tmp39571 = ~(s2 ? tmp39572 : tmp39581);
  assign tmp39564 = s3 ? tmp39565 : tmp39571;
  assign tmp39593 = l1 ? 1 : tmp39567;
  assign tmp39594 = ~(l1 ? tmp39384 : 1);
  assign tmp39592 = s0 ? tmp39593 : tmp39594;
  assign tmp39596 = l1 ? tmp39587 : tmp39588;
  assign tmp39595 = ~(s0 ? tmp39596 : tmp39576);
  assign tmp39591 = s1 ? tmp39592 : tmp39595;
  assign tmp39598 = s0 ? tmp39566 : tmp39487;
  assign tmp39597 = s1 ? tmp39598 : tmp39477;
  assign tmp39590 = s2 ? tmp39591 : tmp39597;
  assign tmp39600 = s1 ? tmp39569 : tmp39531;
  assign tmp39604 = l2 ? tmp39378 : tmp39430;
  assign tmp39603 = l1 ? tmp39434 : tmp39604;
  assign tmp39602 = s0 ? tmp39603 : tmp39585;
  assign tmp39601 = ~(s1 ? tmp39585 : tmp39602);
  assign tmp39599 = ~(s2 ? tmp39600 : tmp39601);
  assign tmp39589 = s3 ? tmp39590 : tmp39599;
  assign tmp39563 = s4 ? tmp39564 : tmp39589;
  assign tmp39611 = l1 ? tmp39527 : tmp39567;
  assign tmp39610 = s0 ? tmp39611 : tmp39487;
  assign tmp39612 = ~(l1 ? tmp39575 : 1);
  assign tmp39609 = s1 ? tmp39610 : tmp39612;
  assign tmp39616 = ~(l3 ? 1 : 0);
  assign tmp39615 = ~(l2 ? tmp39379 : tmp39616);
  assign tmp39614 = l1 ? tmp39527 : tmp39615;
  assign tmp39617 = s0 ? tmp39585 : 0;
  assign tmp39613 = s1 ? tmp39614 : tmp39617;
  assign tmp39608 = s2 ? tmp39609 : tmp39613;
  assign tmp39621 = l2 ? tmp39376 : tmp39403;
  assign tmp39620 = l1 ? tmp39621 : tmp39375;
  assign tmp39623 = ~(l2 ? tmp39430 : tmp39616);
  assign tmp39622 = ~(l1 ? tmp39434 : tmp39623);
  assign tmp39619 = s1 ? tmp39620 : tmp39622;
  assign tmp39626 = l1 ? tmp39434 : tmp39501;
  assign tmp39625 = s0 ? tmp39603 : tmp39626;
  assign tmp39628 = l1 ? tmp39587 : tmp39532;
  assign tmp39630 = l2 ? tmp39430 : tmp39403;
  assign tmp39629 = l1 ? tmp39630 : tmp39532;
  assign tmp39627 = ~(s0 ? tmp39628 : tmp39629);
  assign tmp39624 = ~(s1 ? tmp39625 : tmp39627);
  assign tmp39618 = ~(s2 ? tmp39619 : tmp39624);
  assign tmp39607 = s3 ? tmp39608 : tmp39618;
  assign tmp39635 = l1 ? tmp39378 : tmp39604;
  assign tmp39637 = ~(l2 ? tmp39440 : tmp39616);
  assign tmp39636 = l1 ? tmp39577 : tmp39637;
  assign tmp39634 = s0 ? tmp39635 : tmp39636;
  assign tmp39639 = ~(l1 ? tmp39480 : tmp39375);
  assign tmp39638 = s0 ? tmp39477 : tmp39639;
  assign tmp39633 = s1 ? tmp39634 : tmp39638;
  assign tmp39642 = l1 ? tmp39575 : tmp39429;
  assign tmp39641 = ~(s0 ? tmp39642 : tmp39487);
  assign tmp39640 = s1 ? tmp39483 : tmp39641;
  assign tmp39632 = s2 ? tmp39633 : tmp39640;
  assign tmp39646 = l1 ? tmp39630 : tmp39429;
  assign tmp39647 = ~(l1 ? tmp39378 : tmp39541);
  assign tmp39645 = s0 ? tmp39646 : tmp39647;
  assign tmp39649 = l2 ? tmp39378 : tmp39376;
  assign tmp39648 = ~(l1 ? tmp39434 : tmp39649);
  assign tmp39644 = s1 ? tmp39645 : tmp39648;
  assign tmp39651 = l1 ? 1 : tmp39513;
  assign tmp39650 = s1 ? tmp39651 : tmp39531;
  assign tmp39643 = ~(s2 ? tmp39644 : tmp39650);
  assign tmp39631 = s3 ? tmp39632 : tmp39643;
  assign tmp39606 = s4 ? tmp39607 : tmp39631;
  assign tmp39657 = l1 ? tmp39434 : tmp39623;
  assign tmp39656 = s0 ? tmp39657 : 0;
  assign tmp39658 = ~(l1 ? tmp39429 : tmp39375);
  assign tmp39655 = s1 ? tmp39656 : tmp39658;
  assign tmp39660 = l1 ? 1 : tmp39518;
  assign tmp39661 = ~(l1 ? tmp39630 : 1);
  assign tmp39659 = s1 ? tmp39660 : tmp39661;
  assign tmp39654 = s2 ? tmp39655 : tmp39659;
  assign tmp39664 = ~(l1 ? tmp39527 : tmp39501);
  assign tmp39663 = s1 ? tmp39651 : tmp39664;
  assign tmp39666 = l1 ? tmp39378 : tmp39435;
  assign tmp39667 = ~(l1 ? tmp39630 : tmp39429);
  assign tmp39665 = ~(s1 ? tmp39666 : tmp39667);
  assign tmp39662 = ~(s2 ? tmp39663 : tmp39665);
  assign tmp39653 = s3 ? tmp39654 : tmp39662;
  assign tmp39671 = l1 ? tmp39527 : tmp39435;
  assign tmp39670 = s1 ? tmp39671 : tmp39603;
  assign tmp39669 = s2 ? tmp39670 : tmp39667;
  assign tmp39673 = l1 ? tmp39527 : tmp39604;
  assign tmp39674 = ~(l1 ? tmp39630 : tmp39532);
  assign tmp39672 = s1 ? tmp39673 : tmp39674;
  assign tmp39668 = s3 ? tmp39669 : tmp39672;
  assign tmp39652 = s4 ? tmp39653 : tmp39668;
  assign tmp39605 = s5 ? tmp39606 : tmp39652;
  assign tmp39562 = s6 ? tmp39563 : tmp39605;
  assign tmp39369 = s7 ? tmp39370 : tmp39562;
  assign tmp39681 = l2 ? tmp39460 : tmp39378;
  assign tmp39680 = l1 ? tmp39681 : tmp39567;
  assign tmp39684 = l2 ? tmp39403 : tmp39379;
  assign tmp39683 = ~(l1 ? tmp39684 : tmp39567);
  assign tmp39682 = ~(s0 ? tmp39569 : tmp39683);
  assign tmp39679 = s1 ? tmp39680 : tmp39682;
  assign tmp39688 = l1 ? tmp39587 : tmp39402;
  assign tmp39690 = ~(l2 ? tmp39376 : tmp39378);
  assign tmp39689 = ~(l1 ? tmp39577 : tmp39690);
  assign tmp39687 = s0 ? tmp39688 : tmp39689;
  assign tmp39692 = l1 ? tmp39587 : tmp39375;
  assign tmp39691 = s0 ? tmp39692 : tmp39689;
  assign tmp39686 = s1 ? tmp39687 : tmp39691;
  assign tmp39695 = ~(l1 ? tmp39402 : tmp39386);
  assign tmp39694 = s0 ? tmp39692 : tmp39695;
  assign tmp39697 = l1 ? tmp39577 : tmp39690;
  assign tmp39696 = ~(s0 ? tmp39697 : tmp39586);
  assign tmp39693 = s1 ? tmp39694 : tmp39696;
  assign tmp39685 = ~(s2 ? tmp39686 : tmp39693);
  assign tmp39678 = s3 ? tmp39679 : tmp39685;
  assign tmp39702 = l1 ? tmp39402 : tmp39567;
  assign tmp39701 = s0 ? tmp39702 : tmp39594;
  assign tmp39703 = ~(s0 ? tmp39596 : tmp39689);
  assign tmp39700 = s1 ? tmp39701 : tmp39703;
  assign tmp39705 = s0 ? tmp39680 : tmp39487;
  assign tmp39704 = s1 ? tmp39705 : tmp39477;
  assign tmp39699 = s2 ? tmp39700 : tmp39704;
  assign tmp39708 = s0 ? tmp39603 : tmp39697;
  assign tmp39707 = ~(s1 ? tmp39697 : tmp39708);
  assign tmp39706 = ~(s2 ? tmp39600 : tmp39707);
  assign tmp39698 = s3 ? tmp39699 : tmp39706;
  assign tmp39677 = s4 ? tmp39678 : tmp39698;
  assign tmp39715 = l1 ? tmp39684 : tmp39567;
  assign tmp39714 = s0 ? tmp39715 : tmp39487;
  assign tmp39716 = ~(l1 ? tmp39587 : tmp39402);
  assign tmp39713 = s1 ? tmp39714 : tmp39716;
  assign tmp39718 = l1 ? tmp39684 : tmp39637;
  assign tmp39720 = ~(l1 ? 1 : tmp39402);
  assign tmp39719 = s0 ? tmp39697 : tmp39720;
  assign tmp39717 = s1 ? tmp39718 : tmp39719;
  assign tmp39712 = s2 ? tmp39713 : tmp39717;
  assign tmp39723 = l1 ? tmp39630 : tmp39375;
  assign tmp39725 = ~(l2 ? tmp39376 : tmp39616);
  assign tmp39724 = ~(l1 ? tmp39434 : tmp39725);
  assign tmp39722 = s1 ? tmp39723 : tmp39724;
  assign tmp39728 = l1 ? tmp39630 : tmp39588;
  assign tmp39727 = ~(s0 ? tmp39596 : tmp39728);
  assign tmp39726 = ~(s1 ? tmp39625 : tmp39727);
  assign tmp39721 = ~(s2 ? tmp39722 : tmp39726);
  assign tmp39711 = s3 ? tmp39712 : tmp39721;
  assign tmp39731 = ~(l1 ? tmp39587 : tmp39375);
  assign tmp39730 = s2 ? tmp39633 : tmp39731;
  assign tmp39735 = ~(l1 ? tmp39681 : tmp39541);
  assign tmp39734 = s0 ? tmp39723 : tmp39735;
  assign tmp39733 = s1 ? tmp39734 : tmp39648;
  assign tmp39732 = ~(s2 ? tmp39733 : tmp39650);
  assign tmp39729 = s3 ? tmp39730 : tmp39732;
  assign tmp39710 = s4 ? tmp39711 : tmp39729;
  assign tmp39741 = l1 ? tmp39434 : tmp39725;
  assign tmp39740 = s0 ? tmp39741 : 0;
  assign tmp39739 = s1 ? tmp39740 : tmp39658;
  assign tmp39744 = ~(l2 ? tmp39440 : tmp39389);
  assign tmp39743 = l1 ? 1 : tmp39744;
  assign tmp39742 = s1 ? tmp39743 : tmp39661;
  assign tmp39738 = s2 ? tmp39739 : tmp39742;
  assign tmp39737 = s3 ? tmp39738 : tmp39662;
  assign tmp39747 = ~(l1 ? tmp39630 : tmp39375);
  assign tmp39746 = s2 ? tmp39670 : tmp39747;
  assign tmp39745 = s3 ? tmp39746 : tmp39672;
  assign tmp39736 = s4 ? tmp39737 : tmp39745;
  assign tmp39709 = s5 ? tmp39710 : tmp39736;
  assign tmp39676 = s6 ? tmp39677 : tmp39709;
  assign tmp39675 = s7 ? tmp39370 : tmp39676;
  assign tmp39368 = s8 ? tmp39369 : tmp39675;
  assign tmp39755 = ~(l2 ? tmp39440 : tmp39460);
  assign tmp39754 = l1 ? tmp39378 : tmp39755;
  assign tmp39758 = l2 ? tmp39403 : tmp39381;
  assign tmp39757 = l1 ? tmp39758 : tmp39375;
  assign tmp39759 = ~(l1 ? tmp39527 : tmp39755);
  assign tmp39756 = ~(s0 ? tmp39757 : tmp39759);
  assign tmp39753 = s1 ? tmp39754 : tmp39756;
  assign tmp39763 = l1 ? tmp39575 : tmp39403;
  assign tmp39765 = ~(l2 ? tmp39376 : tmp39460);
  assign tmp39764 = ~(l1 ? tmp39434 : tmp39765);
  assign tmp39762 = s0 ? tmp39763 : tmp39764;
  assign tmp39767 = l1 ? tmp39575 : tmp39621;
  assign tmp39766 = s0 ? tmp39767 : tmp39764;
  assign tmp39761 = s1 ? tmp39762 : tmp39766;
  assign tmp39770 = ~(l1 ? 1 : tmp39386);
  assign tmp39769 = s0 ? tmp39767 : tmp39770;
  assign tmp39772 = l1 ? tmp39434 : tmp39765;
  assign tmp39773 = ~(l1 ? tmp39575 : tmp39493);
  assign tmp39771 = ~(s0 ? tmp39772 : tmp39773);
  assign tmp39768 = s1 ? tmp39769 : tmp39771;
  assign tmp39760 = ~(s2 ? tmp39761 : tmp39768);
  assign tmp39752 = s3 ? tmp39753 : tmp39760;
  assign tmp39778 = l1 ? 1 : tmp39755;
  assign tmp39779 = ~(l1 ? tmp39758 : 1);
  assign tmp39777 = s0 ? tmp39778 : tmp39779;
  assign tmp39781 = l1 ? tmp39575 : tmp39493;
  assign tmp39780 = ~(s0 ? tmp39781 : tmp39764);
  assign tmp39776 = s1 ? tmp39777 : tmp39780;
  assign tmp39785 = l2 ? tmp39403 : tmp39386;
  assign tmp39784 = ~(l1 ? tmp39785 : 1);
  assign tmp39783 = s0 ? tmp39754 : tmp39784;
  assign tmp39786 = l1 ? 1 : tmp39478;
  assign tmp39782 = s1 ? tmp39783 : tmp39786;
  assign tmp39775 = s2 ? tmp39776 : tmp39782;
  assign tmp39788 = s1 ? tmp39757 : tmp39531;
  assign tmp39790 = s0 ? tmp39603 : tmp39772;
  assign tmp39789 = ~(s1 ? tmp39772 : tmp39790);
  assign tmp39787 = ~(s2 ? tmp39788 : tmp39789);
  assign tmp39774 = s3 ? tmp39775 : tmp39787;
  assign tmp39751 = s4 ? tmp39752 : tmp39774;
  assign tmp39797 = l1 ? tmp39527 : tmp39755;
  assign tmp39796 = s0 ? tmp39797 : tmp39487;
  assign tmp39798 = ~(l1 ? tmp39575 : tmp39403);
  assign tmp39795 = s1 ? tmp39796 : tmp39798;
  assign tmp39801 = ~(l2 ? tmp39440 : tmp39398);
  assign tmp39800 = l1 ? tmp39527 : tmp39801;
  assign tmp39803 = ~(l2 ? tmp39403 : 1);
  assign tmp39802 = s0 ? tmp39772 : tmp39803;
  assign tmp39799 = s1 ? tmp39800 : tmp39802;
  assign tmp39794 = s2 ? tmp39795 : tmp39799;
  assign tmp39807 = ~(l2 ? tmp39376 : tmp39398);
  assign tmp39806 = ~(l1 ? tmp39434 : tmp39807);
  assign tmp39805 = s1 ? tmp39621 : tmp39806;
  assign tmp39810 = l1 ? tmp39575 : tmp39588;
  assign tmp39811 = l1 ? tmp39621 : tmp39588;
  assign tmp39809 = ~(s0 ? tmp39810 : tmp39811);
  assign tmp39808 = ~(s1 ? tmp39625 : tmp39809);
  assign tmp39804 = ~(s2 ? tmp39805 : tmp39808);
  assign tmp39793 = s3 ? tmp39794 : tmp39804;
  assign tmp39816 = l1 ? tmp39434 : tmp39801;
  assign tmp39815 = s0 ? tmp39635 : tmp39816;
  assign tmp39818 = ~(l1 ? tmp39403 : tmp39375);
  assign tmp39817 = s0 ? tmp39786 : tmp39818;
  assign tmp39814 = s1 ? tmp39815 : tmp39817;
  assign tmp39819 = ~(l1 ? tmp39575 : tmp39621);
  assign tmp39813 = s2 ? tmp39814 : tmp39819;
  assign tmp39823 = l1 ? tmp39630 : tmp39621;
  assign tmp39824 = ~(l1 ? tmp39378 : tmp39435);
  assign tmp39822 = s0 ? tmp39823 : tmp39824;
  assign tmp39821 = s1 ? tmp39822 : tmp39648;
  assign tmp39820 = ~(s2 ? tmp39821 : tmp39650);
  assign tmp39812 = s3 ? tmp39813 : tmp39820;
  assign tmp39792 = s4 ? tmp39793 : tmp39812;
  assign tmp39830 = l1 ? tmp39434 : tmp39807;
  assign tmp39829 = s0 ? tmp39830 : 0;
  assign tmp39828 = s1 ? tmp39829 : tmp39658;
  assign tmp39831 = s1 ? tmp39786 : tmp39661;
  assign tmp39827 = s2 ? tmp39828 : tmp39831;
  assign tmp39834 = ~(l2 ? tmp39430 : tmp39403);
  assign tmp39833 = ~(s1 ? tmp39666 : tmp39834);
  assign tmp39832 = ~(s2 ? tmp39663 : tmp39833);
  assign tmp39826 = s3 ? tmp39827 : tmp39832;
  assign tmp39837 = ~(l1 ? tmp39630 : tmp39621);
  assign tmp39836 = s2 ? tmp39670 : tmp39837;
  assign tmp39840 = l2 ? tmp39430 : tmp39460;
  assign tmp39839 = ~(l1 ? tmp39630 : tmp39840);
  assign tmp39838 = s1 ? tmp39673 : tmp39839;
  assign tmp39835 = s3 ? tmp39836 : tmp39838;
  assign tmp39825 = s4 ? tmp39826 : tmp39835;
  assign tmp39791 = s5 ? tmp39792 : tmp39825;
  assign tmp39750 = s6 ? tmp39751 : tmp39791;
  assign tmp39749 = s7 ? tmp39370 : tmp39750;
  assign tmp39748 = s8 ? tmp39675 : tmp39749;
  assign tmp39367 = s9 ? tmp39368 : tmp39748;
  assign tmp39848 = ~(s0 ? tmp39757 : tmp39570);
  assign tmp39847 = s1 ? tmp39566 : tmp39848;
  assign tmp39852 = l1 ? tmp39575 : tmp39402;
  assign tmp39853 = ~(l1 ? tmp39434 : tmp39690);
  assign tmp39851 = s0 ? tmp39852 : tmp39853;
  assign tmp39854 = s0 ? tmp39580 : tmp39853;
  assign tmp39850 = s1 ? tmp39851 : tmp39854;
  assign tmp39856 = s0 ? tmp39580 : tmp39770;
  assign tmp39858 = l1 ? tmp39434 : tmp39690;
  assign tmp39859 = ~(l1 ? tmp39575 : tmp39588);
  assign tmp39857 = ~(s0 ? tmp39858 : tmp39859);
  assign tmp39855 = s1 ? tmp39856 : tmp39857;
  assign tmp39849 = ~(s2 ? tmp39850 : tmp39855);
  assign tmp39846 = s3 ? tmp39847 : tmp39849;
  assign tmp39863 = s0 ? tmp39593 : tmp39779;
  assign tmp39864 = ~(s0 ? tmp39810 : tmp39853);
  assign tmp39862 = s1 ? tmp39863 : tmp39864;
  assign tmp39866 = s0 ? tmp39566 : tmp39784;
  assign tmp39865 = s1 ? tmp39866 : tmp39786;
  assign tmp39861 = s2 ? tmp39862 : tmp39865;
  assign tmp39869 = s0 ? tmp39603 : tmp39858;
  assign tmp39868 = ~(s1 ? tmp39858 : tmp39869);
  assign tmp39867 = ~(s2 ? tmp39788 : tmp39868);
  assign tmp39860 = s3 ? tmp39861 : tmp39867;
  assign tmp39845 = s4 ? tmp39846 : tmp39860;
  assign tmp39875 = ~(l1 ? tmp39575 : tmp39402);
  assign tmp39874 = s1 ? tmp39610 : tmp39875;
  assign tmp39877 = l1 ? tmp39527 : tmp39637;
  assign tmp39878 = s0 ? tmp39858 : tmp39803;
  assign tmp39876 = s1 ? tmp39877 : tmp39878;
  assign tmp39873 = s2 ? tmp39874 : tmp39876;
  assign tmp39880 = s1 ? tmp39620 : tmp39724;
  assign tmp39879 = ~(s2 ? tmp39880 : tmp39808);
  assign tmp39872 = s3 ? tmp39873 : tmp39879;
  assign tmp39885 = l1 ? tmp39434 : tmp39637;
  assign tmp39884 = s0 ? tmp39635 : tmp39885;
  assign tmp39883 = s1 ? tmp39884 : tmp39817;
  assign tmp39886 = ~(l1 ? tmp39575 : tmp39375);
  assign tmp39882 = s2 ? tmp39883 : tmp39886;
  assign tmp39889 = s0 ? tmp39723 : tmp39647;
  assign tmp39888 = s1 ? tmp39889 : tmp39648;
  assign tmp39887 = ~(s2 ? tmp39888 : tmp39650);
  assign tmp39881 = s3 ? tmp39882 : tmp39887;
  assign tmp39871 = s4 ? tmp39872 : tmp39881;
  assign tmp39870 = s5 ? tmp39871 : tmp39736;
  assign tmp39844 = s6 ? tmp39845 : tmp39870;
  assign tmp39843 = s7 ? tmp39370 : tmp39844;
  assign tmp39842 = s8 ? tmp39843 : tmp39370;
  assign tmp39898 = ~(l1 ? tmp39575 : tmp39429);
  assign tmp39897 = s1 ? tmp39483 : tmp39898;
  assign tmp39896 = s2 ? tmp39633 : tmp39897;
  assign tmp39895 = s3 ? tmp39896 : tmp39643;
  assign tmp39894 = s4 ? tmp39607 : tmp39895;
  assign tmp39893 = s5 ? tmp39894 : tmp39652;
  assign tmp39892 = s6 ? tmp39563 : tmp39893;
  assign tmp39891 = s7 ? tmp39892 : tmp39750;
  assign tmp39899 = s7 ? tmp39676 : tmp39844;
  assign tmp39890 = s8 ? tmp39891 : tmp39899;
  assign tmp39841 = s9 ? tmp39842 : tmp39890;
  assign tmp39366 = s10 ? tmp39367 : tmp39841;
  assign tmp39903 = s7 ? tmp39562 : tmp39750;
  assign tmp39902 = s8 ? tmp39903 : tmp39899;
  assign tmp39901 = s9 ? tmp39842 : tmp39902;
  assign tmp39900 = s10 ? tmp39367 : tmp39901;
  assign tmp39365 = s11 ? tmp39366 : tmp39900;
  assign tmp39915 = l2 ? tmp39378 : tmp39460;
  assign tmp39914 = l1 ? tmp39915 : tmp39801;
  assign tmp39918 = l2 ? tmp39376 : tmp39386;
  assign tmp39917 = l1 ? tmp39785 : tmp39918;
  assign tmp39919 = ~(l1 ? tmp39547 : tmp39801);
  assign tmp39916 = ~(s0 ? tmp39917 : tmp39919);
  assign tmp39913 = s1 ? tmp39914 : tmp39916;
  assign tmp39923 = l1 ? tmp39918 : tmp39384;
  assign tmp39925 = l2 ? tmp39460 : tmp39440;
  assign tmp39926 = ~(l2 ? tmp39430 : tmp39398);
  assign tmp39924 = ~(l1 ? tmp39925 : tmp39926);
  assign tmp39922 = s0 ? tmp39923 : tmp39924;
  assign tmp39928 = l1 ? tmp39918 : tmp39575;
  assign tmp39927 = s0 ? tmp39928 : tmp39924;
  assign tmp39921 = s1 ? tmp39922 : tmp39927;
  assign tmp39930 = s0 ? tmp39928 : tmp39401;
  assign tmp39932 = l1 ? tmp39925 : tmp39926;
  assign tmp39934 = l2 ? tmp39376 : tmp39398;
  assign tmp39933 = ~(l1 ? tmp39918 : tmp39934);
  assign tmp39931 = ~(s0 ? tmp39932 : tmp39933);
  assign tmp39929 = s1 ? tmp39930 : tmp39931;
  assign tmp39920 = ~(s2 ? tmp39921 : tmp39929);
  assign tmp39912 = s3 ? tmp39913 : tmp39920;
  assign tmp39939 = l1 ? tmp39480 : tmp39801;
  assign tmp39940 = ~(l1 ? tmp39785 : tmp39385);
  assign tmp39938 = s0 ? tmp39939 : tmp39940;
  assign tmp39942 = l1 ? tmp39918 : tmp39934;
  assign tmp39941 = ~(s0 ? tmp39942 : tmp39924);
  assign tmp39937 = s1 ? tmp39938 : tmp39941;
  assign tmp39944 = s0 ? tmp39914 : tmp39420;
  assign tmp39946 = l1 ? tmp39480 : tmp39478;
  assign tmp39945 = s0 ? tmp39946 : tmp39424;
  assign tmp39943 = s1 ? tmp39944 : tmp39945;
  assign tmp39936 = s2 ? tmp39937 : tmp39943;
  assign tmp39949 = s0 ? tmp39432 : tmp39531;
  assign tmp39948 = s1 ? tmp39917 : tmp39949;
  assign tmp39951 = s0 ? tmp39603 : tmp39932;
  assign tmp39950 = ~(s1 ? tmp39932 : tmp39951);
  assign tmp39947 = ~(s2 ? tmp39948 : tmp39950);
  assign tmp39935 = s3 ? tmp39936 : tmp39947;
  assign tmp39911 = s4 ? tmp39912 : tmp39935;
  assign tmp39958 = l1 ? tmp39547 : tmp39801;
  assign tmp39957 = s0 ? tmp39958 : tmp39420;
  assign tmp39959 = ~(s0 ? tmp39448 : tmp39923);
  assign tmp39956 = s1 ? tmp39957 : tmp39959;
  assign tmp39961 = s0 ? tmp39448 : tmp39919;
  assign tmp39962 = ~(s0 ? tmp39932 : tmp39452);
  assign tmp39960 = ~(s1 ? tmp39961 : tmp39962);
  assign tmp39955 = s2 ? tmp39956 : tmp39960;
  assign tmp39966 = l1 ? tmp39375 : tmp39575;
  assign tmp39965 = s0 ? tmp39456 : tmp39966;
  assign tmp39968 = ~(l1 ? tmp39469 : tmp39926);
  assign tmp39967 = s0 ? tmp39456 : tmp39968;
  assign tmp39964 = s1 ? tmp39965 : tmp39967;
  assign tmp39972 = l2 ? tmp39430 : tmp39386;
  assign tmp39971 = l1 ? tmp39972 : tmp39840;
  assign tmp39973 = l1 ? tmp39429 : tmp39840;
  assign tmp39970 = ~(s0 ? tmp39971 : tmp39973);
  assign tmp39969 = ~(s1 ? tmp39625 : tmp39970);
  assign tmp39963 = ~(s2 ? tmp39964 : tmp39969);
  assign tmp39954 = s3 ? tmp39955 : tmp39963;
  assign tmp39978 = l1 ? tmp39469 : tmp39801;
  assign tmp39977 = s0 ? tmp39635 : tmp39978;
  assign tmp39980 = ~(l1 ? tmp39402 : tmp39375);
  assign tmp39979 = s0 ? tmp39946 : tmp39980;
  assign tmp39976 = s1 ? tmp39977 : tmp39979;
  assign tmp39981 = ~(l1 ? tmp39918 : tmp39621);
  assign tmp39975 = s2 ? tmp39976 : tmp39981;
  assign tmp39985 = l1 ? tmp39429 : tmp39621;
  assign tmp39986 = ~(l1 ? tmp39915 : tmp39435);
  assign tmp39984 = s0 ? tmp39985 : tmp39986;
  assign tmp39987 = ~(l1 ? tmp39469 : tmp39604);
  assign tmp39983 = s1 ? tmp39984 : tmp39987;
  assign tmp39982 = ~(s2 ? tmp39983 : tmp39650);
  assign tmp39974 = s3 ? tmp39975 : tmp39982;
  assign tmp39953 = s4 ? tmp39954 : tmp39974;
  assign tmp39993 = l1 ? tmp39469 : tmp39926;
  assign tmp39992 = s0 ? tmp39993 : 0;
  assign tmp39991 = s1 ? tmp39992 : tmp39658;
  assign tmp39995 = l1 ? tmp39480 : tmp39404;
  assign tmp39996 = ~(l1 ? tmp39429 : tmp39480);
  assign tmp39994 = s1 ? tmp39995 : tmp39996;
  assign tmp39990 = s2 ? tmp39991 : tmp39994;
  assign tmp39999 = ~(l1 ? tmp39429 : tmp39630);
  assign tmp39998 = ~(s1 ? tmp39666 : tmp39999);
  assign tmp39997 = ~(s2 ? tmp39663 : tmp39998);
  assign tmp39989 = s3 ? tmp39990 : tmp39997;
  assign tmp40002 = ~(l1 ? tmp39429 : tmp39621);
  assign tmp40001 = s2 ? tmp39670 : tmp40002;
  assign tmp40004 = ~(l1 ? tmp39429 : tmp39840);
  assign tmp40003 = s1 ? tmp39673 : tmp40004;
  assign tmp40000 = s3 ? tmp40001 : tmp40003;
  assign tmp39988 = s4 ? tmp39989 : tmp40000;
  assign tmp39952 = s5 ? tmp39953 : tmp39988;
  assign tmp39910 = s6 ? tmp39911 : tmp39952;
  assign tmp39909 = s7 ? tmp39370 : tmp39910;
  assign tmp40010 = l1 ? tmp39460 : tmp39801;
  assign tmp40012 = l1 ? tmp39385 : tmp39918;
  assign tmp40014 = l2 ? tmp39403 : tmp39440;
  assign tmp40013 = ~(l1 ? tmp40014 : tmp39801);
  assign tmp40011 = ~(s0 ? tmp40012 : tmp40013);
  assign tmp40009 = s1 ? tmp40010 : tmp40011;
  assign tmp40018 = l1 ? tmp39972 : tmp39758;
  assign tmp40019 = ~(l1 ? tmp39925 : tmp39807);
  assign tmp40017 = s0 ? tmp40018 : tmp40019;
  assign tmp40021 = l1 ? tmp39972 : tmp39575;
  assign tmp40020 = s0 ? tmp40021 : tmp40019;
  assign tmp40016 = s1 ? tmp40017 : tmp40020;
  assign tmp40024 = ~(l1 ? tmp39402 : tmp39478);
  assign tmp40023 = s0 ? tmp40021 : tmp40024;
  assign tmp40026 = l1 ? tmp39925 : tmp39807;
  assign tmp40027 = ~(l1 ? tmp39972 : tmp39934);
  assign tmp40025 = ~(s0 ? tmp40026 : tmp40027);
  assign tmp40022 = s1 ? tmp40023 : tmp40025;
  assign tmp40015 = ~(s2 ? tmp40016 : tmp40022);
  assign tmp40008 = s3 ? tmp40009 : tmp40015;
  assign tmp40032 = l1 ? tmp39403 : tmp39801;
  assign tmp40031 = s0 ? tmp40032 : tmp39420;
  assign tmp40034 = l1 ? tmp39972 : tmp39934;
  assign tmp40033 = ~(s0 ? tmp40034 : tmp40019);
  assign tmp40030 = s1 ? tmp40031 : tmp40033;
  assign tmp40036 = s0 ? tmp40010 : tmp39420;
  assign tmp40037 = l1 ? tmp39403 : tmp39478;
  assign tmp40035 = s1 ? tmp40036 : tmp40037;
  assign tmp40029 = s2 ? tmp40030 : tmp40035;
  assign tmp40039 = s1 ? tmp40012 : tmp39531;
  assign tmp40041 = s0 ? tmp39603 : tmp40026;
  assign tmp40040 = ~(s1 ? tmp40026 : tmp40041);
  assign tmp40038 = ~(s2 ? tmp40039 : tmp40040);
  assign tmp40028 = s3 ? tmp40029 : tmp40038;
  assign tmp40007 = s4 ? tmp40008 : tmp40028;
  assign tmp40048 = l1 ? tmp40014 : tmp39801;
  assign tmp40047 = s0 ? tmp40048 : tmp39420;
  assign tmp40049 = ~(s0 ? tmp39448 : tmp40018);
  assign tmp40046 = s1 ? tmp40047 : tmp40049;
  assign tmp40051 = s0 ? tmp39448 : tmp40013;
  assign tmp40053 = ~(l1 ? 1 : tmp39785);
  assign tmp40052 = ~(s0 ? tmp40026 : tmp40053);
  assign tmp40050 = ~(s1 ? tmp40051 : tmp40052);
  assign tmp40045 = s2 ? tmp40046 : tmp40050;
  assign tmp40056 = l1 ? tmp39429 : tmp39575;
  assign tmp40057 = ~(l1 ? tmp39469 : tmp39807);
  assign tmp40055 = s1 ? tmp40056 : tmp40057;
  assign tmp40060 = l1 ? tmp39972 : tmp39493;
  assign tmp40061 = l1 ? tmp39429 : tmp39493;
  assign tmp40059 = ~(s0 ? tmp40060 : tmp40061);
  assign tmp40058 = ~(s1 ? tmp39625 : tmp40059);
  assign tmp40054 = ~(s2 ? tmp40055 : tmp40058);
  assign tmp40044 = s3 ? tmp40045 : tmp40054;
  assign tmp40066 = l1 ? tmp39925 : tmp39801;
  assign tmp40065 = s0 ? tmp39635 : tmp40066;
  assign tmp40068 = ~(l1 ? 1 : tmp39375);
  assign tmp40067 = s0 ? tmp40037 : tmp40068;
  assign tmp40064 = s1 ? tmp40065 : tmp40067;
  assign tmp40069 = ~(l1 ? tmp39972 : tmp39621);
  assign tmp40063 = s2 ? tmp40064 : tmp40069;
  assign tmp40073 = ~(l1 ? tmp39460 : tmp39435);
  assign tmp40072 = s0 ? tmp39985 : tmp40073;
  assign tmp40071 = s1 ? tmp40072 : tmp39987;
  assign tmp40070 = ~(s2 ? tmp40071 : tmp39650);
  assign tmp40062 = s3 ? tmp40063 : tmp40070;
  assign tmp40043 = s4 ? tmp40044 : tmp40062;
  assign tmp40079 = l1 ? tmp39469 : tmp39807;
  assign tmp40078 = s0 ? tmp40079 : 0;
  assign tmp40077 = s1 ? tmp40078 : tmp39658;
  assign tmp40080 = s1 ? tmp39946 : tmp39996;
  assign tmp40076 = s2 ? tmp40077 : tmp40080;
  assign tmp40075 = s3 ? tmp40076 : tmp39997;
  assign tmp40074 = s4 ? tmp40075 : tmp40000;
  assign tmp40042 = s5 ? tmp40043 : tmp40074;
  assign tmp40006 = s6 ? tmp40007 : tmp40042;
  assign tmp40005 = s7 ? tmp39370 : tmp40006;
  assign tmp39908 = s8 ? tmp39909 : tmp40005;
  assign tmp40087 = l1 ? tmp39915 : tmp39637;
  assign tmp40086 = s1 ? tmp40087 : tmp39916;
  assign tmp40091 = l1 ? tmp39918 : tmp39785;
  assign tmp40092 = ~(l1 ? tmp39469 : tmp39725);
  assign tmp40090 = s0 ? tmp40091 : tmp40092;
  assign tmp40093 = s0 ? tmp39918 : tmp40092;
  assign tmp40089 = s1 ? tmp40090 : tmp40093;
  assign tmp40096 = ~(l1 ? 1 : tmp39478);
  assign tmp40095 = s0 ? tmp39918 : tmp40096;
  assign tmp40098 = l1 ? tmp39469 : tmp39725;
  assign tmp40100 = l2 ? tmp39376 : tmp39616;
  assign tmp40099 = ~(l1 ? tmp39918 : tmp40100);
  assign tmp40097 = ~(s0 ? tmp40098 : tmp40099);
  assign tmp40094 = s1 ? tmp40095 : tmp40097;
  assign tmp40088 = ~(s2 ? tmp40089 : tmp40094);
  assign tmp40085 = s3 ? tmp40086 : tmp40088;
  assign tmp40105 = l1 ? tmp39918 : tmp40100;
  assign tmp40104 = ~(s0 ? tmp40105 : tmp40092);
  assign tmp40103 = s1 ? tmp39938 : tmp40104;
  assign tmp40107 = s0 ? tmp40087 : tmp39940;
  assign tmp40106 = s1 ? tmp40107 : tmp39946;
  assign tmp40102 = s2 ? tmp40103 : tmp40106;
  assign tmp40109 = s1 ? tmp39917 : tmp39531;
  assign tmp40111 = s0 ? tmp39603 : tmp40098;
  assign tmp40110 = ~(s1 ? tmp40098 : tmp40111);
  assign tmp40108 = ~(s2 ? tmp40109 : tmp40110);
  assign tmp40101 = s3 ? tmp40102 : tmp40108;
  assign tmp40084 = s4 ? tmp40085 : tmp40101;
  assign tmp40117 = ~(s0 ? tmp39448 : tmp40091);
  assign tmp40116 = s1 ? tmp39957 : tmp40117;
  assign tmp40120 = ~(l1 ? tmp39402 : tmp39785);
  assign tmp40119 = ~(s0 ? tmp40098 : tmp40120);
  assign tmp40118 = ~(s1 ? tmp39961 : tmp40119);
  assign tmp40115 = s2 ? tmp40116 : tmp40118;
  assign tmp40123 = l1 ? tmp39375 : tmp39918;
  assign tmp40122 = s1 ? tmp40123 : tmp40057;
  assign tmp40126 = l1 ? tmp39918 : tmp39493;
  assign tmp40127 = l1 ? tmp39375 : tmp39493;
  assign tmp40125 = ~(s0 ? tmp40126 : tmp40127);
  assign tmp40124 = ~(s1 ? tmp39625 : tmp40125);
  assign tmp40121 = ~(s2 ? tmp40122 : tmp40124);
  assign tmp40114 = s3 ? tmp40115 : tmp40121;
  assign tmp40113 = s4 ? tmp40114 : tmp39974;
  assign tmp40112 = s5 ? tmp40113 : tmp40074;
  assign tmp40083 = s6 ? tmp40084 : tmp40112;
  assign tmp40082 = s7 ? tmp39370 : tmp40083;
  assign tmp40081 = s8 ? tmp40005 : tmp40082;
  assign tmp39907 = s9 ? tmp39908 : tmp40081;
  assign tmp40137 = l1 ? tmp39918 : tmp39758;
  assign tmp40136 = s0 ? tmp40137 : tmp40057;
  assign tmp40138 = s0 ? tmp39928 : tmp40057;
  assign tmp40135 = s1 ? tmp40136 : tmp40138;
  assign tmp40140 = s0 ? tmp39928 : tmp40096;
  assign tmp40141 = ~(s0 ? tmp40079 : tmp39933);
  assign tmp40139 = s1 ? tmp40140 : tmp40141;
  assign tmp40134 = ~(s2 ? tmp40135 : tmp40139);
  assign tmp40133 = s3 ? tmp39913 : tmp40134;
  assign tmp40145 = ~(s0 ? tmp39942 : tmp40057);
  assign tmp40144 = s1 ? tmp39938 : tmp40145;
  assign tmp40147 = s0 ? tmp39914 : tmp39940;
  assign tmp40146 = s1 ? tmp40147 : tmp39946;
  assign tmp40143 = s2 ? tmp40144 : tmp40146;
  assign tmp40150 = s0 ? tmp39603 : tmp40079;
  assign tmp40149 = ~(s1 ? tmp40079 : tmp40150);
  assign tmp40148 = ~(s2 ? tmp40109 : tmp40149);
  assign tmp40142 = s3 ? tmp40143 : tmp40148;
  assign tmp40132 = s4 ? tmp40133 : tmp40142;
  assign tmp40156 = ~(s0 ? tmp39448 : tmp40137);
  assign tmp40155 = s1 ? tmp39957 : tmp40156;
  assign tmp40158 = ~(s0 ? tmp40079 : tmp40120);
  assign tmp40157 = ~(s1 ? tmp39961 : tmp40158);
  assign tmp40154 = s2 ? tmp40155 : tmp40157;
  assign tmp40160 = s1 ? tmp39966 : tmp40057;
  assign tmp40159 = ~(s2 ? tmp40160 : tmp40124);
  assign tmp40153 = s3 ? tmp40154 : tmp40159;
  assign tmp40152 = s4 ? tmp40153 : tmp39974;
  assign tmp40151 = s5 ? tmp40152 : tmp40074;
  assign tmp40131 = s6 ? tmp40132 : tmp40151;
  assign tmp40130 = s7 ? tmp39370 : tmp40131;
  assign tmp40129 = s8 ? tmp40130 : tmp39370;
  assign tmp40166 = ~(s2 ? tmp40109 : tmp39950);
  assign tmp40165 = s3 ? tmp39936 : tmp40166;
  assign tmp40164 = s4 ? tmp39912 : tmp40165;
  assign tmp40172 = s0 ? tmp39932 : tmp39452;
  assign tmp40171 = s1 ? tmp39958 : tmp40172;
  assign tmp40170 = s2 ? tmp39956 : tmp40171;
  assign tmp40174 = s1 ? tmp39965 : tmp39968;
  assign tmp40173 = ~(s2 ? tmp40174 : tmp39969);
  assign tmp40169 = s3 ? tmp40170 : tmp40173;
  assign tmp40168 = s4 ? tmp40169 : tmp39974;
  assign tmp40167 = s5 ? tmp40168 : tmp39988;
  assign tmp40163 = s6 ? tmp40164 : tmp40167;
  assign tmp40181 = s0 ? tmp40098 : tmp40120;
  assign tmp40180 = s1 ? tmp39958 : tmp40181;
  assign tmp40179 = s2 ? tmp40116 : tmp40180;
  assign tmp40178 = s3 ? tmp40179 : tmp40121;
  assign tmp40177 = s4 ? tmp40178 : tmp39974;
  assign tmp40176 = s5 ? tmp40177 : tmp40074;
  assign tmp40175 = s6 ? tmp40084 : tmp40176;
  assign tmp40162 = s7 ? tmp40163 : tmp40175;
  assign tmp40189 = s0 ? tmp40026 : tmp40053;
  assign tmp40188 = s1 ? tmp40048 : tmp40189;
  assign tmp40187 = s2 ? tmp40046 : tmp40188;
  assign tmp40186 = s3 ? tmp40187 : tmp40054;
  assign tmp40185 = s4 ? tmp40186 : tmp40062;
  assign tmp40184 = s5 ? tmp40185 : tmp40074;
  assign tmp40183 = s6 ? tmp40007 : tmp40184;
  assign tmp40196 = s0 ? tmp40079 : tmp40120;
  assign tmp40195 = s1 ? tmp39958 : tmp40196;
  assign tmp40194 = s2 ? tmp40155 : tmp40195;
  assign tmp40193 = s3 ? tmp40194 : tmp40159;
  assign tmp40192 = s4 ? tmp40193 : tmp39974;
  assign tmp40191 = s5 ? tmp40192 : tmp40074;
  assign tmp40190 = s6 ? tmp40132 : tmp40191;
  assign tmp40182 = s7 ? tmp40183 : tmp40190;
  assign tmp40161 = s8 ? tmp40162 : tmp40182;
  assign tmp40128 = s9 ? tmp40129 : tmp40161;
  assign tmp39906 = s10 ? tmp39907 : tmp40128;
  assign tmp40200 = s7 ? tmp39910 : tmp40083;
  assign tmp40201 = s7 ? tmp40006 : tmp40131;
  assign tmp40199 = s8 ? tmp40200 : tmp40201;
  assign tmp40198 = s9 ? tmp40129 : tmp40199;
  assign tmp40197 = s10 ? tmp39907 : tmp40198;
  assign tmp39905 = s11 ? tmp39906 : tmp40197;
  assign tmp40211 = l1 ? tmp39915 : tmp39435;
  assign tmp40214 = ~(l2 ? tmp39378 : tmp39440);
  assign tmp40213 = l1 ? tmp39785 : tmp40214;
  assign tmp40215 = ~(l1 ? tmp39547 : tmp39435);
  assign tmp40212 = ~(s0 ? tmp40213 : tmp40215);
  assign tmp40210 = s1 ? tmp40211 : tmp40212;
  assign tmp40219 = l1 ? tmp39918 : tmp39381;
  assign tmp40218 = s0 ? tmp40219 : tmp39987;
  assign tmp40222 = ~(l2 ? tmp39378 : tmp39379);
  assign tmp40221 = l1 ? tmp39918 : tmp40222;
  assign tmp40220 = s0 ? tmp40221 : tmp39987;
  assign tmp40217 = s1 ? tmp40218 : tmp40220;
  assign tmp40225 = ~(l1 ? tmp39402 : 1);
  assign tmp40224 = s0 ? tmp40221 : tmp40225;
  assign tmp40227 = l1 ? tmp39469 : tmp39604;
  assign tmp40229 = ~(l2 ? tmp39378 : tmp39430);
  assign tmp40228 = ~(l1 ? tmp39918 : tmp40229);
  assign tmp40226 = ~(s0 ? tmp40227 : tmp40228);
  assign tmp40223 = s1 ? tmp40224 : tmp40226;
  assign tmp40216 = ~(s2 ? tmp40217 : tmp40223);
  assign tmp40209 = s3 ? tmp40210 : tmp40216;
  assign tmp40234 = ~(l1 ? tmp39785 : tmp39386);
  assign tmp40233 = s0 ? tmp39491 : tmp40234;
  assign tmp40236 = l1 ? tmp39918 : tmp40229;
  assign tmp40235 = ~(s0 ? tmp40236 : tmp39987);
  assign tmp40232 = s1 ? tmp40233 : tmp40235;
  assign tmp40238 = s0 ? tmp40211 : tmp39420;
  assign tmp40239 = s0 ? tmp39520 : tmp39424;
  assign tmp40237 = s1 ? tmp40238 : tmp40239;
  assign tmp40231 = s2 ? tmp40232 : tmp40237;
  assign tmp40241 = s1 ? tmp40213 : tmp39949;
  assign tmp40243 = s0 ? tmp39603 : tmp40227;
  assign tmp40242 = ~(s1 ? tmp40227 : tmp40243);
  assign tmp40240 = ~(s2 ? tmp40241 : tmp40242);
  assign tmp40230 = s3 ? tmp40231 : tmp40240;
  assign tmp40208 = s4 ? tmp40209 : tmp40230;
  assign tmp40250 = ~(l1 ? tmp39385 : tmp39386);
  assign tmp40249 = s0 ? tmp39546 : tmp40250;
  assign tmp40251 = ~(l1 ? tmp39918 : tmp39381);
  assign tmp40248 = s1 ? tmp40249 : tmp40251;
  assign tmp40253 = s0 ? tmp40227 : tmp39583;
  assign tmp40252 = s1 ? tmp39546 : tmp40253;
  assign tmp40247 = s2 ? tmp40248 : tmp40252;
  assign tmp40256 = l1 ? tmp39375 : tmp40222;
  assign tmp40255 = s1 ? tmp40256 : tmp39987;
  assign tmp40259 = l1 ? tmp39918 : tmp39377;
  assign tmp40258 = ~(s0 ? tmp40259 : tmp40127);
  assign tmp40257 = ~(s1 ? tmp39625 : tmp40258);
  assign tmp40254 = ~(s2 ? tmp40255 : tmp40257);
  assign tmp40246 = s3 ? tmp40247 : tmp40254;
  assign tmp40263 = s0 ? tmp39635 : tmp39468;
  assign tmp40264 = s0 ? tmp39520 : tmp39980;
  assign tmp40262 = s1 ? tmp40263 : tmp40264;
  assign tmp40265 = ~(l1 ? tmp39918 : tmp39388);
  assign tmp40261 = s2 ? tmp40262 : tmp40265;
  assign tmp40269 = l1 ? tmp39429 : tmp39388;
  assign tmp40268 = s0 ? tmp40269 : tmp39986;
  assign tmp40267 = s1 ? tmp40268 : tmp39987;
  assign tmp40266 = ~(s2 ? tmp40267 : tmp39650);
  assign tmp40260 = s3 ? tmp40261 : tmp40266;
  assign tmp40245 = s4 ? tmp40246 : tmp40260;
  assign tmp40274 = s0 ? tmp40227 : 0;
  assign tmp40273 = s1 ? tmp40274 : tmp39658;
  assign tmp40275 = s1 ? tmp39520 : tmp39996;
  assign tmp40272 = s2 ? tmp40273 : tmp40275;
  assign tmp40271 = s3 ? tmp40272 : tmp39997;
  assign tmp40278 = ~(l1 ? tmp39429 : tmp39388);
  assign tmp40277 = s2 ? tmp39670 : tmp40278;
  assign tmp40276 = s3 ? tmp40277 : tmp40003;
  assign tmp40270 = s4 ? tmp40271 : tmp40276;
  assign tmp40244 = s5 ? tmp40245 : tmp40270;
  assign tmp40207 = s6 ? tmp40208 : tmp40244;
  assign tmp40206 = s7 ? tmp39370 : tmp40207;
  assign tmp40284 = l1 ? tmp39460 : tmp39435;
  assign tmp40286 = l1 ? tmp39385 : tmp40214;
  assign tmp40287 = ~(l1 ? tmp40014 : tmp39435);
  assign tmp40285 = ~(s0 ? tmp40286 : tmp40287);
  assign tmp40283 = s1 ? tmp40284 : tmp40285;
  assign tmp40291 = l1 ? tmp39972 : tmp39381;
  assign tmp40292 = ~(l1 ? tmp39925 : tmp39604);
  assign tmp40290 = s0 ? tmp40291 : tmp40292;
  assign tmp40294 = l1 ? tmp39972 : tmp40222;
  assign tmp40293 = s0 ? tmp40294 : tmp40292;
  assign tmp40289 = s1 ? tmp40290 : tmp40293;
  assign tmp40296 = s0 ? tmp40294 : tmp40225;
  assign tmp40298 = l1 ? tmp39925 : tmp39604;
  assign tmp40299 = ~(l1 ? tmp39972 : tmp40229);
  assign tmp40297 = ~(s0 ? tmp40298 : tmp40299);
  assign tmp40295 = s1 ? tmp40296 : tmp40297;
  assign tmp40288 = ~(s2 ? tmp40289 : tmp40295);
  assign tmp40282 = s3 ? tmp40283 : tmp40288;
  assign tmp40304 = l1 ? tmp39403 : tmp39435;
  assign tmp40303 = s0 ? tmp40304 : tmp40250;
  assign tmp40306 = l1 ? tmp39972 : tmp40229;
  assign tmp40305 = ~(s0 ? tmp40306 : tmp40292);
  assign tmp40302 = s1 ? tmp40303 : tmp40305;
  assign tmp40308 = s0 ? tmp40284 : tmp39420;
  assign tmp40309 = l1 ? tmp39403 : 1;
  assign tmp40307 = s1 ? tmp40308 : tmp40309;
  assign tmp40301 = s2 ? tmp40302 : tmp40307;
  assign tmp40311 = s1 ? tmp40286 : tmp39531;
  assign tmp40313 = s0 ? tmp39603 : tmp40298;
  assign tmp40312 = ~(s1 ? tmp40298 : tmp40313);
  assign tmp40310 = ~(s2 ? tmp40311 : tmp40312);
  assign tmp40300 = s3 ? tmp40301 : tmp40310;
  assign tmp40281 = s4 ? tmp40282 : tmp40300;
  assign tmp40320 = l1 ? tmp40014 : tmp39435;
  assign tmp40319 = s0 ? tmp40320 : tmp40250;
  assign tmp40321 = ~(l1 ? tmp39972 : tmp39381);
  assign tmp40318 = s1 ? tmp40319 : tmp40321;
  assign tmp40324 = ~(l1 ? 1 : tmp39457);
  assign tmp40323 = s0 ? tmp40298 : tmp40324;
  assign tmp40322 = s1 ? tmp40320 : tmp40323;
  assign tmp40317 = s2 ? tmp40318 : tmp40322;
  assign tmp40327 = l1 ? tmp39429 : tmp40222;
  assign tmp40326 = s1 ? tmp40327 : tmp39987;
  assign tmp40330 = l1 ? tmp39972 : tmp39377;
  assign tmp40329 = ~(s0 ? tmp40330 : tmp40061);
  assign tmp40328 = ~(s1 ? tmp39625 : tmp40329);
  assign tmp40325 = ~(s2 ? tmp40326 : tmp40328);
  assign tmp40316 = s3 ? tmp40317 : tmp40325;
  assign tmp40335 = l1 ? tmp39925 : tmp39435;
  assign tmp40334 = s0 ? tmp39635 : tmp40335;
  assign tmp40336 = s0 ? tmp40309 : tmp40068;
  assign tmp40333 = s1 ? tmp40334 : tmp40336;
  assign tmp40337 = ~(l1 ? tmp39972 : tmp39388);
  assign tmp40332 = s2 ? tmp40333 : tmp40337;
  assign tmp40340 = s0 ? tmp40269 : tmp40073;
  assign tmp40339 = s1 ? tmp40340 : tmp39987;
  assign tmp40338 = ~(s2 ? tmp40339 : tmp39650);
  assign tmp40331 = s3 ? tmp40332 : tmp40338;
  assign tmp40315 = s4 ? tmp40316 : tmp40331;
  assign tmp40314 = s5 ? tmp40315 : tmp40270;
  assign tmp40280 = s6 ? tmp40281 : tmp40314;
  assign tmp40279 = s7 ? tmp39370 : tmp40280;
  assign tmp40205 = s8 ? tmp40206 : tmp40279;
  assign tmp40347 = l1 ? tmp39915 : tmp39541;
  assign tmp40346 = s1 ? tmp40347 : tmp40212;
  assign tmp40351 = l1 ? tmp39918 : tmp39457;
  assign tmp40352 = ~(l1 ? tmp39469 : tmp39649);
  assign tmp40350 = s0 ? tmp40351 : tmp40352;
  assign tmp40354 = l1 ? tmp39918 : tmp40214;
  assign tmp40353 = s0 ? tmp40354 : tmp40352;
  assign tmp40349 = s1 ? tmp40350 : tmp40353;
  assign tmp40356 = s0 ? tmp40354 : 0;
  assign tmp40358 = l1 ? tmp39469 : tmp39649;
  assign tmp40360 = ~(l2 ? tmp39378 : tmp39376);
  assign tmp40359 = ~(l1 ? tmp39918 : tmp40360);
  assign tmp40357 = ~(s0 ? tmp40358 : tmp40359);
  assign tmp40355 = s1 ? tmp40356 : tmp40357;
  assign tmp40348 = ~(s2 ? tmp40349 : tmp40355);
  assign tmp40345 = s3 ? tmp40346 : tmp40348;
  assign tmp40365 = l1 ? tmp39918 : tmp40360;
  assign tmp40364 = ~(s0 ? tmp40365 : tmp40352);
  assign tmp40363 = s1 ? tmp40233 : tmp40364;
  assign tmp40367 = s0 ? tmp40347 : tmp39940;
  assign tmp40366 = s1 ? tmp40367 : tmp39520;
  assign tmp40362 = s2 ? tmp40363 : tmp40366;
  assign tmp40369 = s1 ? tmp40213 : tmp39531;
  assign tmp40371 = s0 ? tmp39603 : tmp40358;
  assign tmp40370 = ~(s1 ? tmp40358 : tmp40371);
  assign tmp40368 = ~(s2 ? tmp40369 : tmp40370);
  assign tmp40361 = s3 ? tmp40362 : tmp40368;
  assign tmp40344 = s4 ? tmp40345 : tmp40361;
  assign tmp40377 = ~(l1 ? tmp39918 : tmp39457);
  assign tmp40376 = s1 ? tmp40249 : tmp40377;
  assign tmp40379 = s0 ? tmp40358 : tmp39583;
  assign tmp40378 = s1 ? tmp39546 : tmp40379;
  assign tmp40375 = s2 ? tmp40376 : tmp40378;
  assign tmp40382 = l1 ? tmp39375 : tmp40214;
  assign tmp40381 = s1 ? tmp40382 : tmp39987;
  assign tmp40380 = ~(s2 ? tmp40381 : tmp40257);
  assign tmp40374 = s3 ? tmp40375 : tmp40380;
  assign tmp40373 = s4 ? tmp40374 : tmp40260;
  assign tmp40372 = s5 ? tmp40373 : tmp40270;
  assign tmp40343 = s6 ? tmp40344 : tmp40372;
  assign tmp40342 = s7 ? tmp39370 : tmp40343;
  assign tmp40341 = s8 ? tmp40279 : tmp40342;
  assign tmp40204 = s9 ? tmp40205 : tmp40341;
  assign tmp40391 = s0 ? tmp40221 : 0;
  assign tmp40390 = s1 ? tmp40391 : tmp40226;
  assign tmp40389 = ~(s2 ? tmp40217 : tmp40390);
  assign tmp40388 = s3 ? tmp40210 : tmp40389;
  assign tmp40395 = s0 ? tmp40211 : tmp39940;
  assign tmp40394 = s1 ? tmp40395 : tmp39520;
  assign tmp40393 = s2 ? tmp40232 : tmp40394;
  assign tmp40396 = ~(s2 ? tmp40369 : tmp40242);
  assign tmp40392 = s3 ? tmp40393 : tmp40396;
  assign tmp40387 = s4 ? tmp40388 : tmp40392;
  assign tmp40386 = s6 ? tmp40387 : tmp40244;
  assign tmp40385 = s7 ? tmp39370 : tmp40386;
  assign tmp40384 = s8 ? tmp40385 : tmp39370;
  assign tmp40401 = s3 ? tmp40231 : tmp40396;
  assign tmp40400 = s4 ? tmp40209 : tmp40401;
  assign tmp40399 = s6 ? tmp40400 : tmp40244;
  assign tmp40398 = s7 ? tmp40399 : tmp40343;
  assign tmp40402 = s7 ? tmp40280 : tmp40386;
  assign tmp40397 = s8 ? tmp40398 : tmp40402;
  assign tmp40383 = s9 ? tmp40384 : tmp40397;
  assign tmp40203 = s10 ? tmp40204 : tmp40383;
  assign tmp40406 = s7 ? tmp40207 : tmp40343;
  assign tmp40405 = s8 ? tmp40406 : tmp40402;
  assign tmp40404 = s9 ? tmp40384 : tmp40405;
  assign tmp40403 = s10 ? tmp40204 : tmp40404;
  assign tmp40202 = s11 ? tmp40203 : tmp40403;
  assign tmp39904 = s12 ? tmp39905 : tmp40202;
  assign tmp39364 = s13 ? tmp39365 : tmp39904;
  assign tmp40419 = l2 ? tmp39378 : tmp39398;
  assign tmp40418 = l1 ? tmp40419 : tmp39801;
  assign tmp40421 = l1 ? tmp39402 : tmp39918;
  assign tmp40423 = l2 ? 1 : 0;
  assign tmp40422 = ~(l1 ? tmp40423 : tmp39801);
  assign tmp40420 = ~(s0 ? tmp40421 : tmp40422);
  assign tmp40417 = s1 ? tmp40418 : tmp40420;
  assign tmp40427 = l1 ? tmp39375 : tmp39384;
  assign tmp40428 = ~(l1 ? tmp39408 : tmp39926);
  assign tmp40426 = s0 ? tmp40427 : tmp40428;
  assign tmp40429 = s0 ? tmp39966 : tmp40428;
  assign tmp40425 = s1 ? tmp40426 : tmp40429;
  assign tmp40432 = ~(l1 ? tmp39385 : tmp39404);
  assign tmp40431 = s0 ? tmp39966 : tmp40432;
  assign tmp40434 = l1 ? tmp39408 : tmp39926;
  assign tmp40435 = ~(l1 ? tmp39375 : tmp39934);
  assign tmp40433 = ~(s0 ? tmp40434 : tmp40435);
  assign tmp40430 = s1 ? tmp40431 : tmp40433;
  assign tmp40424 = ~(s2 ? tmp40425 : tmp40430);
  assign tmp40416 = s3 ? tmp40417 : tmp40424;
  assign tmp40440 = l1 ? tmp39384 : tmp39801;
  assign tmp40439 = s0 ? tmp40440 : tmp39424;
  assign tmp40442 = l1 ? tmp39375 : tmp39934;
  assign tmp40441 = ~(s0 ? tmp40442 : tmp40428);
  assign tmp40438 = s1 ? tmp40439 : tmp40441;
  assign tmp40444 = s0 ? tmp40418 : tmp39424;
  assign tmp40445 = l1 ? tmp39384 : tmp39478;
  assign tmp40443 = s1 ? tmp40444 : tmp40445;
  assign tmp40437 = s2 ? tmp40438 : tmp40443;
  assign tmp40447 = s1 ? tmp40421 : tmp39531;
  assign tmp40449 = s0 ? tmp40434 : tmp39932;
  assign tmp40450 = s0 ? tmp39603 : tmp40434;
  assign tmp40448 = ~(s1 ? tmp40449 : tmp40450);
  assign tmp40446 = ~(s2 ? tmp40447 : tmp40448);
  assign tmp40436 = s3 ? tmp40437 : tmp40446;
  assign tmp40415 = s4 ? tmp40416 : tmp40436;
  assign tmp40457 = l1 ? tmp40423 : tmp39801;
  assign tmp40456 = s0 ? tmp40457 : tmp39452;
  assign tmp40458 = ~(l1 ? tmp39375 : tmp39384);
  assign tmp40455 = s1 ? tmp40456 : tmp40458;
  assign tmp40459 = s1 ? tmp40457 : tmp40172;
  assign tmp40454 = s2 ? tmp40455 : tmp40459;
  assign tmp40463 = l1 ? tmp39375 : tmp39840;
  assign tmp40462 = ~(s0 ? tmp40463 : tmp40127);
  assign tmp40461 = ~(s1 ? tmp39625 : tmp40462);
  assign tmp40460 = ~(s2 ? tmp39964 : tmp40461);
  assign tmp40453 = s3 ? tmp40454 : tmp40460;
  assign tmp40468 = l1 ? tmp39408 : tmp39801;
  assign tmp40467 = s0 ? tmp39635 : tmp40468;
  assign tmp40469 = s0 ? tmp40445 : tmp39980;
  assign tmp40466 = s1 ? tmp40467 : tmp40469;
  assign tmp40470 = ~(l1 ? tmp39375 : tmp39621);
  assign tmp40465 = s2 ? tmp40466 : tmp40470;
  assign tmp40464 = s3 ? tmp40465 : tmp39982;
  assign tmp40452 = s4 ? tmp40453 : tmp40464;
  assign tmp40451 = s5 ? tmp40452 : tmp39988;
  assign tmp40414 = s6 ? tmp40415 : tmp40451;
  assign tmp40413 = s7 ? tmp39370 : tmp40414;
  assign tmp40477 = ~(l2 ? tmp39379 : tmp39398);
  assign tmp40476 = l1 ? tmp40419 : tmp40477;
  assign tmp40479 = l1 ? tmp39402 : tmp39972;
  assign tmp40480 = ~(l1 ? tmp40423 : tmp40477);
  assign tmp40478 = ~(s0 ? tmp40479 : tmp40480);
  assign tmp40475 = s1 ? tmp40476 : tmp40478;
  assign tmp40484 = l1 ? tmp39375 : tmp39587;
  assign tmp40483 = s0 ? tmp40484 : tmp40428;
  assign tmp40482 = s1 ? tmp40426 : tmp40483;
  assign tmp40486 = s0 ? tmp40484 : tmp40432;
  assign tmp40489 = l2 ? tmp39430 : tmp39398;
  assign tmp40488 = ~(l1 ? tmp39375 : tmp40489);
  assign tmp40487 = ~(s0 ? tmp40434 : tmp40488);
  assign tmp40485 = s1 ? tmp40486 : tmp40487;
  assign tmp40481 = ~(s2 ? tmp40482 : tmp40485);
  assign tmp40474 = s3 ? tmp40475 : tmp40481;
  assign tmp40494 = l1 ? tmp39384 : tmp40477;
  assign tmp40493 = s0 ? tmp40494 : tmp39424;
  assign tmp40496 = l1 ? tmp39375 : tmp40489;
  assign tmp40495 = ~(s0 ? tmp40496 : tmp40428);
  assign tmp40492 = s1 ? tmp40493 : tmp40495;
  assign tmp40498 = s0 ? tmp40476 : tmp39424;
  assign tmp40499 = l1 ? tmp39384 : tmp39404;
  assign tmp40497 = s1 ? tmp40498 : tmp40499;
  assign tmp40491 = s2 ? tmp40492 : tmp40497;
  assign tmp40501 = s1 ? tmp40479 : tmp39531;
  assign tmp40503 = s0 ? tmp40434 : tmp39993;
  assign tmp40506 = l2 ? tmp39460 : tmp39430;
  assign tmp40505 = l1 ? tmp39434 : tmp40506;
  assign tmp40504 = s0 ? tmp40505 : tmp40434;
  assign tmp40502 = ~(s1 ? tmp40503 : tmp40504);
  assign tmp40500 = ~(s2 ? tmp40501 : tmp40502);
  assign tmp40490 = s3 ? tmp40491 : tmp40500;
  assign tmp40473 = s4 ? tmp40474 : tmp40490;
  assign tmp40513 = l1 ? tmp40423 : tmp40477;
  assign tmp40512 = s0 ? tmp40513 : tmp39452;
  assign tmp40511 = s1 ? tmp40512 : tmp40458;
  assign tmp40515 = s0 ? tmp39993 : tmp39424;
  assign tmp40514 = s1 ? tmp40513 : tmp40515;
  assign tmp40510 = s2 ? tmp40511 : tmp40514;
  assign tmp40517 = s1 ? tmp40484 : tmp39968;
  assign tmp40519 = s0 ? tmp40505 : tmp39626;
  assign tmp40520 = ~(l1 ? tmp39375 : tmp39840);
  assign tmp40518 = ~(s1 ? tmp40519 : tmp40520);
  assign tmp40516 = ~(s2 ? tmp40517 : tmp40518);
  assign tmp40509 = s3 ? tmp40510 : tmp40516;
  assign tmp40525 = l1 ? tmp39408 : tmp40477;
  assign tmp40524 = s0 ? tmp39635 : tmp40525;
  assign tmp40527 = ~(l1 ? tmp39402 : tmp39429);
  assign tmp40526 = s0 ? tmp40445 : tmp40527;
  assign tmp40523 = s1 ? tmp40524 : tmp40526;
  assign tmp40528 = ~(l1 ? tmp39375 : tmp39630);
  assign tmp40522 = s2 ? tmp40523 : tmp40528;
  assign tmp40532 = l1 ? tmp39429 : tmp39630;
  assign tmp40534 = l2 ? tmp39403 : tmp39430;
  assign tmp40533 = ~(l1 ? tmp39915 : tmp40534);
  assign tmp40531 = s0 ? tmp40532 : tmp40533;
  assign tmp40530 = s1 ? tmp40531 : tmp39987;
  assign tmp40529 = ~(s2 ? tmp40530 : tmp39650);
  assign tmp40521 = s3 ? tmp40522 : tmp40529;
  assign tmp40508 = s4 ? tmp40509 : tmp40521;
  assign tmp40539 = ~(l2 ? tmp39430 : 1);
  assign tmp40538 = s1 ? tmp39992 : tmp40539;
  assign tmp40537 = s2 ? tmp40538 : tmp39994;
  assign tmp40536 = s3 ? tmp40537 : tmp39997;
  assign tmp40542 = s1 ? tmp39671 : tmp40505;
  assign tmp40541 = s2 ? tmp40542 : tmp39999;
  assign tmp40540 = s3 ? tmp40541 : tmp40003;
  assign tmp40535 = s4 ? tmp40536 : tmp40540;
  assign tmp40507 = s5 ? tmp40508 : tmp40535;
  assign tmp40472 = s6 ? tmp40473 : tmp40507;
  assign tmp40471 = s7 ? tmp39370 : tmp40472;
  assign tmp40412 = s8 ? tmp40413 : tmp40471;
  assign tmp40549 = l1 ? tmp40419 : tmp39615;
  assign tmp40551 = ~(l1 ? tmp40423 : tmp39615);
  assign tmp40550 = ~(s0 ? tmp40479 : tmp40551);
  assign tmp40548 = s1 ? tmp40549 : tmp40550;
  assign tmp40555 = l1 ? tmp39375 : tmp39385;
  assign tmp40556 = ~(l1 ? tmp39408 : tmp39623);
  assign tmp40554 = s0 ? tmp40555 : tmp40556;
  assign tmp40558 = l1 ? tmp39375 : tmp39972;
  assign tmp40557 = s0 ? tmp40558 : tmp40556;
  assign tmp40553 = s1 ? tmp40554 : tmp40557;
  assign tmp40560 = s0 ? tmp40558 : tmp40432;
  assign tmp40562 = l1 ? tmp39408 : tmp39623;
  assign tmp40564 = l2 ? tmp39430 : tmp39616;
  assign tmp40563 = ~(l1 ? tmp39375 : tmp40564);
  assign tmp40561 = ~(s0 ? tmp40562 : tmp40563);
  assign tmp40559 = s1 ? tmp40560 : tmp40561;
  assign tmp40552 = ~(s2 ? tmp40553 : tmp40559);
  assign tmp40547 = s3 ? tmp40548 : tmp40552;
  assign tmp40569 = l1 ? tmp39384 : tmp39615;
  assign tmp40568 = s0 ? tmp40569 : tmp39424;
  assign tmp40571 = l1 ? tmp39375 : tmp40564;
  assign tmp40570 = ~(s0 ? tmp40571 : tmp40556);
  assign tmp40567 = s1 ? tmp40568 : tmp40570;
  assign tmp40573 = s0 ? tmp40549 : tmp39424;
  assign tmp40572 = s1 ? tmp40573 : tmp40499;
  assign tmp40566 = s2 ? tmp40567 : tmp40572;
  assign tmp40577 = l1 ? tmp39469 : tmp39623;
  assign tmp40576 = s0 ? tmp40562 : tmp40577;
  assign tmp40578 = s0 ? tmp40505 : tmp40562;
  assign tmp40575 = ~(s1 ? tmp40576 : tmp40578);
  assign tmp40574 = ~(s2 ? tmp40501 : tmp40575);
  assign tmp40565 = s3 ? tmp40566 : tmp40574;
  assign tmp40546 = s4 ? tmp40547 : tmp40565;
  assign tmp40585 = l1 ? tmp40423 : tmp39615;
  assign tmp40584 = s0 ? tmp40585 : tmp39452;
  assign tmp40586 = ~(l1 ? tmp39375 : tmp39385);
  assign tmp40583 = s1 ? tmp40584 : tmp40586;
  assign tmp40588 = s0 ? tmp40577 : tmp39424;
  assign tmp40587 = s1 ? tmp40585 : tmp40588;
  assign tmp40582 = s2 ? tmp40583 : tmp40587;
  assign tmp40591 = ~(l1 ? tmp39469 : tmp39623);
  assign tmp40590 = s1 ? tmp40558 : tmp40591;
  assign tmp40593 = ~(l1 ? tmp39375 : tmp39532);
  assign tmp40592 = ~(s1 ? tmp40519 : tmp40593);
  assign tmp40589 = ~(s2 ? tmp40590 : tmp40592);
  assign tmp40581 = s3 ? tmp40582 : tmp40589;
  assign tmp40596 = ~(l1 ? tmp39375 : tmp39429);
  assign tmp40595 = s2 ? tmp40523 : tmp40596;
  assign tmp40599 = s0 ? tmp39429 : tmp40533;
  assign tmp40598 = s1 ? tmp40599 : tmp39987;
  assign tmp40597 = ~(s2 ? tmp40598 : tmp39650);
  assign tmp40594 = s3 ? tmp40595 : tmp40597;
  assign tmp40580 = s4 ? tmp40581 : tmp40594;
  assign tmp40604 = s0 ? tmp40577 : 0;
  assign tmp40603 = s1 ? tmp40604 : tmp40539;
  assign tmp40606 = l1 ? tmp39480 : tmp39518;
  assign tmp40605 = s1 ? tmp40606 : tmp39996;
  assign tmp40602 = s2 ? tmp40603 : tmp40605;
  assign tmp40601 = s3 ? tmp40602 : tmp39997;
  assign tmp40608 = s2 ? tmp40542 : tmp40539;
  assign tmp40607 = s3 ? tmp40608 : tmp40003;
  assign tmp40600 = s4 ? tmp40601 : tmp40607;
  assign tmp40579 = s5 ? tmp40580 : tmp40600;
  assign tmp40545 = s6 ? tmp40546 : tmp40579;
  assign tmp40544 = s7 ? tmp39370 : tmp40545;
  assign tmp40543 = s8 ? tmp40471 : tmp40544;
  assign tmp40411 = s9 ? tmp40412 : tmp40543;
  assign tmp40610 = s8 ? tmp40471 : tmp39370;
  assign tmp40617 = ~(s2 ? tmp40174 : tmp40461);
  assign tmp40616 = s3 ? tmp40454 : tmp40617;
  assign tmp40615 = s4 ? tmp40616 : tmp40464;
  assign tmp40614 = s5 ? tmp40615 : tmp39988;
  assign tmp40613 = s6 ? tmp40415 : tmp40614;
  assign tmp40612 = s7 ? tmp40613 : tmp40545;
  assign tmp40611 = s8 ? tmp40612 : tmp40472;
  assign tmp40609 = s9 ? tmp40610 : tmp40611;
  assign tmp40410 = s10 ? tmp40411 : tmp40609;
  assign tmp40621 = s7 ? tmp40414 : tmp40545;
  assign tmp40620 = s8 ? tmp40621 : tmp40472;
  assign tmp40619 = s9 ? tmp40610 : tmp40620;
  assign tmp40618 = s10 ? tmp40411 : tmp40619;
  assign tmp40409 = s11 ? tmp40410 : tmp40618;
  assign tmp40632 = l2 ? tmp39378 : tmp39616;
  assign tmp40634 = ~(l3 ? tmp39379 : 1);
  assign tmp40633 = l2 ? tmp39376 : tmp40634;
  assign tmp40631 = l1 ? tmp40632 : tmp40633;
  assign tmp40637 = l2 ? 1 : tmp39389;
  assign tmp40636 = ~(l1 ? tmp40637 : tmp40633);
  assign tmp40635 = ~(s0 ? tmp39946 : tmp40636);
  assign tmp40630 = s1 ? tmp40631 : tmp40635;
  assign tmp40640 = l1 ? tmp39621 : tmp39478;
  assign tmp40642 = l2 ? tmp39378 : tmp39389;
  assign tmp40643 = l2 ? tmp39440 : tmp40634;
  assign tmp40641 = ~(l1 ? tmp40642 : tmp40643);
  assign tmp40639 = s0 ? tmp40640 : tmp40641;
  assign tmp40645 = s0 ? tmp40640 : tmp39420;
  assign tmp40647 = l1 ? tmp40642 : tmp40643;
  assign tmp40649 = ~(l2 ? tmp39440 : tmp40634);
  assign tmp40648 = ~(l1 ? tmp39621 : tmp40649);
  assign tmp40646 = ~(s0 ? tmp40647 : tmp40648);
  assign tmp40644 = s1 ? tmp40645 : tmp40646;
  assign tmp40638 = ~(s2 ? tmp40639 : tmp40644);
  assign tmp40629 = s3 ? tmp40630 : tmp40638;
  assign tmp40654 = l1 ? tmp39385 : tmp40633;
  assign tmp40655 = ~(l1 ? tmp39480 : tmp39478);
  assign tmp40653 = s0 ? tmp40654 : tmp40655;
  assign tmp40657 = l1 ? tmp39621 : tmp40649;
  assign tmp40656 = ~(s0 ? tmp40657 : tmp40641);
  assign tmp40652 = s1 ? tmp40653 : tmp40656;
  assign tmp40659 = s0 ? tmp40631 : tmp40225;
  assign tmp40660 = l1 ? tmp39785 : tmp39375;
  assign tmp40658 = s1 ? tmp40659 : tmp40660;
  assign tmp40651 = s2 ? tmp40652 : tmp40658;
  assign tmp40662 = s1 ? tmp39946 : tmp39651;
  assign tmp40665 = l1 ? tmp39577 : tmp40643;
  assign tmp40664 = s0 ? tmp40647 : tmp40665;
  assign tmp40668 = l2 ? tmp39440 : tmp39430;
  assign tmp40667 = l1 ? tmp39434 : tmp40668;
  assign tmp40666 = s0 ? tmp40667 : tmp40647;
  assign tmp40663 = ~(s1 ? tmp40664 : tmp40666);
  assign tmp40661 = ~(s2 ? tmp40662 : tmp40663);
  assign tmp40650 = s3 ? tmp40651 : tmp40661;
  assign tmp40628 = s4 ? tmp40629 : tmp40650;
  assign tmp40675 = l1 ? tmp40637 : tmp40633;
  assign tmp40674 = s0 ? tmp40675 : tmp40096;
  assign tmp40676 = ~(l1 ? tmp39621 : tmp39478);
  assign tmp40673 = s1 ? tmp40674 : tmp40676;
  assign tmp40678 = l1 ? tmp40637 : tmp39376;
  assign tmp40679 = s0 ? tmp40665 : tmp39401;
  assign tmp40677 = s1 ? tmp40678 : tmp40679;
  assign tmp40672 = s2 ? tmp40673 : tmp40677;
  assign tmp40683 = l2 ? tmp39440 : tmp39376;
  assign tmp40682 = ~(l1 ? tmp39434 : tmp40683);
  assign tmp40681 = s1 ? tmp40640 : tmp40682;
  assign tmp40685 = s0 ? tmp40667 : tmp39626;
  assign tmp40687 = l1 ? tmp39630 : tmp39513;
  assign tmp40686 = ~(s0 ? tmp40657 : tmp40687);
  assign tmp40684 = ~(s1 ? tmp40685 : tmp40686);
  assign tmp40680 = ~(s2 ? tmp40681 : tmp40684);
  assign tmp40671 = s3 ? tmp40672 : tmp40680;
  assign tmp40693 = l2 ? tmp39379 : tmp39430;
  assign tmp40692 = l1 ? tmp39378 : tmp40693;
  assign tmp40694 = l1 ? tmp40642 : tmp39376;
  assign tmp40691 = s0 ? tmp40692 : tmp40694;
  assign tmp40696 = l1 ? tmp39785 : 1;
  assign tmp40695 = s0 ? tmp40696 : tmp39479;
  assign tmp40690 = s1 ? tmp40691 : tmp40695;
  assign tmp40697 = ~(s1 ? tmp39495 : tmp40640);
  assign tmp40689 = s2 ? tmp40690 : tmp40697;
  assign tmp40701 = l1 ? tmp39630 : tmp39478;
  assign tmp40702 = ~(l1 ? tmp39378 : tmp39376);
  assign tmp40700 = s0 ? tmp40701 : tmp40702;
  assign tmp40705 = l2 ? tmp39379 : tmp39376;
  assign tmp40704 = ~(l1 ? tmp39434 : tmp40705);
  assign tmp40703 = s0 ? tmp39495 : tmp40704;
  assign tmp40699 = s1 ? tmp40700 : tmp40703;
  assign tmp40698 = ~(s2 ? tmp40699 : tmp39651);
  assign tmp40688 = s3 ? tmp40689 : tmp40698;
  assign tmp40670 = s4 ? tmp40671 : tmp40688;
  assign tmp40711 = l1 ? tmp39434 : tmp40683;
  assign tmp40710 = s0 ? tmp40711 : 0;
  assign tmp40709 = s1 ? tmp40710 : tmp39521;
  assign tmp40713 = l1 ? 1 : tmp39480;
  assign tmp40712 = s1 ? tmp40713 : tmp39661;
  assign tmp40708 = s2 ? tmp40709 : tmp40712;
  assign tmp40716 = l1 ? tmp39378 : tmp39430;
  assign tmp40715 = ~(s1 ? tmp40716 : tmp39661);
  assign tmp40714 = ~(s2 ? tmp39663 : tmp40715);
  assign tmp40707 = s3 ? tmp40708 : tmp40714;
  assign tmp40719 = s1 ? tmp39671 : tmp40667;
  assign tmp40720 = ~(l1 ? tmp39630 : tmp39478);
  assign tmp40718 = s2 ? tmp40719 : tmp40720;
  assign tmp40722 = ~(l1 ? tmp39630 : tmp39513);
  assign tmp40721 = s1 ? tmp39673 : tmp40722;
  assign tmp40717 = s3 ? tmp40718 : tmp40721;
  assign tmp40706 = s4 ? tmp40707 : tmp40717;
  assign tmp40669 = s5 ? tmp40670 : tmp40706;
  assign tmp40627 = s6 ? tmp40628 : tmp40669;
  assign tmp40626 = s7 ? tmp39370 : tmp40627;
  assign tmp40729 = l2 ? tmp39430 : tmp40634;
  assign tmp40728 = l1 ? tmp40632 : tmp40729;
  assign tmp40731 = l1 ? tmp39403 : tmp39404;
  assign tmp40732 = ~(l1 ? tmp40637 : tmp40729);
  assign tmp40730 = ~(s0 ? tmp40731 : tmp40732);
  assign tmp40727 = s1 ? tmp40728 : tmp40730;
  assign tmp40735 = l1 ? tmp39621 : tmp39404;
  assign tmp40737 = l2 ? tmp39379 : tmp40634;
  assign tmp40736 = ~(l1 ? tmp40642 : tmp40737);
  assign tmp40734 = s0 ? tmp40735 : tmp40736;
  assign tmp40739 = s0 ? tmp40735 : tmp39420;
  assign tmp40741 = l1 ? tmp40642 : tmp40737;
  assign tmp40743 = ~(l2 ? tmp39379 : tmp40634);
  assign tmp40742 = ~(l1 ? tmp39621 : tmp40743);
  assign tmp40740 = ~(s0 ? tmp40741 : tmp40742);
  assign tmp40738 = s1 ? tmp40739 : tmp40740;
  assign tmp40733 = ~(s2 ? tmp40734 : tmp40738);
  assign tmp40726 = s3 ? tmp40727 : tmp40733;
  assign tmp40748 = l1 ? tmp39385 : tmp40729;
  assign tmp40749 = ~(l1 ? tmp39403 : tmp39478);
  assign tmp40747 = s0 ? tmp40748 : tmp40749;
  assign tmp40751 = l1 ? tmp39621 : tmp40743;
  assign tmp40750 = ~(s0 ? tmp40751 : tmp40736);
  assign tmp40746 = s1 ? tmp40747 : tmp40750;
  assign tmp40753 = s0 ? tmp40728 : tmp40225;
  assign tmp40752 = s1 ? tmp40753 : tmp39428;
  assign tmp40745 = s2 ? tmp40746 : tmp40752;
  assign tmp40755 = s1 ? tmp40731 : tmp39651;
  assign tmp40758 = l1 ? tmp39434 : tmp40737;
  assign tmp40757 = s0 ? tmp40741 : tmp40758;
  assign tmp40760 = l1 ? tmp39434 : tmp40693;
  assign tmp40759 = s0 ? tmp40760 : tmp40741;
  assign tmp40756 = ~(s1 ? tmp40757 : tmp40759);
  assign tmp40754 = ~(s2 ? tmp40755 : tmp40756);
  assign tmp40744 = s3 ? tmp40745 : tmp40754;
  assign tmp40725 = s4 ? tmp40726 : tmp40744;
  assign tmp40767 = l1 ? tmp40637 : tmp40729;
  assign tmp40766 = s0 ? tmp40767 : tmp40096;
  assign tmp40768 = ~(l1 ? tmp39621 : tmp39404);
  assign tmp40765 = s1 ? tmp40766 : tmp40768;
  assign tmp40771 = l2 ? tmp39430 : tmp39376;
  assign tmp40770 = l1 ? tmp40637 : tmp40771;
  assign tmp40772 = s0 ? tmp40758 : tmp39401;
  assign tmp40769 = s1 ? tmp40770 : tmp40772;
  assign tmp40764 = s2 ? tmp40765 : tmp40769;
  assign tmp40774 = s1 ? tmp40735 : tmp40704;
  assign tmp40776 = s0 ? tmp40760 : tmp39626;
  assign tmp40779 = l2 ? tmp39403 : tmp39378;
  assign tmp40778 = l1 ? tmp39621 : tmp40779;
  assign tmp40777 = ~(s0 ? tmp40751 : tmp40778);
  assign tmp40775 = ~(s1 ? tmp40776 : tmp40777);
  assign tmp40773 = ~(s2 ? tmp40774 : tmp40775);
  assign tmp40763 = s3 ? tmp40764 : tmp40773;
  assign tmp40784 = l1 ? tmp40642 : tmp40771;
  assign tmp40783 = s0 ? tmp40692 : tmp40784;
  assign tmp40782 = s1 ? tmp40783 : tmp39482;
  assign tmp40781 = s2 ? tmp40782 : tmp40768;
  assign tmp40788 = l1 ? tmp39630 : tmp39404;
  assign tmp40789 = ~(l1 ? tmp39378 : tmp40771);
  assign tmp40787 = s0 ? tmp40788 : tmp40789;
  assign tmp40786 = s1 ? tmp40787 : tmp40704;
  assign tmp40785 = ~(s2 ? tmp40786 : tmp39651);
  assign tmp40780 = s3 ? tmp40781 : tmp40785;
  assign tmp40762 = s4 ? tmp40763 : tmp40780;
  assign tmp40795 = l1 ? tmp39434 : tmp40705;
  assign tmp40794 = s0 ? tmp40795 : 0;
  assign tmp40796 = ~(l1 ? tmp39429 : tmp39402);
  assign tmp40793 = s1 ? tmp40794 : tmp40796;
  assign tmp40792 = s2 ? tmp40793 : tmp40712;
  assign tmp40791 = s3 ? tmp40792 : tmp40714;
  assign tmp40799 = s1 ? tmp39671 : tmp40760;
  assign tmp40800 = ~(l1 ? tmp39630 : tmp39404);
  assign tmp40798 = s2 ? tmp40799 : tmp40800;
  assign tmp40797 = s3 ? tmp40798 : tmp40721;
  assign tmp40790 = s4 ? tmp40791 : tmp40797;
  assign tmp40761 = s5 ? tmp40762 : tmp40790;
  assign tmp40724 = s6 ? tmp40725 : tmp40761;
  assign tmp40723 = s7 ? tmp39370 : tmp40724;
  assign tmp40625 = s8 ? tmp40626 : tmp40723;
  assign tmp40624 = s9 ? tmp40625 : tmp40723;
  assign tmp40802 = s8 ? tmp40723 : tmp39370;
  assign tmp40810 = s1 ? tmp40700 : tmp40704;
  assign tmp40809 = ~(s2 ? tmp40810 : tmp39651);
  assign tmp40808 = s3 ? tmp40689 : tmp40809;
  assign tmp40807 = s4 ? tmp40671 : tmp40808;
  assign tmp40806 = s5 ? tmp40807 : tmp40706;
  assign tmp40805 = s6 ? tmp40628 : tmp40806;
  assign tmp40816 = l2 ? tmp39430 : tmp39380;
  assign tmp40815 = l1 ? tmp40632 : tmp40816;
  assign tmp40818 = ~(l1 ? tmp40637 : tmp40816);
  assign tmp40817 = ~(s0 ? tmp40731 : tmp40818);
  assign tmp40814 = s1 ? tmp40815 : tmp40817;
  assign tmp40821 = l1 ? tmp39621 : tmp39518;
  assign tmp40823 = l2 ? tmp39379 : tmp39380;
  assign tmp40822 = ~(l1 ? tmp40642 : tmp40823);
  assign tmp40820 = s0 ? tmp40821 : tmp40822;
  assign tmp40825 = s0 ? tmp40821 : tmp39420;
  assign tmp40827 = l1 ? tmp40642 : tmp40823;
  assign tmp40829 = ~(l2 ? tmp39379 : tmp39380);
  assign tmp40828 = ~(l1 ? tmp39621 : tmp40829);
  assign tmp40826 = ~(s0 ? tmp40827 : tmp40828);
  assign tmp40824 = s1 ? tmp40825 : tmp40826;
  assign tmp40819 = ~(s2 ? tmp40820 : tmp40824);
  assign tmp40813 = s3 ? tmp40814 : tmp40819;
  assign tmp40834 = l1 ? tmp39385 : tmp40816;
  assign tmp40833 = s0 ? tmp40834 : tmp40749;
  assign tmp40836 = l1 ? tmp39621 : tmp40829;
  assign tmp40835 = ~(s0 ? tmp40836 : tmp40822);
  assign tmp40832 = s1 ? tmp40833 : tmp40835;
  assign tmp40838 = s0 ? tmp40815 : tmp40225;
  assign tmp40837 = s1 ? tmp40838 : tmp39428;
  assign tmp40831 = s2 ? tmp40832 : tmp40837;
  assign tmp40842 = l1 ? tmp39434 : tmp40823;
  assign tmp40841 = s0 ? tmp40827 : tmp40842;
  assign tmp40843 = s0 ? tmp40760 : tmp40827;
  assign tmp40840 = ~(s1 ? tmp40841 : tmp40843);
  assign tmp40839 = ~(s2 ? tmp40755 : tmp40840);
  assign tmp40830 = s3 ? tmp40831 : tmp40839;
  assign tmp40812 = s4 ? tmp40813 : tmp40830;
  assign tmp40850 = l1 ? tmp40637 : tmp40816;
  assign tmp40849 = s0 ? tmp40850 : tmp40096;
  assign tmp40851 = ~(l1 ? tmp39621 : tmp39518);
  assign tmp40848 = s1 ? tmp40849 : tmp40851;
  assign tmp40853 = l1 ? tmp40637 : tmp39430;
  assign tmp40854 = s0 ? tmp40842 : tmp39401;
  assign tmp40852 = s1 ? tmp40853 : tmp40854;
  assign tmp40847 = s2 ? tmp40848 : tmp40852;
  assign tmp40857 = ~(l1 ? tmp39434 : tmp40693);
  assign tmp40856 = s1 ? tmp40821 : tmp40857;
  assign tmp40861 = l2 ? tmp39403 : tmp39460;
  assign tmp40860 = l1 ? tmp39621 : tmp40861;
  assign tmp40859 = ~(s0 ? tmp40836 : tmp40860);
  assign tmp40858 = ~(s1 ? tmp40776 : tmp40859);
  assign tmp40855 = ~(s2 ? tmp40856 : tmp40858);
  assign tmp40846 = s3 ? tmp40847 : tmp40855;
  assign tmp40866 = l1 ? tmp40642 : tmp39430;
  assign tmp40865 = s0 ? tmp40692 : tmp40866;
  assign tmp40864 = s1 ? tmp40865 : tmp39482;
  assign tmp40863 = s2 ? tmp40864 : tmp40851;
  assign tmp40870 = l1 ? tmp39630 : tmp39518;
  assign tmp40871 = ~(l1 ? tmp39378 : tmp39430);
  assign tmp40869 = s0 ? tmp40870 : tmp40871;
  assign tmp40868 = s1 ? tmp40869 : tmp40857;
  assign tmp40867 = ~(s2 ? tmp40868 : tmp39651);
  assign tmp40862 = s3 ? tmp40863 : tmp40867;
  assign tmp40845 = s4 ? tmp40846 : tmp40862;
  assign tmp40876 = s0 ? tmp40760 : 0;
  assign tmp40875 = s1 ? tmp40876 : tmp40796;
  assign tmp40877 = s1 ? 1 : tmp39661;
  assign tmp40874 = s2 ? tmp40875 : tmp40877;
  assign tmp40880 = ~(l1 ? tmp39630 : tmp39480);
  assign tmp40879 = ~(s1 ? tmp40716 : tmp40880);
  assign tmp40878 = ~(s2 ? tmp39663 : tmp40879);
  assign tmp40873 = s3 ? tmp40874 : tmp40878;
  assign tmp40883 = ~(l1 ? tmp39630 : tmp39518);
  assign tmp40882 = s2 ? tmp40799 : tmp40883;
  assign tmp40885 = ~(l1 ? tmp39630 : tmp39459);
  assign tmp40884 = s1 ? tmp39673 : tmp40885;
  assign tmp40881 = s3 ? tmp40882 : tmp40884;
  assign tmp40872 = s4 ? tmp40873 : tmp40881;
  assign tmp40844 = s5 ? tmp40845 : tmp40872;
  assign tmp40811 = s6 ? tmp40812 : tmp40844;
  assign tmp40804 = s7 ? tmp40805 : tmp40811;
  assign tmp40803 = s8 ? tmp40804 : tmp40724;
  assign tmp40801 = s9 ? tmp40802 : tmp40803;
  assign tmp40623 = s10 ? tmp40624 : tmp40801;
  assign tmp40889 = s7 ? tmp40627 : tmp40811;
  assign tmp40888 = s8 ? tmp40889 : tmp40724;
  assign tmp40887 = s9 ? tmp40802 : tmp40888;
  assign tmp40886 = s10 ? tmp40624 : tmp40887;
  assign tmp40622 = s11 ? tmp40623 : tmp40886;
  assign tmp40408 = s12 ? tmp40409 : tmp40622;
  assign tmp40901 = l2 ? tmp39440 : tmp39616;
  assign tmp40900 = l1 ? tmp40901 : tmp39567;
  assign tmp40903 = l1 ? tmp39480 : tmp39375;
  assign tmp40905 = l2 ? tmp39376 : tmp39389;
  assign tmp40904 = ~(l1 ? tmp40905 : tmp39567);
  assign tmp40902 = ~(s0 ? tmp40903 : tmp40904);
  assign tmp40899 = s1 ? tmp40900 : tmp40902;
  assign tmp40910 = l2 ? tmp39440 : tmp39389;
  assign tmp40909 = ~(l1 ? tmp40910 : tmp39578);
  assign tmp40908 = s0 ? tmp39520 : tmp40909;
  assign tmp40911 = s0 ? tmp40903 : tmp40909;
  assign tmp40907 = s1 ? tmp40908 : tmp40911;
  assign tmp40914 = ~(l1 ? tmp39785 : tmp39457);
  assign tmp40913 = s0 ? tmp40903 : tmp40914;
  assign tmp40916 = l1 ? tmp40910 : tmp39578;
  assign tmp40917 = ~(l1 ? tmp39480 : tmp39588);
  assign tmp40915 = ~(s0 ? tmp40916 : tmp40917);
  assign tmp40912 = s1 ? tmp40913 : tmp40915;
  assign tmp40906 = ~(s2 ? tmp40907 : tmp40912);
  assign tmp40898 = s3 ? tmp40899 : tmp40906;
  assign tmp40922 = l1 ? tmp39918 : tmp39567;
  assign tmp40921 = s0 ? tmp40922 : tmp39479;
  assign tmp40924 = l1 ? tmp39480 : tmp39588;
  assign tmp40923 = ~(s0 ? tmp40924 : tmp40909);
  assign tmp40920 = s1 ? tmp40921 : tmp40923;
  assign tmp40926 = s0 ? tmp40900 : tmp40225;
  assign tmp40927 = l1 ? tmp39785 : tmp39478;
  assign tmp40925 = s1 ? tmp40926 : tmp40927;
  assign tmp40919 = s2 ? tmp40920 : tmp40925;
  assign tmp40929 = s1 ? tmp40903 : tmp39531;
  assign tmp40933 = l2 ? tmp39440 : tmp39379;
  assign tmp40932 = l1 ? tmp40933 : tmp39578;
  assign tmp40931 = s0 ? tmp40916 : tmp40932;
  assign tmp40935 = l1 ? tmp39379 : tmp39604;
  assign tmp40934 = s0 ? tmp40935 : tmp40916;
  assign tmp40930 = ~(s1 ? tmp40931 : tmp40934);
  assign tmp40928 = ~(s2 ? tmp40929 : tmp40930);
  assign tmp40918 = s3 ? tmp40919 : tmp40928;
  assign tmp40897 = s4 ? tmp40898 : tmp40918;
  assign tmp40942 = l1 ? tmp40905 : tmp39567;
  assign tmp40941 = s0 ? tmp40942 : 0;
  assign tmp40940 = s1 ? tmp40941 : tmp39479;
  assign tmp40944 = l1 ? tmp40905 : tmp39615;
  assign tmp40945 = s0 ? tmp40932 : 0;
  assign tmp40943 = s1 ? tmp40944 : tmp40945;
  assign tmp40939 = s2 ? tmp40940 : tmp40943;
  assign tmp40948 = ~(l1 ? tmp39379 : tmp39623);
  assign tmp40947 = s1 ? tmp40903 : tmp40948;
  assign tmp40950 = s0 ? tmp40935 : tmp39626;
  assign tmp40951 = ~(l1 ? tmp39480 : tmp39532);
  assign tmp40949 = ~(s1 ? tmp40950 : tmp40951);
  assign tmp40946 = ~(s2 ? tmp40947 : tmp40949);
  assign tmp40938 = s3 ? tmp40939 : tmp40946;
  assign tmp40956 = l1 ? tmp40910 : tmp39637;
  assign tmp40955 = s0 ? tmp39635 : tmp40956;
  assign tmp40957 = s0 ? tmp40927 : tmp39639;
  assign tmp40954 = s1 ? tmp40955 : tmp40957;
  assign tmp40958 = ~(l1 ? tmp39480 : tmp39429);
  assign tmp40953 = s2 ? tmp40954 : tmp40958;
  assign tmp40962 = l1 ? tmp39480 : tmp39429;
  assign tmp40963 = ~(l1 ? tmp39439 : tmp39541);
  assign tmp40961 = s0 ? tmp40962 : tmp40963;
  assign tmp40964 = ~(l1 ? tmp39379 : tmp39649);
  assign tmp40960 = s1 ? tmp40961 : tmp40964;
  assign tmp40959 = ~(s2 ? tmp40960 : tmp39650);
  assign tmp40952 = s3 ? tmp40953 : tmp40959;
  assign tmp40937 = s4 ? tmp40938 : tmp40952;
  assign tmp40970 = l1 ? tmp39379 : tmp39623;
  assign tmp40969 = s0 ? tmp40970 : 0;
  assign tmp40968 = s1 ? tmp40969 : tmp40068;
  assign tmp40972 = l1 ? tmp39429 : tmp39518;
  assign tmp40973 = ~(s0 ? tmp39520 : tmp39521);
  assign tmp40971 = s1 ? tmp40972 : tmp40973;
  assign tmp40967 = s2 ? tmp40968 : tmp40971;
  assign tmp40976 = s0 ? tmp39480 : tmp39651;
  assign tmp40975 = s1 ? tmp40976 : tmp39664;
  assign tmp40977 = ~(s1 ? tmp39666 : tmp40958);
  assign tmp40974 = ~(s2 ? tmp40975 : tmp40977);
  assign tmp40966 = s3 ? tmp40967 : tmp40974;
  assign tmp40982 = l2 ? tmp39430 : tmp39379;
  assign tmp40981 = l1 ? tmp40982 : tmp39435;
  assign tmp40980 = s1 ? tmp40981 : tmp40935;
  assign tmp40983 = ~(s1 ? tmp40962 : tmp39548);
  assign tmp40979 = s2 ? tmp40980 : tmp40983;
  assign tmp40985 = l1 ? tmp40982 : tmp39604;
  assign tmp40984 = s1 ? tmp40985 : tmp40951;
  assign tmp40978 = s3 ? tmp40979 : tmp40984;
  assign tmp40965 = s4 ? tmp40966 : tmp40978;
  assign tmp40936 = s5 ? tmp40937 : tmp40965;
  assign tmp40896 = s6 ? tmp40897 : tmp40936;
  assign tmp40895 = s7 ? tmp39370 : tmp40896;
  assign tmp40992 = l2 ? tmp39379 : tmp39616;
  assign tmp40993 = ~(l2 ? tmp39379 : tmp39378);
  assign tmp40991 = l1 ? tmp40992 : tmp40993;
  assign tmp40995 = l1 ? tmp39403 : tmp39429;
  assign tmp40997 = l2 ? tmp39430 : tmp39389;
  assign tmp40996 = ~(l1 ? tmp40997 : tmp40993);
  assign tmp40994 = ~(s0 ? tmp40995 : tmp40996);
  assign tmp40990 = s1 ? tmp40991 : tmp40994;
  assign tmp41002 = l2 ? tmp39379 : tmp39389;
  assign tmp41001 = ~(l1 ? tmp41002 : tmp39578);
  assign tmp41000 = s0 ? tmp40309 : tmp41001;
  assign tmp41003 = s0 ? tmp40995 : tmp41001;
  assign tmp40999 = s1 ? tmp41000 : tmp41003;
  assign tmp41006 = ~(l1 ? tmp39385 : tmp39457);
  assign tmp41005 = s0 ? tmp40995 : tmp41006;
  assign tmp41008 = l1 ? tmp41002 : tmp39578;
  assign tmp41009 = ~(l1 ? tmp39403 : tmp39532);
  assign tmp41007 = ~(s0 ? tmp41008 : tmp41009);
  assign tmp41004 = s1 ? tmp41005 : tmp41007;
  assign tmp40998 = ~(s2 ? tmp40999 : tmp41004);
  assign tmp40989 = s3 ? tmp40990 : tmp40998;
  assign tmp41014 = l1 ? tmp39972 : tmp40993;
  assign tmp41015 = ~(l1 ? tmp39403 : 1);
  assign tmp41013 = s0 ? tmp41014 : tmp41015;
  assign tmp41017 = l1 ? tmp39403 : tmp39532;
  assign tmp41016 = ~(s0 ? tmp41017 : tmp41001);
  assign tmp41012 = s1 ? tmp41013 : tmp41016;
  assign tmp41019 = s0 ? tmp40991 : tmp40225;
  assign tmp41020 = l1 ? tmp39385 : tmp39404;
  assign tmp41018 = s1 ? tmp41019 : tmp41020;
  assign tmp41011 = s2 ? tmp41012 : tmp41018;
  assign tmp41022 = s1 ? tmp40995 : tmp39531;
  assign tmp41025 = l1 ? tmp39379 : tmp39578;
  assign tmp41024 = s0 ? tmp41008 : tmp41025;
  assign tmp41027 = l1 ? tmp39379 : tmp40506;
  assign tmp41026 = s0 ? tmp41027 : tmp41008;
  assign tmp41023 = ~(s1 ? tmp41024 : tmp41026);
  assign tmp41021 = ~(s2 ? tmp41022 : tmp41023);
  assign tmp41010 = s3 ? tmp41011 : tmp41021;
  assign tmp40988 = s4 ? tmp40989 : tmp41010;
  assign tmp41034 = l1 ? tmp40997 : tmp40993;
  assign tmp41033 = s0 ? tmp41034 : 0;
  assign tmp41032 = s1 ? tmp41033 : tmp41015;
  assign tmp41036 = l1 ? tmp40997 : tmp39615;
  assign tmp41037 = s0 ? tmp41025 : tmp40225;
  assign tmp41035 = s1 ? tmp41036 : tmp41037;
  assign tmp41031 = s2 ? tmp41032 : tmp41035;
  assign tmp41039 = s1 ? tmp40995 : tmp40948;
  assign tmp41041 = s0 ? tmp41027 : tmp39626;
  assign tmp41040 = ~(s1 ? tmp41041 : tmp41009);
  assign tmp41038 = ~(s2 ? tmp41039 : tmp41040);
  assign tmp41030 = s3 ? tmp41031 : tmp41038;
  assign tmp41046 = l1 ? tmp41002 : tmp39615;
  assign tmp41045 = s0 ? tmp39635 : tmp41046;
  assign tmp41048 = l1 ? tmp39385 : tmp39478;
  assign tmp41049 = ~(l1 ? tmp39403 : tmp39429);
  assign tmp41047 = s0 ? tmp41048 : tmp41049;
  assign tmp41044 = s1 ? tmp41045 : tmp41047;
  assign tmp41043 = s2 ? tmp41044 : tmp41049;
  assign tmp41054 = l2 ? tmp39403 : tmp39376;
  assign tmp41053 = ~(l1 ? tmp39475 : tmp41054);
  assign tmp41052 = s0 ? tmp40962 : tmp41053;
  assign tmp41051 = s1 ? tmp41052 : tmp40964;
  assign tmp41050 = ~(s2 ? tmp41051 : tmp39650);
  assign tmp41042 = s3 ? tmp41043 : tmp41050;
  assign tmp41029 = s4 ? tmp41030 : tmp41042;
  assign tmp41059 = ~(l1 ? 1 : tmp39429);
  assign tmp41058 = s1 ? tmp40969 : tmp41059;
  assign tmp41060 = s1 ? tmp40972 : tmp39479;
  assign tmp41057 = s2 ? tmp41058 : tmp41060;
  assign tmp41056 = s3 ? tmp41057 : tmp40974;
  assign tmp41063 = s1 ? tmp40981 : tmp41027;
  assign tmp41064 = ~(s1 ? tmp40962 : tmp39480);
  assign tmp41062 = s2 ? tmp41063 : tmp41064;
  assign tmp41061 = s3 ? tmp41062 : tmp40984;
  assign tmp41055 = s4 ? tmp41056 : tmp41061;
  assign tmp41028 = s5 ? tmp41029 : tmp41055;
  assign tmp40987 = s6 ? tmp40988 : tmp41028;
  assign tmp40986 = s7 ? tmp39370 : tmp40987;
  assign tmp40894 = s8 ? tmp40895 : tmp40986;
  assign tmp41071 = l1 ? tmp40992 : tmp39755;
  assign tmp41073 = l1 ? tmp39403 : tmp39375;
  assign tmp41074 = ~(l1 ? tmp40997 : tmp39755);
  assign tmp41072 = ~(s0 ? tmp41073 : tmp41074);
  assign tmp41070 = s1 ? tmp41071 : tmp41072;
  assign tmp41078 = ~(l1 ? tmp41002 : tmp39765);
  assign tmp41077 = s0 ? tmp39495 : tmp41078;
  assign tmp41080 = l1 ? tmp39403 : tmp39621;
  assign tmp41079 = s0 ? tmp41080 : tmp41078;
  assign tmp41076 = s1 ? tmp41077 : tmp41079;
  assign tmp41082 = s0 ? tmp41080 : tmp40250;
  assign tmp41084 = l1 ? tmp41002 : tmp39765;
  assign tmp41085 = ~(l1 ? tmp39403 : tmp39493);
  assign tmp41083 = ~(s0 ? tmp41084 : tmp41085);
  assign tmp41081 = s1 ? tmp41082 : tmp41083;
  assign tmp41075 = ~(s2 ? tmp41076 : tmp41081);
  assign tmp41069 = s3 ? tmp41070 : tmp41075;
  assign tmp41090 = l1 ? tmp39972 : tmp39755;
  assign tmp41089 = s0 ? tmp41090 : tmp41015;
  assign tmp41092 = l1 ? tmp39403 : tmp39493;
  assign tmp41091 = ~(s0 ? tmp41092 : tmp41078);
  assign tmp41088 = s1 ? tmp41089 : tmp41091;
  assign tmp41094 = s0 ? tmp41071 : tmp40225;
  assign tmp41093 = s1 ? tmp41094 : tmp41048;
  assign tmp41087 = s2 ? tmp41088 : tmp41093;
  assign tmp41096 = s1 ? tmp41073 : tmp39531;
  assign tmp41099 = l1 ? tmp39379 : tmp39765;
  assign tmp41098 = s0 ? tmp41084 : tmp41099;
  assign tmp41100 = s0 ? tmp40935 : tmp41084;
  assign tmp41097 = ~(s1 ? tmp41098 : tmp41100);
  assign tmp41095 = ~(s2 ? tmp41096 : tmp41097);
  assign tmp41086 = s3 ? tmp41087 : tmp41095;
  assign tmp41068 = s4 ? tmp41069 : tmp41086;
  assign tmp41107 = l1 ? tmp40997 : tmp39755;
  assign tmp41106 = s0 ? tmp41107 : 0;
  assign tmp41105 = s1 ? tmp41106 : tmp39484;
  assign tmp41109 = l1 ? tmp40997 : tmp39801;
  assign tmp41110 = s0 ? tmp41099 : tmp39803;
  assign tmp41108 = s1 ? tmp41109 : tmp41110;
  assign tmp41104 = s2 ? tmp41105 : tmp41108;
  assign tmp41113 = ~(l1 ? tmp39379 : tmp39807);
  assign tmp41112 = s1 ? tmp41080 : tmp41113;
  assign tmp41114 = ~(s1 ? tmp40950 : tmp41085);
  assign tmp41111 = ~(s2 ? tmp41112 : tmp41114);
  assign tmp41103 = s3 ? tmp41104 : tmp41111;
  assign tmp41119 = l1 ? tmp41002 : tmp39801;
  assign tmp41118 = s0 ? tmp39635 : tmp41119;
  assign tmp41120 = s0 ? tmp41048 : tmp39818;
  assign tmp41117 = s1 ? tmp41118 : tmp41120;
  assign tmp41121 = ~(l1 ? tmp39403 : tmp39621);
  assign tmp41116 = s2 ? tmp41117 : tmp41121;
  assign tmp41125 = l1 ? tmp39480 : tmp39621;
  assign tmp41126 = ~(l1 ? tmp39475 : tmp39435);
  assign tmp41124 = s0 ? tmp41125 : tmp41126;
  assign tmp41127 = ~(l1 ? tmp39379 : tmp39604);
  assign tmp41123 = s1 ? tmp41124 : tmp41127;
  assign tmp41122 = ~(s2 ? tmp41123 : tmp39650);
  assign tmp41115 = s3 ? tmp41116 : tmp41122;
  assign tmp41102 = s4 ? tmp41103 : tmp41115;
  assign tmp41133 = l1 ? tmp39379 : tmp39807;
  assign tmp41132 = s0 ? tmp41133 : 0;
  assign tmp41131 = s1 ? tmp41132 : tmp40068;
  assign tmp41135 = l1 ? tmp39429 : tmp39478;
  assign tmp41134 = s1 ? tmp41135 : tmp39479;
  assign tmp41130 = s2 ? tmp41131 : tmp41134;
  assign tmp41138 = ~(l1 ? tmp39480 : tmp39630);
  assign tmp41137 = ~(s1 ? tmp39666 : tmp41138);
  assign tmp41136 = ~(s2 ? tmp40975 : tmp41137);
  assign tmp41129 = s3 ? tmp41130 : tmp41136;
  assign tmp41141 = ~(s1 ? tmp41125 : tmp39480);
  assign tmp41140 = s2 ? tmp40980 : tmp41141;
  assign tmp41143 = ~(l1 ? tmp39480 : tmp39840);
  assign tmp41142 = s1 ? tmp40985 : tmp41143;
  assign tmp41139 = s3 ? tmp41140 : tmp41142;
  assign tmp41128 = s4 ? tmp41129 : tmp41139;
  assign tmp41101 = s5 ? tmp41102 : tmp41128;
  assign tmp41067 = s6 ? tmp41068 : tmp41101;
  assign tmp41066 = s7 ? tmp39370 : tmp41067;
  assign tmp41065 = s8 ? tmp40986 : tmp41066;
  assign tmp40893 = s9 ? tmp40894 : tmp41065;
  assign tmp41151 = l1 ? tmp40992 : tmp39567;
  assign tmp41153 = ~(l1 ? tmp40997 : tmp39567);
  assign tmp41152 = ~(s0 ? tmp41073 : tmp41153);
  assign tmp41150 = s1 ? tmp41151 : tmp41152;
  assign tmp41157 = ~(l1 ? tmp41002 : tmp39690);
  assign tmp41156 = s0 ? tmp39495 : tmp41157;
  assign tmp41158 = s0 ? tmp41073 : tmp41157;
  assign tmp41155 = s1 ? tmp41156 : tmp41158;
  assign tmp41160 = s0 ? tmp41073 : tmp40250;
  assign tmp41162 = l1 ? tmp41002 : tmp39690;
  assign tmp41163 = ~(l1 ? tmp39403 : tmp39588);
  assign tmp41161 = ~(s0 ? tmp41162 : tmp41163);
  assign tmp41159 = s1 ? tmp41160 : tmp41161;
  assign tmp41154 = ~(s2 ? tmp41155 : tmp41159);
  assign tmp41149 = s3 ? tmp41150 : tmp41154;
  assign tmp41168 = l1 ? tmp39972 : tmp39567;
  assign tmp41167 = s0 ? tmp41168 : tmp41015;
  assign tmp41170 = l1 ? tmp39403 : tmp39588;
  assign tmp41169 = ~(s0 ? tmp41170 : tmp41157);
  assign tmp41166 = s1 ? tmp41167 : tmp41169;
  assign tmp41172 = s0 ? tmp41151 : tmp40225;
  assign tmp41171 = s1 ? tmp41172 : tmp41048;
  assign tmp41165 = s2 ? tmp41166 : tmp41171;
  assign tmp41176 = l1 ? tmp39379 : tmp39690;
  assign tmp41175 = s0 ? tmp41162 : tmp41176;
  assign tmp41177 = s0 ? tmp40935 : tmp41162;
  assign tmp41174 = ~(s1 ? tmp41175 : tmp41177);
  assign tmp41173 = ~(s2 ? tmp41096 : tmp41174);
  assign tmp41164 = s3 ? tmp41165 : tmp41173;
  assign tmp41148 = s4 ? tmp41149 : tmp41164;
  assign tmp41184 = l1 ? tmp40997 : tmp39567;
  assign tmp41183 = s0 ? tmp41184 : 0;
  assign tmp41182 = s1 ? tmp41183 : tmp39484;
  assign tmp41186 = l1 ? tmp40997 : tmp39637;
  assign tmp41187 = s0 ? tmp41176 : tmp39803;
  assign tmp41185 = s1 ? tmp41186 : tmp41187;
  assign tmp41181 = s2 ? tmp41182 : tmp41185;
  assign tmp41190 = ~(l1 ? tmp39379 : tmp39725);
  assign tmp41189 = s1 ? tmp41073 : tmp41190;
  assign tmp41191 = ~(s1 ? tmp40950 : tmp41163);
  assign tmp41188 = ~(s2 ? tmp41189 : tmp41191);
  assign tmp41180 = s3 ? tmp41181 : tmp41188;
  assign tmp41196 = l1 ? tmp41002 : tmp39637;
  assign tmp41195 = s0 ? tmp39635 : tmp41196;
  assign tmp41194 = s1 ? tmp41195 : tmp41120;
  assign tmp41193 = s2 ? tmp41194 : tmp39818;
  assign tmp41200 = ~(l1 ? tmp39475 : tmp39541);
  assign tmp41199 = s0 ? tmp40903 : tmp41200;
  assign tmp41198 = s1 ? tmp41199 : tmp40964;
  assign tmp41197 = ~(s2 ? tmp41198 : tmp39650);
  assign tmp41192 = s3 ? tmp41193 : tmp41197;
  assign tmp41179 = s4 ? tmp41180 : tmp41192;
  assign tmp41206 = l1 ? tmp39379 : tmp39725;
  assign tmp41205 = s0 ? tmp41206 : 0;
  assign tmp41204 = s1 ? tmp41205 : tmp40068;
  assign tmp41208 = l1 ? tmp39429 : tmp39744;
  assign tmp41207 = s1 ? tmp41208 : tmp39479;
  assign tmp41203 = s2 ? tmp41204 : tmp41207;
  assign tmp41202 = s3 ? tmp41203 : tmp40974;
  assign tmp41211 = ~(s1 ? tmp40903 : tmp39480);
  assign tmp41210 = s2 ? tmp40980 : tmp41211;
  assign tmp41209 = s3 ? tmp41210 : tmp40984;
  assign tmp41201 = s4 ? tmp41202 : tmp41209;
  assign tmp41178 = s5 ? tmp41179 : tmp41201;
  assign tmp41147 = s6 ? tmp41148 : tmp41178;
  assign tmp41146 = s7 ? tmp39370 : tmp41147;
  assign tmp41145 = s8 ? tmp41146 : tmp39370;
  assign tmp41218 = s2 ? tmp40980 : tmp40958;
  assign tmp41217 = s3 ? tmp41218 : tmp40984;
  assign tmp41216 = s4 ? tmp40966 : tmp41217;
  assign tmp41215 = s5 ? tmp40937 : tmp41216;
  assign tmp41214 = s6 ? tmp40897 : tmp41215;
  assign tmp41224 = ~(l1 ? tmp39480 : tmp39621);
  assign tmp41223 = s2 ? tmp40980 : tmp41224;
  assign tmp41222 = s3 ? tmp41223 : tmp41142;
  assign tmp41221 = s4 ? tmp41129 : tmp41222;
  assign tmp41220 = s5 ? tmp41102 : tmp41221;
  assign tmp41219 = s6 ? tmp41068 : tmp41220;
  assign tmp41213 = s7 ? tmp41214 : tmp41219;
  assign tmp41230 = s2 ? tmp41063 : tmp40958;
  assign tmp41229 = s3 ? tmp41230 : tmp40984;
  assign tmp41228 = s4 ? tmp41056 : tmp41229;
  assign tmp41227 = s5 ? tmp41029 : tmp41228;
  assign tmp41226 = s6 ? tmp40988 : tmp41227;
  assign tmp41235 = s2 ? tmp40980 : tmp39639;
  assign tmp41234 = s3 ? tmp41235 : tmp40984;
  assign tmp41233 = s4 ? tmp41202 : tmp41234;
  assign tmp41232 = s5 ? tmp41179 : tmp41233;
  assign tmp41231 = s6 ? tmp41148 : tmp41232;
  assign tmp41225 = s7 ? tmp41226 : tmp41231;
  assign tmp41212 = s8 ? tmp41213 : tmp41225;
  assign tmp41144 = s9 ? tmp41145 : tmp41212;
  assign tmp40892 = s10 ? tmp40893 : tmp41144;
  assign tmp41239 = s7 ? tmp40896 : tmp41067;
  assign tmp41240 = s7 ? tmp40987 : tmp41147;
  assign tmp41238 = s8 ? tmp41239 : tmp41240;
  assign tmp41237 = s9 ? tmp41145 : tmp41238;
  assign tmp41236 = s10 ? tmp40893 : tmp41237;
  assign tmp40891 = s11 ? tmp40892 : tmp41236;
  assign tmp41251 = l2 ? 1 : tmp40634;
  assign tmp41250 = l1 ? tmp40901 : tmp41251;
  assign tmp41253 = l1 ? tmp39480 : tmp39423;
  assign tmp41255 = l2 ? tmp39403 : tmp40634;
  assign tmp41254 = ~(l1 ? tmp40905 : tmp41255);
  assign tmp41252 = ~(s0 ? tmp41253 : tmp41254);
  assign tmp41249 = s1 ? tmp41250 : tmp41252;
  assign tmp41260 = l2 ? tmp39460 : tmp40634;
  assign tmp41259 = ~(l1 ? tmp40910 : tmp41260);
  assign tmp41258 = s0 ? tmp39946 : tmp41259;
  assign tmp41261 = s0 ? tmp41253 : tmp41259;
  assign tmp41257 = s1 ? tmp41258 : tmp41261;
  assign tmp41263 = s0 ? tmp41253 : tmp39420;
  assign tmp41265 = l1 ? tmp40910 : tmp41260;
  assign tmp41267 = ~(l2 ? tmp39378 : tmp40634);
  assign tmp41266 = ~(l1 ? tmp39480 : tmp41267);
  assign tmp41264 = ~(s0 ? tmp41265 : tmp41266);
  assign tmp41262 = s1 ? tmp41263 : tmp41264;
  assign tmp41256 = ~(s2 ? tmp41257 : tmp41262);
  assign tmp41248 = s3 ? tmp41249 : tmp41256;
  assign tmp41272 = l1 ? tmp39918 : tmp41255;
  assign tmp41271 = s0 ? tmp41272 : tmp40655;
  assign tmp41274 = l1 ? tmp39480 : tmp41267;
  assign tmp41273 = ~(s0 ? tmp41274 : tmp41259);
  assign tmp41270 = s1 ? tmp41271 : tmp41273;
  assign tmp41276 = s0 ? tmp41250 : tmp40225;
  assign tmp41275 = s1 ? tmp41276 : tmp40696;
  assign tmp41269 = s2 ? tmp41270 : tmp41275;
  assign tmp41278 = s1 ? tmp41253 : tmp39531;
  assign tmp41281 = l1 ? tmp40933 : tmp41260;
  assign tmp41280 = s0 ? tmp41265 : tmp41281;
  assign tmp41282 = s0 ? tmp40935 : tmp41265;
  assign tmp41279 = ~(s1 ? tmp41280 : tmp41282);
  assign tmp41277 = ~(s2 ? tmp41278 : tmp41279);
  assign tmp41268 = s3 ? tmp41269 : tmp41277;
  assign tmp41247 = s4 ? tmp41248 : tmp41268;
  assign tmp41289 = l1 ? tmp40905 : tmp41255;
  assign tmp41288 = s0 ? tmp41289 : tmp40096;
  assign tmp41287 = s1 ? tmp41288 : tmp40655;
  assign tmp41291 = l1 ? tmp40905 : tmp39541;
  assign tmp41292 = s0 ? tmp41281 : tmp39401;
  assign tmp41290 = s1 ? tmp41291 : tmp41292;
  assign tmp41286 = s2 ? tmp41287 : tmp41290;
  assign tmp41294 = s1 ? tmp41253 : tmp40964;
  assign tmp41297 = l1 ? tmp39480 : tmp39532;
  assign tmp41296 = ~(s0 ? tmp41274 : tmp41297);
  assign tmp41295 = ~(s1 ? tmp40950 : tmp41296);
  assign tmp41293 = ~(s2 ? tmp41294 : tmp41295);
  assign tmp41285 = s3 ? tmp41286 : tmp41293;
  assign tmp41302 = l1 ? tmp40910 : tmp39541;
  assign tmp41301 = s0 ? tmp39635 : tmp41302;
  assign tmp41303 = s0 ? tmp40696 : tmp39639;
  assign tmp41300 = s1 ? tmp41301 : tmp41303;
  assign tmp41304 = ~(l1 ? tmp39480 : tmp39423);
  assign tmp41299 = s2 ? tmp41300 : tmp41304;
  assign tmp41307 = s0 ? tmp41253 : tmp40963;
  assign tmp41306 = s1 ? tmp41307 : tmp40964;
  assign tmp41305 = ~(s2 ? tmp41306 : tmp39650);
  assign tmp41298 = s3 ? tmp41299 : tmp41305;
  assign tmp41284 = s4 ? tmp41285 : tmp41298;
  assign tmp41313 = l1 ? tmp39379 : tmp39649;
  assign tmp41312 = s0 ? tmp41313 : 0;
  assign tmp41311 = s1 ? tmp41312 : tmp40068;
  assign tmp41315 = l1 ? tmp39429 : tmp39480;
  assign tmp41314 = s1 ? tmp41315 : tmp39479;
  assign tmp41310 = s2 ? tmp41311 : tmp41314;
  assign tmp41309 = s3 ? tmp41310 : tmp40974;
  assign tmp41318 = ~(s1 ? tmp41253 : tmp39480);
  assign tmp41317 = s2 ? tmp40980 : tmp41318;
  assign tmp41316 = s3 ? tmp41317 : tmp40984;
  assign tmp41308 = s4 ? tmp41309 : tmp41316;
  assign tmp41283 = s5 ? tmp41284 : tmp41308;
  assign tmp41246 = s6 ? tmp41247 : tmp41283;
  assign tmp41245 = s7 ? tmp39370 : tmp41246;
  assign tmp41324 = l1 ? tmp40992 : tmp41255;
  assign tmp41327 = ~(l2 ? tmp39460 : 0);
  assign tmp41326 = l1 ? tmp39403 : tmp41327;
  assign tmp41328 = ~(l1 ? tmp40997 : tmp41255);
  assign tmp41325 = ~(s0 ? tmp41326 : tmp41328);
  assign tmp41323 = s1 ? tmp41324 : tmp41325;
  assign tmp41332 = ~(l1 ? tmp41002 : tmp41260);
  assign tmp41331 = s0 ? tmp40037 : tmp41332;
  assign tmp41333 = s0 ? tmp41326 : tmp41332;
  assign tmp41330 = s1 ? tmp41331 : tmp41333;
  assign tmp41336 = ~(l1 ? tmp39385 : tmp39785);
  assign tmp41335 = s0 ? tmp41326 : tmp41336;
  assign tmp41338 = l1 ? tmp41002 : tmp41260;
  assign tmp41340 = ~(l2 ? tmp39460 : tmp40634);
  assign tmp41339 = ~(l1 ? tmp39403 : tmp41340);
  assign tmp41337 = ~(s0 ? tmp41338 : tmp41339);
  assign tmp41334 = s1 ? tmp41335 : tmp41337;
  assign tmp41329 = ~(s2 ? tmp41330 : tmp41334);
  assign tmp41322 = s3 ? tmp41323 : tmp41329;
  assign tmp41345 = l1 ? tmp39972 : tmp41255;
  assign tmp41344 = s0 ? tmp41345 : tmp40749;
  assign tmp41347 = l1 ? tmp39403 : tmp41340;
  assign tmp41346 = ~(s0 ? tmp41347 : tmp41332);
  assign tmp41343 = s1 ? tmp41344 : tmp41346;
  assign tmp41349 = s0 ? tmp41324 : tmp40225;
  assign tmp41350 = l1 ? tmp39385 : tmp39402;
  assign tmp41348 = s1 ? tmp41349 : tmp41350;
  assign tmp41342 = s2 ? tmp41343 : tmp41348;
  assign tmp41352 = s1 ? tmp41326 : tmp39531;
  assign tmp41355 = l1 ? tmp39379 : tmp41260;
  assign tmp41354 = s0 ? tmp41338 : tmp41355;
  assign tmp41356 = s0 ? tmp41027 : tmp41338;
  assign tmp41353 = ~(s1 ? tmp41354 : tmp41356);
  assign tmp41351 = ~(s2 ? tmp41352 : tmp41353);
  assign tmp41341 = s3 ? tmp41342 : tmp41351;
  assign tmp41321 = s4 ? tmp41322 : tmp41341;
  assign tmp41363 = l1 ? tmp40997 : tmp41255;
  assign tmp41362 = s0 ? tmp41363 : tmp40096;
  assign tmp41361 = s1 ? tmp41362 : tmp40749;
  assign tmp41365 = l1 ? tmp40997 : tmp41054;
  assign tmp41366 = s0 ? tmp41355 : tmp40024;
  assign tmp41364 = s1 ? tmp41365 : tmp41366;
  assign tmp41360 = s2 ? tmp41361 : tmp41364;
  assign tmp41370 = l2 ? tmp39460 : tmp39376;
  assign tmp41369 = ~(l1 ? tmp39379 : tmp41370);
  assign tmp41368 = s1 ? tmp41326 : tmp41369;
  assign tmp41372 = ~(s0 ? tmp41347 : tmp41017);
  assign tmp41371 = ~(s1 ? tmp41041 : tmp41372);
  assign tmp41367 = ~(s2 ? tmp41368 : tmp41371);
  assign tmp41359 = s3 ? tmp41360 : tmp41367;
  assign tmp41377 = l1 ? tmp41002 : tmp41054;
  assign tmp41376 = s0 ? tmp39635 : tmp41377;
  assign tmp41378 = s0 ? tmp39483 : tmp41049;
  assign tmp41375 = s1 ? tmp41376 : tmp41378;
  assign tmp41379 = ~(l1 ? tmp39403 : tmp41327);
  assign tmp41374 = s2 ? tmp41375 : tmp41379;
  assign tmp41383 = l1 ? tmp39480 : tmp41327;
  assign tmp41382 = s0 ? tmp41383 : tmp41053;
  assign tmp41381 = s1 ? tmp41382 : tmp40964;
  assign tmp41380 = ~(s2 ? tmp41381 : tmp39650);
  assign tmp41373 = s3 ? tmp41374 : tmp41380;
  assign tmp41358 = s4 ? tmp41359 : tmp41373;
  assign tmp41389 = l1 ? tmp39379 : tmp41370;
  assign tmp41388 = s0 ? tmp41389 : 0;
  assign tmp41387 = s1 ? tmp41388 : tmp41059;
  assign tmp41391 = l1 ? tmp39429 : tmp39403;
  assign tmp41390 = s1 ? tmp41391 : tmp39479;
  assign tmp41386 = s2 ? tmp41387 : tmp41390;
  assign tmp41385 = s3 ? tmp41386 : tmp40974;
  assign tmp41394 = ~(s1 ? tmp41383 : tmp39480);
  assign tmp41393 = s2 ? tmp41063 : tmp41394;
  assign tmp41392 = s3 ? tmp41393 : tmp40984;
  assign tmp41384 = s4 ? tmp41385 : tmp41392;
  assign tmp41357 = s5 ? tmp41358 : tmp41384;
  assign tmp41320 = s6 ? tmp41321 : tmp41357;
  assign tmp41319 = s7 ? tmp39370 : tmp41320;
  assign tmp41244 = s8 ? tmp41245 : tmp41319;
  assign tmp41401 = l1 ? tmp40992 : tmp39409;
  assign tmp41403 = l1 ? tmp39403 : tmp39423;
  assign tmp41404 = ~(l1 ? tmp40997 : tmp39409);
  assign tmp41402 = ~(s0 ? tmp41403 : tmp41404);
  assign tmp41400 = s1 ? tmp41401 : tmp41402;
  assign tmp41408 = l1 ? tmp39403 : tmp39518;
  assign tmp41410 = l2 ? tmp39378 : tmp39380;
  assign tmp41409 = ~(l1 ? tmp41002 : tmp41410);
  assign tmp41407 = s0 ? tmp41408 : tmp41409;
  assign tmp41412 = l1 ? tmp39403 : tmp39388;
  assign tmp41411 = s0 ? tmp41412 : tmp41409;
  assign tmp41406 = s1 ? tmp41407 : tmp41411;
  assign tmp41414 = s0 ? tmp41412 : tmp39420;
  assign tmp41416 = l1 ? tmp41002 : tmp41410;
  assign tmp41417 = ~(l1 ? tmp39403 : tmp39377);
  assign tmp41415 = ~(s0 ? tmp41416 : tmp41417);
  assign tmp41413 = s1 ? tmp41414 : tmp41415;
  assign tmp41405 = ~(s2 ? tmp41406 : tmp41413);
  assign tmp41399 = s3 ? tmp41400 : tmp41405;
  assign tmp41422 = l1 ? tmp39972 : tmp39409;
  assign tmp41421 = s0 ? tmp41422 : tmp40749;
  assign tmp41424 = l1 ? tmp39403 : tmp39377;
  assign tmp41423 = ~(s0 ? tmp41424 : tmp41409);
  assign tmp41420 = s1 ? tmp41421 : tmp41423;
  assign tmp41426 = s0 ? tmp41401 : tmp40225;
  assign tmp41425 = s1 ? tmp41426 : tmp39483;
  assign tmp41419 = s2 ? tmp41420 : tmp41425;
  assign tmp41428 = s1 ? tmp41403 : tmp39531;
  assign tmp41431 = l1 ? tmp39379 : tmp41410;
  assign tmp41430 = s0 ? tmp41416 : tmp41431;
  assign tmp41432 = s0 ? tmp40935 : tmp41416;
  assign tmp41429 = ~(s1 ? tmp41430 : tmp41432);
  assign tmp41427 = ~(s2 ? tmp41428 : tmp41429);
  assign tmp41418 = s3 ? tmp41419 : tmp41427;
  assign tmp41398 = s4 ? tmp41399 : tmp41418;
  assign tmp41439 = l1 ? tmp40997 : tmp39409;
  assign tmp41438 = s0 ? tmp41439 : tmp40096;
  assign tmp41440 = ~(l1 ? tmp39403 : tmp39518);
  assign tmp41437 = s1 ? tmp41438 : tmp41440;
  assign tmp41442 = l1 ? tmp40997 : tmp39435;
  assign tmp41443 = s0 ? tmp41431 : tmp39401;
  assign tmp41441 = s1 ? tmp41442 : tmp41443;
  assign tmp41436 = s2 ? tmp41437 : tmp41441;
  assign tmp41445 = s1 ? tmp41412 : tmp41127;
  assign tmp41447 = ~(s0 ? tmp41424 : tmp41092);
  assign tmp41446 = ~(s1 ? tmp40950 : tmp41447);
  assign tmp41444 = ~(s2 ? tmp41445 : tmp41446);
  assign tmp41435 = s3 ? tmp41436 : tmp41444;
  assign tmp41452 = l1 ? tmp41002 : tmp39435;
  assign tmp41451 = s0 ? tmp39635 : tmp41452;
  assign tmp41453 = s0 ? tmp39483 : tmp39818;
  assign tmp41450 = s1 ? tmp41451 : tmp41453;
  assign tmp41454 = ~(l1 ? tmp39403 : tmp39388);
  assign tmp41449 = s2 ? tmp41450 : tmp41454;
  assign tmp41458 = l1 ? tmp39480 : tmp39388;
  assign tmp41457 = s0 ? tmp41458 : tmp41126;
  assign tmp41456 = s1 ? tmp41457 : tmp41127;
  assign tmp41455 = ~(s2 ? tmp41456 : tmp39650);
  assign tmp41448 = s3 ? tmp41449 : tmp41455;
  assign tmp41434 = s4 ? tmp41435 : tmp41448;
  assign tmp41463 = s0 ? tmp40935 : 0;
  assign tmp41462 = s1 ? tmp41463 : tmp40068;
  assign tmp41464 = s1 ? tmp39549 : tmp39479;
  assign tmp41461 = s2 ? tmp41462 : tmp41464;
  assign tmp41460 = s3 ? tmp41461 : tmp41136;
  assign tmp41467 = ~(s1 ? tmp41458 : tmp39480);
  assign tmp41466 = s2 ? tmp40980 : tmp41467;
  assign tmp41465 = s3 ? tmp41466 : tmp41142;
  assign tmp41459 = s4 ? tmp41460 : tmp41465;
  assign tmp41433 = s5 ? tmp41434 : tmp41459;
  assign tmp41397 = s6 ? tmp41398 : tmp41433;
  assign tmp41396 = s7 ? tmp39370 : tmp41397;
  assign tmp41395 = s8 ? tmp41319 : tmp41396;
  assign tmp41243 = s9 ? tmp41244 : tmp41395;
  assign tmp41475 = l1 ? tmp40992 : tmp41251;
  assign tmp41477 = ~(l1 ? tmp40997 : tmp41251);
  assign tmp41476 = ~(s0 ? tmp41403 : tmp41477);
  assign tmp41474 = s1 ? tmp41475 : tmp41476;
  assign tmp41482 = l2 ? tmp39378 : tmp40634;
  assign tmp41481 = ~(l1 ? tmp41002 : tmp41482);
  assign tmp41480 = s0 ? tmp40731 : tmp41481;
  assign tmp41483 = s0 ? tmp41403 : tmp41481;
  assign tmp41479 = s1 ? tmp41480 : tmp41483;
  assign tmp41485 = s0 ? tmp41403 : tmp39420;
  assign tmp41487 = l1 ? tmp41002 : tmp41482;
  assign tmp41488 = ~(l1 ? tmp39403 : tmp41267);
  assign tmp41486 = ~(s0 ? tmp41487 : tmp41488);
  assign tmp41484 = s1 ? tmp41485 : tmp41486;
  assign tmp41478 = ~(s2 ? tmp41479 : tmp41484);
  assign tmp41473 = s3 ? tmp41474 : tmp41478;
  assign tmp41493 = l1 ? tmp39972 : tmp41251;
  assign tmp41492 = s0 ? tmp41493 : tmp40749;
  assign tmp41495 = l1 ? tmp39403 : tmp41267;
  assign tmp41494 = ~(s0 ? tmp41495 : tmp41481);
  assign tmp41491 = s1 ? tmp41492 : tmp41494;
  assign tmp41497 = s0 ? tmp41475 : tmp40225;
  assign tmp41496 = s1 ? tmp41497 : tmp39483;
  assign tmp41490 = s2 ? tmp41491 : tmp41496;
  assign tmp41501 = l1 ? tmp39379 : tmp41482;
  assign tmp41500 = s0 ? tmp41487 : tmp41501;
  assign tmp41502 = s0 ? tmp40935 : tmp41487;
  assign tmp41499 = ~(s1 ? tmp41500 : tmp41502);
  assign tmp41498 = ~(s2 ? tmp41428 : tmp41499);
  assign tmp41489 = s3 ? tmp41490 : tmp41498;
  assign tmp41472 = s4 ? tmp41473 : tmp41489;
  assign tmp41509 = l1 ? tmp40997 : tmp41251;
  assign tmp41508 = s0 ? tmp41509 : tmp40096;
  assign tmp41510 = ~(l1 ? tmp39403 : tmp39404);
  assign tmp41507 = s1 ? tmp41508 : tmp41510;
  assign tmp41512 = l1 ? tmp40997 : tmp39541;
  assign tmp41513 = s0 ? tmp41501 : tmp39401;
  assign tmp41511 = s1 ? tmp41512 : tmp41513;
  assign tmp41506 = s2 ? tmp41507 : tmp41511;
  assign tmp41515 = s1 ? tmp41403 : tmp40964;
  assign tmp41517 = ~(s0 ? tmp41495 : tmp41170);
  assign tmp41516 = ~(s1 ? tmp40950 : tmp41517);
  assign tmp41514 = ~(s2 ? tmp41515 : tmp41516);
  assign tmp41505 = s3 ? tmp41506 : tmp41514;
  assign tmp41522 = l1 ? tmp41002 : tmp39541;
  assign tmp41521 = s0 ? tmp39635 : tmp41522;
  assign tmp41520 = s1 ? tmp41521 : tmp41453;
  assign tmp41523 = ~(l1 ? tmp39403 : tmp39423);
  assign tmp41519 = s2 ? tmp41520 : tmp41523;
  assign tmp41526 = s0 ? tmp41253 : tmp41200;
  assign tmp41525 = s1 ? tmp41526 : tmp40964;
  assign tmp41524 = ~(s2 ? tmp41525 : tmp39650);
  assign tmp41518 = s3 ? tmp41519 : tmp41524;
  assign tmp41504 = s4 ? tmp41505 : tmp41518;
  assign tmp41503 = s5 ? tmp41504 : tmp41308;
  assign tmp41471 = s6 ? tmp41472 : tmp41503;
  assign tmp41470 = s7 ? tmp39370 : tmp41471;
  assign tmp41469 = s8 ? tmp41470 : tmp39370;
  assign tmp41533 = s2 ? tmp40980 : tmp41304;
  assign tmp41532 = s3 ? tmp41533 : tmp40984;
  assign tmp41531 = s4 ? tmp41309 : tmp41532;
  assign tmp41530 = s5 ? tmp41284 : tmp41531;
  assign tmp41529 = s6 ? tmp41247 : tmp41530;
  assign tmp41539 = ~(l1 ? tmp39480 : tmp39388);
  assign tmp41538 = s2 ? tmp40980 : tmp41539;
  assign tmp41537 = s3 ? tmp41538 : tmp41142;
  assign tmp41536 = s4 ? tmp41460 : tmp41537;
  assign tmp41535 = s5 ? tmp41434 : tmp41536;
  assign tmp41534 = s6 ? tmp41398 : tmp41535;
  assign tmp41528 = s7 ? tmp41529 : tmp41534;
  assign tmp41546 = ~(l1 ? tmp39480 : tmp41327);
  assign tmp41545 = s2 ? tmp41063 : tmp41546;
  assign tmp41544 = s3 ? tmp41545 : tmp40984;
  assign tmp41543 = s4 ? tmp41385 : tmp41544;
  assign tmp41542 = s5 ? tmp41358 : tmp41543;
  assign tmp41541 = s6 ? tmp41321 : tmp41542;
  assign tmp41548 = s5 ? tmp41504 : tmp41531;
  assign tmp41547 = s6 ? tmp41472 : tmp41548;
  assign tmp41540 = s7 ? tmp41541 : tmp41547;
  assign tmp41527 = s8 ? tmp41528 : tmp41540;
  assign tmp41468 = s9 ? tmp41469 : tmp41527;
  assign tmp41242 = s10 ? tmp41243 : tmp41468;
  assign tmp41552 = s7 ? tmp41246 : tmp41397;
  assign tmp41553 = s7 ? tmp41320 : tmp41471;
  assign tmp41551 = s8 ? tmp41552 : tmp41553;
  assign tmp41550 = s9 ? tmp41469 : tmp41551;
  assign tmp41549 = s10 ? tmp41243 : tmp41550;
  assign tmp41241 = s11 ? tmp41242 : tmp41549;
  assign tmp40890 = s12 ? tmp40891 : tmp41241;
  assign tmp40407 = s13 ? tmp40408 : tmp40890;
  assign tmp39363 = s14 ? tmp39364 : tmp40407;
  assign tmp41564 = l1 ? tmp39384 : tmp39409;
  assign tmp41566 = ~(l1 ? tmp41251 : tmp39409);
  assign tmp41565 = ~(s0 ? tmp39422 : tmp41566);
  assign tmp41563 = s1 ? tmp41564 : tmp41565;
  assign tmp41570 = l1 ? tmp39375 : tmp39518;
  assign tmp41571 = ~(l1 ? tmp41251 : tmp41410);
  assign tmp41569 = s0 ? tmp41570 : tmp41571;
  assign tmp41573 = l1 ? tmp39588 : tmp39388;
  assign tmp41572 = s0 ? tmp41573 : tmp41571;
  assign tmp41568 = s1 ? tmp41569 : tmp41572;
  assign tmp41575 = s0 ? tmp41573 : tmp39420;
  assign tmp41577 = l1 ? tmp41251 : tmp41410;
  assign tmp41578 = ~(l1 ? tmp39439 : tmp39377);
  assign tmp41576 = ~(s0 ? tmp41577 : tmp41578);
  assign tmp41574 = s1 ? tmp41575 : tmp41576;
  assign tmp41567 = ~(s2 ? tmp41568 : tmp41574);
  assign tmp41562 = s3 ? tmp41563 : tmp41567;
  assign tmp41582 = s0 ? tmp41564 : tmp40024;
  assign tmp41584 = l1 ? tmp39439 : tmp39377;
  assign tmp41583 = ~(s0 ? tmp41584 : tmp41571);
  assign tmp41581 = s1 ? tmp41582 : tmp41583;
  assign tmp41586 = s0 ? tmp41564 : tmp40225;
  assign tmp41587 = l1 ? tmp39384 : 1;
  assign tmp41585 = s1 ? tmp41586 : tmp41587;
  assign tmp41580 = s2 ? tmp41581 : tmp41585;
  assign tmp41590 = l1 ? tmp39378 : tmp39532;
  assign tmp41589 = s1 ? tmp39422 : tmp41590;
  assign tmp41593 = l1 ? tmp39541 : tmp41410;
  assign tmp41592 = s0 ? tmp41577 : tmp41593;
  assign tmp41595 = l1 ? tmp39435 : tmp39604;
  assign tmp41594 = s0 ? tmp41595 : tmp41577;
  assign tmp41591 = ~(s1 ? tmp41592 : tmp41594);
  assign tmp41588 = ~(s2 ? tmp41589 : tmp41591);
  assign tmp41579 = s3 ? tmp41580 : tmp41588;
  assign tmp41561 = s4 ? tmp41562 : tmp41579;
  assign tmp41602 = l1 ? tmp41251 : tmp39409;
  assign tmp41601 = s0 ? tmp41602 : tmp40096;
  assign tmp41603 = ~(l1 ? tmp39375 : tmp39518);
  assign tmp41600 = s1 ? tmp41601 : tmp41603;
  assign tmp41605 = l1 ? tmp41251 : tmp39435;
  assign tmp41606 = s0 ? tmp41593 : tmp39401;
  assign tmp41604 = s1 ? tmp41605 : tmp41606;
  assign tmp41599 = s2 ? tmp41600 : tmp41604;
  assign tmp41609 = ~(l1 ? tmp39541 : tmp39604);
  assign tmp41608 = s1 ? tmp41573 : tmp41609;
  assign tmp41612 = l1 ? tmp39435 : tmp39501;
  assign tmp41611 = s0 ? tmp41595 : tmp41612;
  assign tmp41614 = l1 ? tmp39439 : tmp39493;
  assign tmp41613 = ~(s0 ? tmp41584 : tmp41614);
  assign tmp41610 = ~(s1 ? tmp41611 : tmp41613);
  assign tmp41607 = ~(s2 ? tmp41608 : tmp41610);
  assign tmp41598 = s3 ? tmp41599 : tmp41607;
  assign tmp41619 = l1 ? 1 : tmp39604;
  assign tmp41618 = s0 ? tmp41619 : tmp41605;
  assign tmp41620 = s0 ? tmp41587 : tmp39980;
  assign tmp41617 = s1 ? tmp41618 : tmp41620;
  assign tmp41616 = s2 ? tmp41617 : tmp39387;
  assign tmp41623 = s0 ? tmp40269 : tmp39535;
  assign tmp41622 = s1 ? tmp41623 : tmp41609;
  assign tmp41625 = l1 ? tmp39501 : tmp39513;
  assign tmp41624 = s1 ? tmp41625 : tmp41590;
  assign tmp41621 = ~(s2 ? tmp41622 : tmp41624);
  assign tmp41615 = s3 ? tmp41616 : tmp41621;
  assign tmp41597 = s4 ? tmp41598 : tmp41615;
  assign tmp41631 = l1 ? tmp39541 : tmp39604;
  assign tmp41630 = s0 ? tmp41631 : tmp39509;
  assign tmp41633 = l1 ? tmp39532 : tmp39375;
  assign tmp41632 = ~(s0 ? tmp39511 : tmp41633);
  assign tmp41629 = s1 ? tmp41630 : tmp41632;
  assign tmp41628 = s2 ? tmp41629 : tmp40275;
  assign tmp41636 = ~(l1 ? tmp39435 : tmp39501);
  assign tmp41635 = s1 ? tmp39651 : tmp41636;
  assign tmp41638 = l1 ? 1 : tmp39435;
  assign tmp41637 = ~(s1 ? tmp41638 : tmp39999);
  assign tmp41634 = ~(s2 ? tmp41635 : tmp41637);
  assign tmp41627 = s3 ? tmp41628 : tmp41634;
  assign tmp41641 = s1 ? tmp39435 : tmp41595;
  assign tmp41643 = l1 ? tmp39532 : tmp39388;
  assign tmp41642 = ~(s0 ? tmp39511 : tmp41643);
  assign tmp41640 = s2 ? tmp41641 : tmp41642;
  assign tmp41645 = ~(l1 ? tmp39475 : tmp39840);
  assign tmp41644 = s1 ? tmp41595 : tmp41645;
  assign tmp41639 = s3 ? tmp41640 : tmp41644;
  assign tmp41626 = s4 ? tmp41627 : tmp41639;
  assign tmp41596 = s5 ? tmp41597 : tmp41626;
  assign tmp41560 = s6 ? tmp41561 : tmp41596;
  assign tmp41559 = s7 ? tmp39370 : tmp41560;
  assign tmp41647 = s8 ? tmp41559 : tmp39370;
  assign tmp41653 = ~(l1 ? tmp39532 : tmp39388);
  assign tmp41652 = s2 ? tmp41641 : tmp41653;
  assign tmp41651 = s3 ? tmp41652 : tmp41644;
  assign tmp41650 = s4 ? tmp41627 : tmp41651;
  assign tmp41649 = s5 ? tmp41597 : tmp41650;
  assign tmp41648 = s6 ? tmp41561 : tmp41649;
  assign tmp41646 = s9 ? tmp41647 : tmp41648;
  assign tmp41558 = s10 ? tmp41559 : tmp41646;
  assign tmp41655 = s9 ? tmp41647 : tmp41560;
  assign tmp41654 = s10 ? tmp41559 : tmp41655;
  assign tmp41557 = s11 ? tmp41558 : tmp41654;
  assign tmp41663 = l1 ? tmp39397 : tmp40637;
  assign tmp41665 = ~(l1 ? tmp40423 : tmp39409);
  assign tmp41664 = ~(s0 ? tmp39422 : tmp41665);
  assign tmp41662 = s1 ? tmp41663 : tmp41664;
  assign tmp41669 = ~(l1 ? tmp40423 : tmp40642);
  assign tmp41668 = s0 ? tmp41570 : tmp41669;
  assign tmp41670 = s0 ? tmp39414 : tmp41669;
  assign tmp41667 = s1 ? tmp41668 : tmp41670;
  assign tmp41673 = l1 ? tmp40423 : tmp40642;
  assign tmp41675 = l2 ? tmp39440 : 1;
  assign tmp41674 = ~(l1 ? tmp41675 : tmp39388);
  assign tmp41672 = ~(s0 ? tmp41673 : tmp41674);
  assign tmp41671 = s1 ? tmp39446 : tmp41672;
  assign tmp41666 = ~(s2 ? tmp41667 : tmp41671);
  assign tmp41661 = s3 ? tmp41662 : tmp41666;
  assign tmp41680 = l1 ? tmp41675 : tmp39388;
  assign tmp41679 = ~(s0 ? tmp41680 : tmp41669);
  assign tmp41678 = s1 ? tmp41582 : tmp41679;
  assign tmp41682 = s0 ? tmp41663 : tmp40225;
  assign tmp41681 = s1 ? tmp41682 : tmp41587;
  assign tmp41677 = s2 ? tmp41678 : tmp41681;
  assign tmp41685 = l1 ? tmp39501 : tmp39429;
  assign tmp41684 = s1 ? tmp39422 : tmp41685;
  assign tmp41688 = l1 ? tmp39547 : tmp40642;
  assign tmp41687 = s0 ? tmp41673 : tmp41688;
  assign tmp41690 = l1 ? tmp39527 : tmp39434;
  assign tmp41689 = s0 ? tmp41690 : tmp41673;
  assign tmp41686 = ~(s1 ? tmp41687 : tmp41689);
  assign tmp41683 = ~(s2 ? tmp41684 : tmp41686);
  assign tmp41676 = s3 ? tmp41677 : tmp41683;
  assign tmp41660 = s4 ? tmp41661 : tmp41676;
  assign tmp41697 = l1 ? tmp40423 : tmp39409;
  assign tmp41696 = s0 ? tmp41697 : tmp40096;
  assign tmp41695 = s1 ? tmp41696 : tmp41603;
  assign tmp41699 = l1 ? tmp40423 : tmp39435;
  assign tmp41700 = s0 ? tmp41688 : tmp39401;
  assign tmp41698 = s1 ? tmp41699 : tmp41700;
  assign tmp41694 = s2 ? tmp41695 : tmp41698;
  assign tmp41703 = ~(l1 ? tmp39547 : tmp39434);
  assign tmp41702 = s1 ? tmp39414 : tmp41703;
  assign tmp41706 = l1 ? tmp39527 : tmp39378;
  assign tmp41705 = s0 ? tmp41690 : tmp41706;
  assign tmp41708 = l1 ? tmp41675 : tmp39621;
  assign tmp41707 = ~(s0 ? tmp41680 : tmp41708);
  assign tmp41704 = ~(s1 ? tmp41705 : tmp41707);
  assign tmp41701 = ~(s2 ? tmp41702 : tmp41704);
  assign tmp41693 = s3 ? tmp41694 : tmp41701;
  assign tmp41713 = l1 ? tmp39513 : tmp39434;
  assign tmp41714 = l1 ? tmp40423 : tmp39527;
  assign tmp41712 = s0 ? tmp41713 : tmp41714;
  assign tmp41711 = s1 ? tmp41712 : tmp41620;
  assign tmp41710 = s2 ? tmp41711 : tmp39387;
  assign tmp41718 = ~(l1 ? tmp39459 : tmp39527);
  assign tmp41717 = s0 ? tmp40269 : tmp41718;
  assign tmp41716 = s1 ? tmp41717 : tmp41703;
  assign tmp41720 = s0 ? tmp41685 : tmp39465;
  assign tmp41719 = s1 ? tmp39499 : tmp41720;
  assign tmp41715 = ~(s2 ? tmp41716 : tmp41719);
  assign tmp41709 = s3 ? tmp41710 : tmp41715;
  assign tmp41692 = s4 ? tmp41693 : tmp41709;
  assign tmp41726 = l1 ? tmp39547 : tmp39434;
  assign tmp41727 = ~(l1 ? tmp39501 : 1);
  assign tmp41725 = s0 ? tmp41726 : tmp41727;
  assign tmp41724 = s1 ? tmp41725 : tmp39658;
  assign tmp41723 = s2 ? tmp41724 : tmp40275;
  assign tmp41730 = ~(l1 ? tmp39527 : tmp39378);
  assign tmp41729 = s1 ? 1 : tmp41730;
  assign tmp41732 = l1 ? tmp39513 : tmp39527;
  assign tmp41731 = ~(s1 ? tmp41732 : tmp39999);
  assign tmp41728 = ~(s2 ? tmp41729 : tmp41731);
  assign tmp41722 = s3 ? tmp41723 : tmp41728;
  assign tmp41735 = s1 ? tmp39671 : tmp41690;
  assign tmp41734 = s2 ? tmp41735 : tmp40278;
  assign tmp41738 = l2 ? tmp39379 : 1;
  assign tmp41737 = ~(l1 ? tmp41738 : tmp39630);
  assign tmp41736 = s1 ? tmp41690 : tmp41737;
  assign tmp41733 = s3 ? tmp41734 : tmp41736;
  assign tmp41721 = s4 ? tmp41722 : tmp41733;
  assign tmp41691 = s5 ? tmp41692 : tmp41721;
  assign tmp41659 = s6 ? tmp41660 : tmp41691;
  assign tmp41658 = s7 ? tmp39370 : tmp41659;
  assign tmp41740 = s8 ? tmp41658 : tmp39370;
  assign tmp41746 = s1 ? tmp39499 : tmp41685;
  assign tmp41745 = ~(s2 ? tmp41716 : tmp41746);
  assign tmp41744 = s3 ? tmp41710 : tmp41745;
  assign tmp41743 = s4 ? tmp41693 : tmp41744;
  assign tmp41742 = s5 ? tmp41743 : tmp41721;
  assign tmp41741 = s6 ? tmp41660 : tmp41742;
  assign tmp41739 = s9 ? tmp41740 : tmp41741;
  assign tmp41657 = s10 ? tmp41658 : tmp41739;
  assign tmp41748 = s9 ? tmp41740 : tmp41659;
  assign tmp41747 = s10 ? tmp41658 : tmp41748;
  assign tmp41656 = s11 ? tmp41657 : tmp41747;
  assign tmp41556 = s12 ? tmp41557 : tmp41656;
  assign tmp41759 = l1 ? tmp39384 : tmp40100;
  assign tmp41761 = ~(l1 ? tmp41251 : tmp39918);
  assign tmp41760 = ~(s0 ? tmp39477 : tmp41761);
  assign tmp41758 = s1 ? tmp41759 : tmp41760;
  assign tmp41765 = l1 ? tmp39375 : tmp39744;
  assign tmp41766 = ~(l1 ? tmp41251 : tmp40901);
  assign tmp41764 = s0 ? tmp41765 : tmp41766;
  assign tmp41768 = l1 ? tmp39588 : tmp39744;
  assign tmp41767 = s0 ? tmp41768 : tmp41766;
  assign tmp41763 = s1 ? tmp41764 : tmp41767;
  assign tmp41770 = s0 ? tmp41768 : tmp39420;
  assign tmp41772 = l1 ? tmp41251 : tmp40901;
  assign tmp41773 = ~(l1 ? tmp39439 : tmp39637);
  assign tmp41771 = ~(s0 ? tmp41772 : tmp41773);
  assign tmp41769 = s1 ? tmp41770 : tmp41771;
  assign tmp41762 = ~(s2 ? tmp41763 : tmp41769);
  assign tmp41757 = s3 ? tmp41758 : tmp41762;
  assign tmp41778 = l1 ? tmp39384 : tmp39918;
  assign tmp41777 = s0 ? tmp41778 : tmp40024;
  assign tmp41780 = l1 ? tmp39439 : tmp39637;
  assign tmp41779 = ~(s0 ? tmp41780 : tmp41766);
  assign tmp41776 = s1 ? tmp41777 : tmp41779;
  assign tmp41782 = s0 ? tmp41759 : tmp40225;
  assign tmp41781 = s1 ? tmp41782 : tmp39569;
  assign tmp41775 = s2 ? tmp41776 : tmp41781;
  assign tmp41784 = s1 ? tmp39477 : tmp39666;
  assign tmp41787 = l1 ? tmp39541 : tmp40901;
  assign tmp41786 = s0 ? tmp41772 : tmp41787;
  assign tmp41789 = l1 ? tmp39435 : tmp39439;
  assign tmp41788 = s0 ? tmp41789 : tmp41772;
  assign tmp41785 = ~(s1 ? tmp41786 : tmp41788);
  assign tmp41783 = ~(s2 ? tmp41784 : tmp41785);
  assign tmp41774 = s3 ? tmp41775 : tmp41783;
  assign tmp41756 = s4 ? tmp41757 : tmp41774;
  assign tmp41796 = l1 ? tmp41251 : tmp39918;
  assign tmp41795 = s0 ? tmp41796 : tmp40096;
  assign tmp41794 = s1 ? tmp41795 : tmp41603;
  assign tmp41798 = l1 ? tmp41251 : tmp39375;
  assign tmp41799 = s0 ? tmp41787 : tmp39401;
  assign tmp41797 = s1 ? tmp41798 : tmp41799;
  assign tmp41793 = s2 ? tmp41794 : tmp41797;
  assign tmp41802 = ~(l1 ? tmp39541 : tmp39439);
  assign tmp41801 = s1 ? tmp41768 : tmp41802;
  assign tmp41805 = l1 ? tmp39435 : tmp39378;
  assign tmp41804 = s0 ? tmp41789 : tmp41805;
  assign tmp41807 = l1 ? tmp39439 : tmp39541;
  assign tmp41806 = ~(s0 ? tmp41780 : tmp41807);
  assign tmp41803 = ~(s1 ? tmp41804 : tmp41806);
  assign tmp41800 = ~(s2 ? tmp41801 : tmp41803);
  assign tmp41792 = s3 ? tmp41793 : tmp41800;
  assign tmp41812 = l1 ? tmp41251 : tmp39588;
  assign tmp41811 = s0 ? tmp39474 : tmp41812;
  assign tmp41813 = s0 ? tmp41587 : tmp40225;
  assign tmp41810 = s1 ? tmp41811 : tmp41813;
  assign tmp41814 = ~(l1 ? tmp39375 : tmp39637);
  assign tmp41809 = s2 ? tmp41810 : tmp41814;
  assign tmp41818 = l1 ? tmp39429 : tmp39637;
  assign tmp41817 = s0 ? tmp41818 : tmp40917;
  assign tmp41819 = ~(l1 ? tmp39541 : tmp39475);
  assign tmp41816 = s1 ? tmp41817 : tmp41819;
  assign tmp41820 = s1 ? tmp39500 : tmp39666;
  assign tmp41815 = ~(s2 ? tmp41816 : tmp41820);
  assign tmp41808 = s3 ? tmp41809 : tmp41815;
  assign tmp41791 = s4 ? tmp41792 : tmp41808;
  assign tmp41826 = l1 ? tmp39541 : tmp39439;
  assign tmp41825 = s0 ? tmp41826 : tmp39509;
  assign tmp41824 = s1 ? tmp41825 : tmp39561;
  assign tmp41823 = s2 ? tmp41824 : tmp40275;
  assign tmp41829 = ~(l1 ? tmp39435 : tmp39378);
  assign tmp41828 = s1 ? tmp41638 : tmp41829;
  assign tmp41832 = ~(l1 ? tmp39429 : tmp39541);
  assign tmp41831 = s0 ? tmp39534 : tmp41832;
  assign tmp41830 = ~(s1 ? tmp39531 : tmp41831);
  assign tmp41827 = ~(s2 ? tmp41828 : tmp41830);
  assign tmp41822 = s3 ? tmp41823 : tmp41827;
  assign tmp41836 = l1 ? tmp39435 : 1;
  assign tmp41835 = s1 ? tmp41836 : tmp41789;
  assign tmp41837 = ~(l1 ? tmp39532 : tmp39637);
  assign tmp41834 = s2 ? tmp41835 : tmp41837;
  assign tmp41839 = s1 ? tmp41805 : tmp41200;
  assign tmp41838 = s2 ? tmp41839 : tmp39534;
  assign tmp41833 = s3 ? tmp41834 : tmp41838;
  assign tmp41821 = s4 ? tmp41822 : tmp41833;
  assign tmp41790 = s5 ? tmp41791 : tmp41821;
  assign tmp41755 = s6 ? tmp41756 : tmp41790;
  assign tmp41754 = s7 ? tmp39370 : tmp41755;
  assign tmp41845 = l1 ? tmp39384 : tmp40564;
  assign tmp41847 = l1 ? tmp39402 : tmp39404;
  assign tmp41848 = ~(l1 ? tmp41251 : tmp39972);
  assign tmp41846 = ~(s0 ? tmp41847 : tmp41848);
  assign tmp41844 = s1 ? tmp41845 : tmp41846;
  assign tmp41852 = ~(l1 ? tmp41251 : tmp40992);
  assign tmp41851 = s0 ? tmp41570 : tmp41852;
  assign tmp41854 = l1 ? tmp39588 : tmp39518;
  assign tmp41853 = s0 ? tmp41854 : tmp41852;
  assign tmp41850 = s1 ? tmp41851 : tmp41853;
  assign tmp41856 = s0 ? tmp41854 : tmp39420;
  assign tmp41858 = l1 ? tmp41251 : tmp40992;
  assign tmp41859 = ~(l1 ? tmp39439 : tmp39615);
  assign tmp41857 = ~(s0 ? tmp41858 : tmp41859);
  assign tmp41855 = s1 ? tmp41856 : tmp41857;
  assign tmp41849 = ~(s2 ? tmp41850 : tmp41855);
  assign tmp41843 = s3 ? tmp41844 : tmp41849;
  assign tmp41864 = l1 ? tmp39384 : tmp39972;
  assign tmp41863 = s0 ? tmp41864 : tmp40024;
  assign tmp41866 = l1 ? tmp39439 : tmp39615;
  assign tmp41865 = ~(s0 ? tmp41866 : tmp41852);
  assign tmp41862 = s1 ? tmp41863 : tmp41865;
  assign tmp41868 = s0 ? tmp41845 : tmp40225;
  assign tmp41869 = l1 ? tmp39384 : tmp39429;
  assign tmp41867 = s1 ? tmp41868 : tmp41869;
  assign tmp41861 = s2 ? tmp41862 : tmp41867;
  assign tmp41871 = s1 ? tmp41847 : tmp39666;
  assign tmp41874 = l1 ? tmp39541 : tmp40992;
  assign tmp41873 = s0 ? tmp41858 : tmp41874;
  assign tmp41876 = l1 ? tmp39435 : tmp39475;
  assign tmp41875 = s0 ? tmp41876 : tmp41858;
  assign tmp41872 = ~(s1 ? tmp41873 : tmp41875);
  assign tmp41870 = ~(s2 ? tmp41871 : tmp41872);
  assign tmp41860 = s3 ? tmp41861 : tmp41870;
  assign tmp41842 = s4 ? tmp41843 : tmp41860;
  assign tmp41883 = l1 ? tmp41251 : tmp39972;
  assign tmp41882 = s0 ? tmp41883 : tmp40096;
  assign tmp41881 = s1 ? tmp41882 : tmp41603;
  assign tmp41885 = l1 ? tmp41251 : tmp39429;
  assign tmp41886 = s0 ? tmp41874 : tmp39401;
  assign tmp41884 = s1 ? tmp41885 : tmp41886;
  assign tmp41880 = s2 ? tmp41881 : tmp41884;
  assign tmp41888 = s1 ? tmp41854 : tmp41819;
  assign tmp41890 = s0 ? tmp41876 : tmp41805;
  assign tmp41892 = l1 ? tmp39439 : tmp41054;
  assign tmp41891 = ~(s0 ? tmp41866 : tmp41892);
  assign tmp41889 = ~(s1 ? tmp41890 : tmp41891);
  assign tmp41887 = ~(s2 ? tmp41888 : tmp41889);
  assign tmp41879 = s3 ? tmp41880 : tmp41887;
  assign tmp41897 = l1 ? tmp41251 : tmp39532;
  assign tmp41896 = s0 ? tmp39474 : tmp41897;
  assign tmp41898 = s0 ? tmp41587 : tmp39803;
  assign tmp41895 = s1 ? tmp41896 : tmp41898;
  assign tmp41899 = ~(l1 ? tmp39375 : tmp39615);
  assign tmp41894 = s2 ? tmp41895 : tmp41899;
  assign tmp41903 = l1 ? tmp39429 : tmp39615;
  assign tmp41902 = s0 ? tmp41903 : tmp40951;
  assign tmp41901 = s1 ? tmp41902 : tmp41819;
  assign tmp41900 = ~(s2 ? tmp41901 : tmp41820);
  assign tmp41893 = s3 ? tmp41894 : tmp41900;
  assign tmp41878 = s4 ? tmp41879 : tmp41893;
  assign tmp41909 = l1 ? tmp39541 : tmp39475;
  assign tmp41908 = s0 ? tmp41909 : tmp39509;
  assign tmp41910 = ~(l1 ? tmp39532 : tmp39402);
  assign tmp41907 = s1 ? tmp41908 : tmp41910;
  assign tmp41906 = s2 ? tmp41907 : tmp40275;
  assign tmp41905 = s3 ? tmp41906 : tmp41827;
  assign tmp41913 = s1 ? tmp41836 : tmp41876;
  assign tmp41914 = ~(l1 ? tmp39532 : tmp39615);
  assign tmp41912 = s2 ? tmp41913 : tmp41914;
  assign tmp41911 = s3 ? tmp41912 : tmp41838;
  assign tmp41904 = s4 ? tmp41905 : tmp41911;
  assign tmp41877 = s5 ? tmp41878 : tmp41904;
  assign tmp41841 = s6 ? tmp41842 : tmp41877;
  assign tmp41840 = s7 ? tmp39370 : tmp41841;
  assign tmp41753 = s8 ? tmp41754 : tmp41840;
  assign tmp41921 = l1 ? tmp39384 : tmp40489;
  assign tmp41923 = ~(l1 ? tmp41251 : tmp39587);
  assign tmp41922 = ~(s0 ? tmp41847 : tmp41923);
  assign tmp41920 = s1 ? tmp41921 : tmp41922;
  assign tmp41928 = l2 ? tmp39379 : tmp39398;
  assign tmp41927 = ~(l1 ? tmp41251 : tmp41928);
  assign tmp41926 = s0 ? tmp41570 : tmp41927;
  assign tmp41929 = s0 ? tmp41854 : tmp41927;
  assign tmp41925 = s1 ? tmp41926 : tmp41929;
  assign tmp41932 = l1 ? tmp41251 : tmp41928;
  assign tmp41933 = ~(l1 ? tmp39439 : tmp40477);
  assign tmp41931 = ~(s0 ? tmp41932 : tmp41933);
  assign tmp41930 = s1 ? tmp41856 : tmp41931;
  assign tmp41924 = ~(s2 ? tmp41925 : tmp41930);
  assign tmp41919 = s3 ? tmp41920 : tmp41924;
  assign tmp41938 = l1 ? tmp39384 : tmp39587;
  assign tmp41937 = s0 ? tmp41938 : tmp40024;
  assign tmp41940 = l1 ? tmp39439 : tmp40477;
  assign tmp41939 = ~(s0 ? tmp41940 : tmp41927);
  assign tmp41936 = s1 ? tmp41937 : tmp41939;
  assign tmp41942 = s0 ? tmp41921 : tmp40225;
  assign tmp41941 = s1 ? tmp41942 : tmp41869;
  assign tmp41935 = s2 ? tmp41936 : tmp41941;
  assign tmp41946 = l1 ? tmp39541 : tmp41928;
  assign tmp41945 = s0 ? tmp41932 : tmp41946;
  assign tmp41947 = s0 ? tmp41876 : tmp41932;
  assign tmp41944 = ~(s1 ? tmp41945 : tmp41947);
  assign tmp41943 = ~(s2 ? tmp41871 : tmp41944);
  assign tmp41934 = s3 ? tmp41935 : tmp41943;
  assign tmp41918 = s4 ? tmp41919 : tmp41934;
  assign tmp41954 = l1 ? tmp41251 : tmp39587;
  assign tmp41953 = s0 ? tmp41954 : tmp40096;
  assign tmp41952 = s1 ? tmp41953 : tmp41603;
  assign tmp41956 = l1 ? tmp41251 : tmp39630;
  assign tmp41957 = s0 ? tmp41946 : tmp39401;
  assign tmp41955 = s1 ? tmp41956 : tmp41957;
  assign tmp41951 = s2 ? tmp41952 : tmp41955;
  assign tmp41960 = ~(l1 ? tmp39541 : tmp39497);
  assign tmp41959 = s1 ? tmp41854 : tmp41960;
  assign tmp41963 = l1 ? tmp39439 : tmp40534;
  assign tmp41962 = ~(s0 ? tmp41940 : tmp41963);
  assign tmp41961 = ~(s1 ? tmp41890 : tmp41962);
  assign tmp41958 = ~(s2 ? tmp41959 : tmp41961);
  assign tmp41950 = s3 ? tmp41951 : tmp41958;
  assign tmp41968 = l1 ? tmp41251 : tmp39840;
  assign tmp41967 = s0 ? tmp39474 : tmp41968;
  assign tmp41966 = s1 ? tmp41967 : tmp41898;
  assign tmp41969 = ~(l1 ? tmp39375 : tmp40477);
  assign tmp41965 = s2 ? tmp41966 : tmp41969;
  assign tmp41973 = l1 ? tmp39429 : tmp40477;
  assign tmp41972 = s0 ? tmp41973 : tmp41143;
  assign tmp41971 = s1 ? tmp41972 : tmp41960;
  assign tmp41970 = ~(s2 ? tmp41971 : tmp41820);
  assign tmp41964 = s3 ? tmp41965 : tmp41970;
  assign tmp41949 = s4 ? tmp41950 : tmp41964;
  assign tmp41979 = l1 ? tmp39541 : tmp39497;
  assign tmp41978 = s0 ? tmp41979 : tmp39509;
  assign tmp41977 = s1 ? tmp41978 : tmp41910;
  assign tmp41976 = s2 ? tmp41977 : tmp40275;
  assign tmp41983 = ~(l1 ? tmp39429 : tmp39435);
  assign tmp41982 = s0 ? tmp39534 : tmp41983;
  assign tmp41981 = ~(s1 ? tmp39531 : tmp41982);
  assign tmp41980 = ~(s2 ? tmp41828 : tmp41981);
  assign tmp41975 = s3 ? tmp41976 : tmp41980;
  assign tmp41986 = ~(l1 ? tmp39532 : tmp40477);
  assign tmp41985 = s2 ? tmp41913 : tmp41986;
  assign tmp41988 = s1 ? tmp41805 : tmp41126;
  assign tmp41987 = s2 ? tmp41988 : tmp39534;
  assign tmp41984 = s3 ? tmp41985 : tmp41987;
  assign tmp41974 = s4 ? tmp41975 : tmp41984;
  assign tmp41948 = s5 ? tmp41949 : tmp41974;
  assign tmp41917 = s6 ? tmp41918 : tmp41948;
  assign tmp41916 = s7 ? tmp39370 : tmp41917;
  assign tmp41915 = s8 ? tmp41840 : tmp41916;
  assign tmp41752 = s9 ? tmp41753 : tmp41915;
  assign tmp41990 = s8 ? tmp41840 : tmp39370;
  assign tmp41996 = s3 ? tmp41834 : tmp41839;
  assign tmp41995 = s4 ? tmp41822 : tmp41996;
  assign tmp41994 = s5 ? tmp41791 : tmp41995;
  assign tmp41993 = s6 ? tmp41756 : tmp41994;
  assign tmp42000 = s3 ? tmp41985 : tmp41988;
  assign tmp41999 = s4 ? tmp41975 : tmp42000;
  assign tmp41998 = s5 ? tmp41949 : tmp41999;
  assign tmp41997 = s6 ? tmp41918 : tmp41998;
  assign tmp41992 = s7 ? tmp41993 : tmp41997;
  assign tmp42004 = s3 ? tmp41912 : tmp41839;
  assign tmp42003 = s4 ? tmp41905 : tmp42004;
  assign tmp42002 = s5 ? tmp41878 : tmp42003;
  assign tmp42001 = s6 ? tmp41842 : tmp42002;
  assign tmp41991 = s8 ? tmp41992 : tmp42001;
  assign tmp41989 = s9 ? tmp41990 : tmp41991;
  assign tmp41751 = s10 ? tmp41752 : tmp41989;
  assign tmp42008 = s7 ? tmp41755 : tmp41917;
  assign tmp42007 = s8 ? tmp42008 : tmp41841;
  assign tmp42006 = s9 ? tmp41990 : tmp42007;
  assign tmp42005 = s10 ? tmp41752 : tmp42006;
  assign tmp41750 = s11 ? tmp41751 : tmp42005;
  assign tmp42017 = l2 ? tmp39378 : tmp39381;
  assign tmp42016 = l1 ? tmp42017 : tmp40637;
  assign tmp42019 = ~(l1 ? tmp39384 : tmp39409);
  assign tmp42018 = ~(s0 ? tmp39422 : tmp42019);
  assign tmp42015 = s1 ? tmp42016 : tmp42018;
  assign tmp42023 = ~(l1 ? tmp42017 : tmp40642);
  assign tmp42022 = s0 ? tmp41570 : tmp42023;
  assign tmp42024 = s0 ? tmp41573 : tmp42023;
  assign tmp42021 = s1 ? tmp42022 : tmp42024;
  assign tmp42027 = l1 ? tmp42017 : tmp40642;
  assign tmp42029 = l2 ? tmp39376 : tmp39379;
  assign tmp42028 = ~(l1 ? tmp42029 : tmp39388);
  assign tmp42026 = ~(s0 ? tmp42027 : tmp42028);
  assign tmp42025 = s1 ? tmp41575 : tmp42026;
  assign tmp42020 = ~(s2 ? tmp42021 : tmp42025);
  assign tmp42014 = s3 ? tmp42015 : tmp42020;
  assign tmp42034 = l1 ? tmp42029 : tmp39388;
  assign tmp42033 = ~(s0 ? tmp42034 : tmp42023);
  assign tmp42032 = s1 ? tmp41582 : tmp42033;
  assign tmp42036 = s0 ? tmp42016 : tmp40225;
  assign tmp42035 = s1 ? tmp42036 : tmp41587;
  assign tmp42031 = s2 ? tmp42032 : tmp42035;
  assign tmp42039 = l1 ? tmp39527 : tmp39429;
  assign tmp42038 = s1 ? tmp39422 : tmp42039;
  assign tmp42043 = l2 ? tmp39378 : tmp39403;
  assign tmp42042 = l1 ? tmp42043 : tmp40642;
  assign tmp42041 = s0 ? tmp42027 : tmp42042;
  assign tmp42045 = l1 ? tmp39501 : tmp39434;
  assign tmp42044 = s0 ? tmp42045 : tmp42027;
  assign tmp42040 = ~(s1 ? tmp42041 : tmp42044);
  assign tmp42037 = ~(s2 ? tmp42038 : tmp42040);
  assign tmp42030 = s3 ? tmp42031 : tmp42037;
  assign tmp42013 = s4 ? tmp42014 : tmp42030;
  assign tmp42051 = s0 ? tmp41564 : tmp40096;
  assign tmp42050 = s1 ? tmp42051 : tmp41603;
  assign tmp42053 = s0 ? tmp42042 : tmp39401;
  assign tmp42052 = s1 ? tmp39486 : tmp42053;
  assign tmp42049 = s2 ? tmp42050 : tmp42052;
  assign tmp42056 = ~(l1 ? tmp42043 : tmp39434);
  assign tmp42055 = s1 ? tmp41573 : tmp42056;
  assign tmp42059 = l1 ? tmp39501 : tmp39378;
  assign tmp42058 = s0 ? tmp42045 : tmp42059;
  assign tmp42061 = l1 ? tmp42029 : tmp39621;
  assign tmp42060 = ~(s0 ? tmp42034 : tmp42061);
  assign tmp42057 = ~(s1 ? tmp42058 : tmp42060);
  assign tmp42054 = ~(s2 ? tmp42055 : tmp42057);
  assign tmp42048 = s3 ? tmp42049 : tmp42054;
  assign tmp42066 = l1 ? tmp42017 : tmp39527;
  assign tmp42065 = s0 ? tmp42045 : tmp42066;
  assign tmp42064 = s1 ? tmp42065 : tmp41620;
  assign tmp42063 = s2 ? tmp42064 : tmp39387;
  assign tmp42070 = ~(l1 ? tmp42043 : tmp39527);
  assign tmp42069 = s0 ? tmp40269 : tmp42070;
  assign tmp42068 = s1 ? tmp42069 : tmp42056;
  assign tmp42071 = s1 ? 1 : tmp42039;
  assign tmp42067 = ~(s2 ? tmp42068 : tmp42071);
  assign tmp42062 = s3 ? tmp42063 : tmp42067;
  assign tmp42047 = s4 ? tmp42048 : tmp42062;
  assign tmp42077 = l1 ? tmp42043 : tmp39434;
  assign tmp42078 = ~(l1 ? tmp39513 : 1);
  assign tmp42076 = s0 ? tmp42077 : tmp42078;
  assign tmp42079 = ~(l1 ? tmp39532 : tmp39375);
  assign tmp42075 = s1 ? tmp42076 : tmp42079;
  assign tmp42074 = s2 ? tmp42075 : tmp40275;
  assign tmp42081 = s1 ? tmp41836 : tmp39528;
  assign tmp42084 = l1 ? tmp39501 : tmp39527;
  assign tmp42083 = s0 ? tmp39512 : tmp42084;
  assign tmp42082 = ~(s1 ? tmp42083 : tmp39999);
  assign tmp42080 = ~(s2 ? tmp42081 : tmp42082);
  assign tmp42073 = s3 ? tmp42074 : tmp42080;
  assign tmp42087 = s1 ? tmp41638 : tmp42045;
  assign tmp42088 = ~(l1 ? tmp40982 : tmp39388);
  assign tmp42086 = s2 ? tmp42087 : tmp42088;
  assign tmp42090 = l1 ? 1 : tmp39434;
  assign tmp42092 = ~(l1 ? tmp40982 : tmp39630);
  assign tmp42091 = s0 ? tmp39512 : tmp42092;
  assign tmp42089 = s1 ? tmp42090 : tmp42091;
  assign tmp42085 = s3 ? tmp42086 : tmp42089;
  assign tmp42072 = s4 ? tmp42073 : tmp42085;
  assign tmp42046 = s5 ? tmp42047 : tmp42072;
  assign tmp42012 = s6 ? tmp42013 : tmp42046;
  assign tmp42011 = s7 ? tmp39370 : tmp42012;
  assign tmp42094 = s8 ? tmp42011 : tmp39370;
  assign tmp42099 = s1 ? tmp42090 : tmp42092;
  assign tmp42098 = s3 ? tmp42086 : tmp42099;
  assign tmp42097 = s4 ? tmp42073 : tmp42098;
  assign tmp42096 = s5 ? tmp42047 : tmp42097;
  assign tmp42095 = s6 ? tmp42013 : tmp42096;
  assign tmp42093 = s9 ? tmp42094 : tmp42095;
  assign tmp42010 = s10 ? tmp42011 : tmp42093;
  assign tmp42101 = s9 ? tmp42094 : tmp42012;
  assign tmp42100 = s10 ? tmp42011 : tmp42101;
  assign tmp42009 = s11 ? tmp42010 : tmp42100;
  assign tmp41749 = s12 ? tmp41750 : tmp42009;
  assign tmp41555 = s13 ? tmp41556 : tmp41749;
  assign tmp42113 = l1 ? tmp40901 : tmp39575;
  assign tmp42115 = ~(l1 ? tmp40905 : tmp39575);
  assign tmp42114 = ~(s0 ? tmp39946 : tmp42115);
  assign tmp42112 = s1 ? tmp42113 : tmp42114;
  assign tmp42119 = l2 ? tmp39440 : tmp39381;
  assign tmp42118 = ~(l1 ? tmp40910 : tmp42119);
  assign tmp42117 = s0 ? tmp39946 : tmp42118;
  assign tmp42121 = s0 ? tmp39946 : tmp39420;
  assign tmp42123 = l1 ? tmp40910 : tmp42119;
  assign tmp42125 = ~(l2 ? tmp39440 : tmp39381);
  assign tmp42124 = ~(l1 ? tmp39480 : tmp42125);
  assign tmp42122 = ~(s0 ? tmp42123 : tmp42124);
  assign tmp42120 = s1 ? tmp42121 : tmp42122;
  assign tmp42116 = ~(s2 ? tmp42117 : tmp42120);
  assign tmp42111 = s3 ? tmp42112 : tmp42116;
  assign tmp42129 = s0 ? tmp39928 : tmp40655;
  assign tmp42131 = l1 ? tmp39480 : tmp42125;
  assign tmp42130 = ~(s0 ? tmp42131 : tmp42118);
  assign tmp42128 = s1 ? tmp42129 : tmp42130;
  assign tmp42133 = s0 ? tmp42113 : tmp40225;
  assign tmp42132 = s1 ? tmp42133 : tmp40660;
  assign tmp42127 = s2 ? tmp42128 : tmp42132;
  assign tmp42136 = l1 ? 1 : tmp39527;
  assign tmp42135 = s1 ? tmp39946 : tmp42136;
  assign tmp42139 = l1 ? tmp40933 : tmp42119;
  assign tmp42138 = s0 ? tmp42123 : tmp42139;
  assign tmp42141 = l1 ? tmp39379 : tmp41675;
  assign tmp42140 = s0 ? tmp42141 : tmp42123;
  assign tmp42137 = ~(s1 ? tmp42138 : tmp42140);
  assign tmp42134 = ~(s2 ? tmp42135 : tmp42137);
  assign tmp42126 = s3 ? tmp42127 : tmp42134;
  assign tmp42110 = s4 ? tmp42111 : tmp42126;
  assign tmp42148 = l1 ? tmp40905 : tmp39575;
  assign tmp42147 = s0 ? tmp42148 : tmp40096;
  assign tmp42146 = s1 ? tmp42147 : tmp40655;
  assign tmp42150 = l1 ? tmp40905 : tmp39621;
  assign tmp42151 = s0 ? tmp42139 : tmp39401;
  assign tmp42149 = s1 ? tmp42150 : tmp42151;
  assign tmp42145 = s2 ? tmp42146 : tmp42149;
  assign tmp42155 = l2 ? tmp39440 : tmp39403;
  assign tmp42154 = ~(l1 ? tmp39379 : tmp42155);
  assign tmp42153 = s1 ? tmp39946 : tmp42154;
  assign tmp42157 = s0 ? tmp42141 : tmp39626;
  assign tmp42159 = l1 ? tmp39480 : tmp39527;
  assign tmp42158 = ~(s0 ? tmp42131 : tmp42159);
  assign tmp42156 = ~(s1 ? tmp42157 : tmp42158);
  assign tmp42152 = ~(s2 ? tmp42153 : tmp42156);
  assign tmp42144 = s3 ? tmp42145 : tmp42152;
  assign tmp42164 = l1 ? tmp39378 : tmp41738;
  assign tmp42165 = l1 ? tmp40910 : tmp39621;
  assign tmp42163 = s0 ? tmp42164 : tmp42165;
  assign tmp42162 = s1 ? tmp42163 : tmp40695;
  assign tmp42166 = ~(s1 ? tmp39495 : tmp39939);
  assign tmp42161 = s2 ? tmp42162 : tmp42166;
  assign tmp42170 = ~(l1 ? tmp39439 : tmp39621);
  assign tmp42169 = s0 ? tmp39939 : tmp42170;
  assign tmp42173 = l2 ? tmp39379 : tmp39403;
  assign tmp42172 = ~(l1 ? tmp39379 : tmp42173);
  assign tmp42171 = s0 ? tmp39495 : tmp42172;
  assign tmp42168 = s1 ? tmp42169 : tmp42171;
  assign tmp42174 = s1 ? tmp39651 : tmp42136;
  assign tmp42167 = ~(s2 ? tmp42168 : tmp42174);
  assign tmp42160 = s3 ? tmp42161 : tmp42167;
  assign tmp42143 = s4 ? tmp42144 : tmp42160;
  assign tmp42180 = l1 ? tmp39379 : tmp42155;
  assign tmp42179 = s0 ? tmp42180 : 0;
  assign tmp42178 = s1 ? tmp42179 : 0;
  assign tmp42177 = s2 ? tmp42178 : tmp41314;
  assign tmp42183 = s0 ? tmp39480 : tmp42136;
  assign tmp42182 = s1 ? tmp42183 : tmp39664;
  assign tmp42184 = ~(s1 ? tmp39534 : tmp39535);
  assign tmp42181 = ~(s2 ? tmp42182 : tmp42184);
  assign tmp42176 = s3 ? tmp42177 : tmp42181;
  assign tmp42189 = ~(l1 ? tmp40982 : 1);
  assign tmp42188 = s0 ? tmp39540 : tmp42189;
  assign tmp42190 = ~(l1 ? tmp39379 : tmp41675);
  assign tmp42187 = s1 ? tmp42188 : tmp42190;
  assign tmp42191 = s1 ? tmp39939 : tmp39480;
  assign tmp42186 = s2 ? tmp42187 : tmp42191;
  assign tmp42194 = l1 ? tmp40982 : tmp39501;
  assign tmp42195 = ~(l1 ? tmp39480 : tmp39527);
  assign tmp42193 = s1 ? tmp42194 : tmp42195;
  assign tmp42192 = ~(s2 ? tmp42193 : tmp39559);
  assign tmp42185 = ~(s3 ? tmp42186 : tmp42192);
  assign tmp42175 = s4 ? tmp42176 : tmp42185;
  assign tmp42142 = s5 ? tmp42143 : tmp42175;
  assign tmp42109 = s6 ? tmp42110 : tmp42142;
  assign tmp42108 = s7 ? tmp39370 : tmp42109;
  assign tmp42201 = l1 ? tmp40992 : tmp39575;
  assign tmp42203 = ~(l1 ? tmp40997 : tmp39575);
  assign tmp42202 = ~(s0 ? tmp40037 : tmp42203);
  assign tmp42200 = s1 ? tmp42201 : tmp42202;
  assign tmp42206 = ~(l1 ? tmp41002 : tmp42119);
  assign tmp42205 = s0 ? tmp40037 : tmp42206;
  assign tmp42208 = s0 ? tmp40037 : tmp41336;
  assign tmp42210 = l1 ? tmp41002 : tmp42119;
  assign tmp42211 = ~(l1 ? tmp39403 : tmp42125);
  assign tmp42209 = ~(s0 ? tmp42210 : tmp42211);
  assign tmp42207 = s1 ? tmp42208 : tmp42209;
  assign tmp42204 = ~(s2 ? tmp42205 : tmp42207);
  assign tmp42199 = s3 ? tmp42200 : tmp42204;
  assign tmp42215 = s0 ? tmp40021 : tmp40749;
  assign tmp42217 = l1 ? tmp39403 : tmp42125;
  assign tmp42216 = ~(s0 ? tmp42217 : tmp42206);
  assign tmp42214 = s1 ? tmp42215 : tmp42216;
  assign tmp42219 = s0 ? tmp42201 : tmp40225;
  assign tmp42220 = l1 ? tmp39385 : tmp39375;
  assign tmp42218 = s1 ? tmp42219 : tmp42220;
  assign tmp42213 = s2 ? tmp42214 : tmp42218;
  assign tmp42222 = s1 ? tmp40037 : tmp42136;
  assign tmp42225 = l1 ? tmp39379 : tmp42119;
  assign tmp42224 = s0 ? tmp42210 : tmp42225;
  assign tmp42226 = s0 ? tmp42141 : tmp42210;
  assign tmp42223 = ~(s1 ? tmp42224 : tmp42226);
  assign tmp42221 = ~(s2 ? tmp42222 : tmp42223);
  assign tmp42212 = s3 ? tmp42213 : tmp42221;
  assign tmp42198 = s4 ? tmp42199 : tmp42212;
  assign tmp42233 = l1 ? tmp40997 : tmp39575;
  assign tmp42232 = s0 ? tmp42233 : tmp40096;
  assign tmp42231 = s1 ? tmp42232 : tmp40749;
  assign tmp42235 = l1 ? tmp40997 : tmp39621;
  assign tmp42236 = s0 ? tmp42225 : tmp40024;
  assign tmp42234 = s1 ? tmp42235 : tmp42236;
  assign tmp42230 = s2 ? tmp42231 : tmp42234;
  assign tmp42238 = s1 ? tmp40037 : tmp42154;
  assign tmp42241 = l1 ? tmp39403 : tmp39527;
  assign tmp42240 = ~(s0 ? tmp42217 : tmp42241);
  assign tmp42239 = ~(s1 ? tmp42157 : tmp42240);
  assign tmp42237 = ~(s2 ? tmp42238 : tmp42239);
  assign tmp42229 = s3 ? tmp42230 : tmp42237;
  assign tmp42246 = l1 ? tmp41002 : tmp39621;
  assign tmp42245 = s0 ? tmp42164 : tmp42246;
  assign tmp42247 = s0 ? tmp39483 : tmp41015;
  assign tmp42244 = s1 ? tmp42245 : tmp42247;
  assign tmp42248 = ~(l1 ? tmp39403 : tmp39801);
  assign tmp42243 = s2 ? tmp42244 : tmp42248;
  assign tmp42252 = ~(l1 ? tmp39475 : tmp39621);
  assign tmp42251 = s0 ? tmp39939 : tmp42252;
  assign tmp42250 = s1 ? tmp42251 : tmp42172;
  assign tmp42249 = ~(s2 ? tmp42250 : tmp42174);
  assign tmp42242 = s3 ? tmp42243 : tmp42249;
  assign tmp42228 = s4 ? tmp42229 : tmp42242;
  assign tmp42255 = s2 ? tmp42178 : tmp41390;
  assign tmp42254 = s3 ? tmp42255 : tmp42181;
  assign tmp42253 = s4 ? tmp42254 : tmp42185;
  assign tmp42227 = s5 ? tmp42228 : tmp42253;
  assign tmp42197 = s6 ? tmp42198 : tmp42227;
  assign tmp42196 = s7 ? tmp39370 : tmp42197;
  assign tmp42107 = s8 ? tmp42108 : tmp42196;
  assign tmp42262 = l1 ? tmp40992 : tmp39587;
  assign tmp42264 = ~(l1 ? tmp40997 : tmp39587);
  assign tmp42263 = ~(s0 ? tmp40731 : tmp42264);
  assign tmp42261 = s1 ? tmp42262 : tmp42263;
  assign tmp42268 = l2 ? tmp39379 : tmp39381;
  assign tmp42267 = ~(l1 ? tmp41002 : tmp42268);
  assign tmp42266 = s0 ? tmp41408 : tmp42267;
  assign tmp42270 = s0 ? tmp41408 : tmp39420;
  assign tmp42272 = l1 ? tmp41002 : tmp42268;
  assign tmp42274 = ~(l2 ? tmp39379 : tmp39381);
  assign tmp42273 = ~(l1 ? tmp39403 : tmp42274);
  assign tmp42271 = ~(s0 ? tmp42272 : tmp42273);
  assign tmp42269 = s1 ? tmp42270 : tmp42271;
  assign tmp42265 = ~(s2 ? tmp42266 : tmp42269);
  assign tmp42260 = s3 ? tmp42261 : tmp42265;
  assign tmp42279 = l1 ? tmp39972 : tmp39587;
  assign tmp42278 = s0 ? tmp42279 : tmp40749;
  assign tmp42281 = l1 ? tmp39403 : tmp42274;
  assign tmp42280 = ~(s0 ? tmp42281 : tmp42267);
  assign tmp42277 = s1 ? tmp42278 : tmp42280;
  assign tmp42283 = s0 ? tmp42262 : tmp40225;
  assign tmp42282 = s1 ? tmp42283 : tmp39428;
  assign tmp42276 = s2 ? tmp42277 : tmp42282;
  assign tmp42285 = s1 ? tmp40731 : tmp42136;
  assign tmp42288 = l1 ? tmp39379 : tmp42268;
  assign tmp42287 = s0 ? tmp42272 : tmp42288;
  assign tmp42290 = l1 ? tmp39379 : tmp41738;
  assign tmp42289 = s0 ? tmp42290 : tmp42272;
  assign tmp42286 = ~(s1 ? tmp42287 : tmp42289);
  assign tmp42284 = ~(s2 ? tmp42285 : tmp42286);
  assign tmp42275 = s3 ? tmp42276 : tmp42284;
  assign tmp42259 = s4 ? tmp42260 : tmp42275;
  assign tmp42297 = l1 ? tmp40997 : tmp39587;
  assign tmp42296 = s0 ? tmp42297 : tmp40096;
  assign tmp42295 = s1 ? tmp42296 : tmp41440;
  assign tmp42299 = l1 ? tmp40997 : tmp39630;
  assign tmp42300 = s0 ? tmp42288 : tmp39401;
  assign tmp42298 = s1 ? tmp42299 : tmp42300;
  assign tmp42294 = s2 ? tmp42295 : tmp42298;
  assign tmp42302 = s1 ? tmp41408 : tmp42172;
  assign tmp42304 = s0 ? tmp42290 : tmp39626;
  assign tmp42306 = l1 ? tmp39403 : tmp39684;
  assign tmp42305 = ~(s0 ? tmp42281 : tmp42306);
  assign tmp42303 = ~(s1 ? tmp42304 : tmp42305);
  assign tmp42301 = ~(s2 ? tmp42302 : tmp42303);
  assign tmp42293 = s3 ? tmp42294 : tmp42301;
  assign tmp42311 = l1 ? tmp41002 : tmp39630;
  assign tmp42310 = s0 ? tmp42164 : tmp42311;
  assign tmp42309 = s1 ? tmp42310 : tmp39482;
  assign tmp42312 = ~(l1 ? tmp39403 : tmp40477);
  assign tmp42308 = s2 ? tmp42309 : tmp42312;
  assign tmp42316 = l1 ? tmp39480 : tmp40477;
  assign tmp42317 = ~(l1 ? tmp39475 : tmp39630);
  assign tmp42315 = s0 ? tmp42316 : tmp42317;
  assign tmp42314 = s1 ? tmp42315 : tmp42172;
  assign tmp42313 = ~(s2 ? tmp42314 : tmp42174);
  assign tmp42307 = s3 ? tmp42308 : tmp42313;
  assign tmp42292 = s4 ? tmp42293 : tmp42307;
  assign tmp42323 = l1 ? tmp39379 : tmp42173;
  assign tmp42322 = s0 ? tmp42323 : 0;
  assign tmp42321 = s1 ? tmp42322 : tmp39720;
  assign tmp42320 = s2 ? tmp42321 : tmp41464;
  assign tmp42319 = s3 ? tmp42320 : tmp42181;
  assign tmp42327 = ~(l1 ? tmp39379 : tmp41738);
  assign tmp42326 = s1 ? tmp42188 : tmp42327;
  assign tmp42328 = s1 ? tmp42316 : tmp39480;
  assign tmp42325 = s2 ? tmp42326 : tmp42328;
  assign tmp42324 = ~(s3 ? tmp42325 : tmp42192);
  assign tmp42318 = s4 ? tmp42319 : tmp42324;
  assign tmp42291 = s5 ? tmp42292 : tmp42318;
  assign tmp42258 = s6 ? tmp42259 : tmp42291;
  assign tmp42257 = s7 ? tmp39370 : tmp42258;
  assign tmp42256 = s8 ? tmp42196 : tmp42257;
  assign tmp42106 = s9 ? tmp42107 : tmp42256;
  assign tmp42336 = s0 ? tmp40731 : tmp42267;
  assign tmp42338 = s0 ? tmp40731 : tmp39420;
  assign tmp42337 = s1 ? tmp42338 : tmp42271;
  assign tmp42335 = ~(s2 ? tmp42336 : tmp42337);
  assign tmp42334 = s3 ? tmp42261 : tmp42335;
  assign tmp42333 = s4 ? tmp42334 : tmp42275;
  assign tmp42343 = s1 ? tmp42296 : tmp41510;
  assign tmp42342 = s2 ? tmp42343 : tmp42298;
  assign tmp42345 = s1 ? tmp40731 : tmp42172;
  assign tmp42344 = ~(s2 ? tmp42345 : tmp42303);
  assign tmp42341 = s3 ? tmp42342 : tmp42344;
  assign tmp42340 = s4 ? tmp42341 : tmp42307;
  assign tmp42348 = s2 ? tmp42321 : tmp41314;
  assign tmp42347 = s3 ? tmp42348 : tmp42181;
  assign tmp42346 = s4 ? tmp42347 : tmp42324;
  assign tmp42339 = s5 ? tmp42340 : tmp42346;
  assign tmp42332 = s6 ? tmp42333 : tmp42339;
  assign tmp42331 = s7 ? tmp39370 : tmp42332;
  assign tmp42330 = s8 ? tmp42331 : tmp39370;
  assign tmp42356 = s1 ? tmp42169 : tmp42172;
  assign tmp42355 = ~(s2 ? tmp42356 : tmp42174);
  assign tmp42354 = s3 ? tmp42161 : tmp42355;
  assign tmp42353 = s4 ? tmp42144 : tmp42354;
  assign tmp42359 = s2 ? tmp42187 : tmp39939;
  assign tmp42360 = ~(s1 ? tmp42194 : tmp42195);
  assign tmp42358 = ~(s3 ? tmp42359 : tmp42360);
  assign tmp42357 = s4 ? tmp42176 : tmp42358;
  assign tmp42352 = s5 ? tmp42353 : tmp42357;
  assign tmp42351 = s6 ? tmp42110 : tmp42352;
  assign tmp42365 = s2 ? tmp42326 : tmp42316;
  assign tmp42364 = ~(s3 ? tmp42365 : tmp42360);
  assign tmp42363 = s4 ? tmp42319 : tmp42364;
  assign tmp42362 = s5 ? tmp42292 : tmp42363;
  assign tmp42361 = s6 ? tmp42259 : tmp42362;
  assign tmp42350 = s7 ? tmp42351 : tmp42361;
  assign tmp42369 = s4 ? tmp42254 : tmp42358;
  assign tmp42368 = s5 ? tmp42228 : tmp42369;
  assign tmp42367 = s6 ? tmp42198 : tmp42368;
  assign tmp42372 = s4 ? tmp42347 : tmp42364;
  assign tmp42371 = s5 ? tmp42340 : tmp42372;
  assign tmp42370 = s6 ? tmp42333 : tmp42371;
  assign tmp42366 = s7 ? tmp42367 : tmp42370;
  assign tmp42349 = s8 ? tmp42350 : tmp42366;
  assign tmp42329 = s9 ? tmp42330 : tmp42349;
  assign tmp42105 = s10 ? tmp42106 : tmp42329;
  assign tmp42376 = s7 ? tmp42109 : tmp42258;
  assign tmp42377 = s7 ? tmp42197 : tmp42332;
  assign tmp42375 = s8 ? tmp42376 : tmp42377;
  assign tmp42374 = s9 ? tmp42330 : tmp42375;
  assign tmp42373 = s10 ? tmp42106 : tmp42374;
  assign tmp42104 = s11 ? tmp42105 : tmp42373;
  assign tmp42387 = l1 ? tmp42119 : tmp40633;
  assign tmp42389 = ~(l2 ? tmp39376 : tmp40634);
  assign tmp42388 = ~(s0 ? tmp39477 : tmp42389);
  assign tmp42386 = s1 ? tmp42387 : tmp42388;
  assign tmp42392 = s0 ? tmp39786 : tmp40649;
  assign tmp42394 = l1 ? tmp39513 : tmp39478;
  assign tmp42393 = s0 ? tmp42394 : tmp40649;
  assign tmp42391 = s1 ? tmp42392 : tmp42393;
  assign tmp42396 = s0 ? tmp42394 : tmp39420;
  assign tmp42398 = ~(l1 ? tmp39513 : tmp40649);
  assign tmp42397 = ~(s0 ? tmp40643 : tmp42398);
  assign tmp42395 = s1 ? tmp42396 : tmp42397;
  assign tmp42390 = ~(s2 ? tmp42391 : tmp42395);
  assign tmp42385 = s3 ? tmp42386 : tmp42390;
  assign tmp42403 = l1 ? tmp39575 : tmp40633;
  assign tmp42402 = s0 ? tmp42403 : tmp40024;
  assign tmp42405 = l1 ? tmp39513 : tmp40649;
  assign tmp42404 = ~(s0 ? tmp42405 : tmp40649);
  assign tmp42401 = s1 ? tmp42402 : tmp42404;
  assign tmp42407 = s0 ? tmp42387 : tmp40225;
  assign tmp42406 = s1 ? tmp42407 : tmp39569;
  assign tmp42400 = s2 ? tmp42401 : tmp42406;
  assign tmp42409 = s1 ? tmp39477 : tmp39513;
  assign tmp42412 = l1 ? tmp40683 : tmp40643;
  assign tmp42411 = s0 ? tmp40643 : tmp42412;
  assign tmp42414 = l1 ? tmp40693 : tmp40668;
  assign tmp42413 = s0 ? tmp42414 : tmp40643;
  assign tmp42410 = ~(s1 ? tmp42411 : tmp42413);
  assign tmp42408 = ~(s2 ? tmp42409 : tmp42410);
  assign tmp42399 = s3 ? tmp42400 : tmp42408;
  assign tmp42384 = s4 ? tmp42385 : tmp42399;
  assign tmp42420 = s0 ? tmp40633 : tmp40096;
  assign tmp42419 = s1 ? tmp42420 : tmp40096;
  assign tmp42422 = l1 ? tmp40633 : tmp39376;
  assign tmp42423 = s0 ? tmp42412 : tmp39401;
  assign tmp42421 = s1 ? tmp42422 : tmp42423;
  assign tmp42418 = s2 ? tmp42419 : tmp42421;
  assign tmp42426 = ~(l1 ? tmp40705 : tmp40683);
  assign tmp42425 = s1 ? tmp42394 : tmp42426;
  assign tmp42429 = l1 ? tmp39604 : tmp39501;
  assign tmp42428 = s0 ? tmp42414 : tmp42429;
  assign tmp42430 = ~(s0 ? tmp42405 : tmp39513);
  assign tmp42427 = ~(s1 ? tmp42428 : tmp42430);
  assign tmp42424 = ~(s2 ? tmp42425 : tmp42427);
  assign tmp42417 = s3 ? tmp42418 : tmp42424;
  assign tmp42435 = l1 ? tmp39501 : tmp40693;
  assign tmp42436 = l1 ? tmp40643 : tmp39376;
  assign tmp42434 = s0 ? tmp42435 : tmp42436;
  assign tmp42433 = s1 ? tmp42434 : tmp41813;
  assign tmp42432 = s2 ? tmp42433 : tmp40096;
  assign tmp42440 = ~(l1 ? tmp42155 : tmp39376);
  assign tmp42439 = s0 ? tmp39786 : tmp42440;
  assign tmp42441 = ~(l2 ? tmp39379 : tmp39376);
  assign tmp42438 = s1 ? tmp42439 : tmp42441;
  assign tmp42442 = s1 ? tmp39651 : tmp39513;
  assign tmp42437 = ~(s2 ? tmp42438 : tmp42442);
  assign tmp42431 = s3 ? tmp42432 : tmp42437;
  assign tmp42416 = s4 ? tmp42417 : tmp42431;
  assign tmp42448 = l1 ? tmp40705 : tmp40683;
  assign tmp42447 = s0 ? tmp42448 : tmp42078;
  assign tmp42446 = s1 ? tmp42447 : tmp42078;
  assign tmp42450 = s0 ? tmp39516 : tmp40880;
  assign tmp42449 = ~(s1 ? tmp42450 : 1);
  assign tmp42445 = s2 ? tmp42446 : tmp42449;
  assign tmp42453 = l1 ? tmp39501 : tmp39430;
  assign tmp42452 = ~(s1 ? tmp42453 : 0);
  assign tmp42451 = ~(s2 ? tmp41635 : tmp42452);
  assign tmp42444 = s3 ? tmp42445 : tmp42451;
  assign tmp42457 = l1 ? tmp39430 : tmp39435;
  assign tmp42456 = s1 ? tmp42457 : tmp42414;
  assign tmp42458 = ~(l1 ? tmp39513 : tmp39478);
  assign tmp42455 = s2 ? tmp42456 : tmp42458;
  assign tmp42461 = ~(l1 ? tmp39430 : tmp39604);
  assign tmp42460 = s0 ? tmp39516 : tmp42461;
  assign tmp42459 = ~(s1 ? tmp42460 : tmp39513);
  assign tmp42454 = s3 ? tmp42455 : tmp42459;
  assign tmp42443 = s4 ? tmp42444 : tmp42454;
  assign tmp42415 = s5 ? tmp42416 : tmp42443;
  assign tmp42383 = s6 ? tmp42384 : tmp42415;
  assign tmp42382 = s7 ? tmp39370 : tmp42383;
  assign tmp42467 = l1 ? tmp42268 : tmp40633;
  assign tmp42469 = ~(l1 ? tmp40729 : tmp40633);
  assign tmp42468 = ~(s0 ? tmp39477 : tmp42469);
  assign tmp42466 = s1 ? tmp42467 : tmp42468;
  assign tmp42473 = ~(l1 ? tmp40737 : tmp40643);
  assign tmp42472 = s0 ? tmp39477 : tmp42473;
  assign tmp42475 = l1 ? tmp40779 : tmp39478;
  assign tmp42474 = s0 ? tmp42475 : tmp42473;
  assign tmp42471 = s1 ? tmp42472 : tmp42474;
  assign tmp42477 = s0 ? tmp42475 : tmp41336;
  assign tmp42479 = l1 ? tmp40737 : tmp40643;
  assign tmp42480 = ~(l1 ? tmp40779 : tmp40649);
  assign tmp42478 = ~(s0 ? tmp42479 : tmp42480);
  assign tmp42476 = s1 ? tmp42477 : tmp42478;
  assign tmp42470 = ~(s2 ? tmp42471 : tmp42476);
  assign tmp42465 = s3 ? tmp42466 : tmp42470;
  assign tmp42485 = l1 ? tmp39587 : tmp40633;
  assign tmp42484 = s0 ? tmp42485 : tmp40024;
  assign tmp42487 = l1 ? tmp40779 : tmp40649;
  assign tmp42486 = ~(s0 ? tmp42487 : tmp42473);
  assign tmp42483 = s1 ? tmp42484 : tmp42486;
  assign tmp42489 = s0 ? tmp42467 : tmp40225;
  assign tmp42488 = s1 ? tmp42489 : tmp39569;
  assign tmp42482 = s2 ? tmp42483 : tmp42488;
  assign tmp42493 = l1 ? tmp40705 : tmp40643;
  assign tmp42492 = s0 ? tmp42479 : tmp42493;
  assign tmp42494 = s0 ? tmp42414 : tmp42479;
  assign tmp42491 = ~(s1 ? tmp42492 : tmp42494);
  assign tmp42490 = ~(s2 ? tmp42409 : tmp42491);
  assign tmp42481 = s3 ? tmp42482 : tmp42490;
  assign tmp42464 = s4 ? tmp42465 : tmp42481;
  assign tmp42501 = l1 ? tmp40729 : tmp40633;
  assign tmp42500 = s0 ? tmp42501 : tmp40096;
  assign tmp42499 = s1 ? tmp42500 : tmp40024;
  assign tmp42503 = l1 ? tmp40729 : tmp39376;
  assign tmp42504 = s0 ? tmp42493 : tmp40024;
  assign tmp42502 = s1 ? tmp42503 : tmp42504;
  assign tmp42498 = s2 ? tmp42499 : tmp42502;
  assign tmp42506 = s1 ? tmp42475 : tmp42426;
  assign tmp42509 = l1 ? tmp40779 : tmp39513;
  assign tmp42508 = ~(s0 ? tmp42487 : tmp42509);
  assign tmp42507 = ~(s1 ? tmp42428 : tmp42508);
  assign tmp42505 = ~(s2 ? tmp42506 : tmp42507);
  assign tmp42497 = s3 ? tmp42498 : tmp42505;
  assign tmp42514 = l1 ? tmp40737 : tmp39376;
  assign tmp42513 = s0 ? tmp42435 : tmp42514;
  assign tmp42512 = s1 ? tmp42513 : tmp41813;
  assign tmp42511 = s2 ? tmp42512 : tmp40024;
  assign tmp42518 = ~(l1 ? tmp42173 : tmp39376);
  assign tmp42517 = s0 ? tmp39786 : tmp42518;
  assign tmp42516 = s1 ? tmp42517 : tmp42441;
  assign tmp42515 = ~(s2 ? tmp42516 : tmp42442);
  assign tmp42510 = s3 ? tmp42511 : tmp42515;
  assign tmp42496 = s4 ? tmp42497 : tmp42510;
  assign tmp42523 = l1 ? tmp39630 : tmp39403;
  assign tmp42522 = s1 ? tmp42523 : 0;
  assign tmp42521 = s2 ? tmp42446 : tmp42522;
  assign tmp42520 = s3 ? tmp42521 : tmp42451;
  assign tmp42526 = l1 ? tmp39430 : tmp39604;
  assign tmp42527 = ~(l2 ? 1 : tmp39378);
  assign tmp42525 = s1 ? tmp42526 : tmp42527;
  assign tmp42524 = s3 ? tmp42455 : tmp42525;
  assign tmp42519 = s4 ? tmp42520 : tmp42524;
  assign tmp42495 = s5 ? tmp42496 : tmp42519;
  assign tmp42463 = s6 ? tmp42464 : tmp42495;
  assign tmp42462 = s7 ? tmp39370 : tmp42463;
  assign tmp42381 = s8 ? tmp42382 : tmp42462;
  assign tmp42534 = l1 ? tmp42268 : tmp40816;
  assign tmp42536 = ~(l1 ? tmp40729 : tmp40816);
  assign tmp42535 = ~(s0 ? tmp41847 : tmp42536);
  assign tmp42533 = s1 ? tmp42534 : tmp42535;
  assign tmp42540 = l1 ? tmp39402 : tmp39518;
  assign tmp42541 = ~(l1 ? tmp40737 : tmp40823);
  assign tmp42539 = s0 ? tmp42540 : tmp42541;
  assign tmp42543 = l1 ? tmp40779 : tmp39518;
  assign tmp42542 = s0 ? tmp42543 : tmp42541;
  assign tmp42538 = s1 ? tmp42539 : tmp42542;
  assign tmp42545 = s0 ? tmp42543 : tmp39420;
  assign tmp42547 = l1 ? tmp40737 : tmp40823;
  assign tmp42548 = ~(l1 ? tmp40779 : tmp40829);
  assign tmp42546 = ~(s0 ? tmp42547 : tmp42548);
  assign tmp42544 = s1 ? tmp42545 : tmp42546;
  assign tmp42537 = ~(s2 ? tmp42538 : tmp42544);
  assign tmp42532 = s3 ? tmp42533 : tmp42537;
  assign tmp42553 = l1 ? tmp39587 : tmp40816;
  assign tmp42552 = s0 ? tmp42553 : tmp40024;
  assign tmp42555 = l1 ? tmp40779 : tmp40829;
  assign tmp42554 = ~(s0 ? tmp42555 : tmp42541);
  assign tmp42551 = s1 ? tmp42552 : tmp42554;
  assign tmp42557 = s0 ? tmp42534 : tmp40225;
  assign tmp42556 = s1 ? tmp42557 : tmp41869;
  assign tmp42550 = s2 ? tmp42551 : tmp42556;
  assign tmp42559 = s1 ? tmp41847 : tmp39513;
  assign tmp42562 = l1 ? tmp40705 : tmp40823;
  assign tmp42561 = s0 ? tmp42547 : tmp42562;
  assign tmp42563 = s0 ? tmp40693 : tmp42547;
  assign tmp42560 = ~(s1 ? tmp42561 : tmp42563);
  assign tmp42558 = ~(s2 ? tmp42559 : tmp42560);
  assign tmp42549 = s3 ? tmp42550 : tmp42558;
  assign tmp42531 = s4 ? tmp42532 : tmp42549;
  assign tmp42570 = l1 ? tmp40729 : tmp40816;
  assign tmp42569 = s0 ? tmp42570 : tmp40096;
  assign tmp42571 = ~(l1 ? tmp39402 : tmp39518);
  assign tmp42568 = s1 ? tmp42569 : tmp42571;
  assign tmp42573 = l1 ? tmp40729 : tmp39430;
  assign tmp42574 = s0 ? tmp42562 : tmp39401;
  assign tmp42572 = s1 ? tmp42573 : tmp42574;
  assign tmp42567 = s2 ? tmp42568 : tmp42572;
  assign tmp42577 = ~(l1 ? tmp40705 : tmp40693);
  assign tmp42576 = s1 ? tmp42543 : tmp42577;
  assign tmp42579 = s0 ? tmp40693 : tmp42429;
  assign tmp42581 = l1 ? tmp40779 : tmp40861;
  assign tmp42580 = ~(s0 ? tmp42555 : tmp42581);
  assign tmp42578 = ~(s1 ? tmp42579 : tmp42580);
  assign tmp42575 = ~(s2 ? tmp42576 : tmp42578);
  assign tmp42566 = s3 ? tmp42567 : tmp42575;
  assign tmp42586 = l1 ? tmp40737 : tmp39430;
  assign tmp42585 = s0 ? tmp42435 : tmp42586;
  assign tmp42584 = s1 ? tmp42585 : tmp41898;
  assign tmp42583 = s2 ? tmp42584 : tmp42571;
  assign tmp42590 = ~(l1 ? tmp42173 : tmp39430);
  assign tmp42589 = s0 ? tmp39660 : tmp42590;
  assign tmp42588 = s1 ? tmp42589 : tmp42577;
  assign tmp42587 = ~(s2 ? tmp42588 : tmp42442);
  assign tmp42582 = s3 ? tmp42583 : tmp42587;
  assign tmp42565 = s4 ? tmp42566 : tmp42582;
  assign tmp42596 = l1 ? tmp40705 : tmp40693;
  assign tmp42595 = s0 ? tmp42596 : tmp42078;
  assign tmp42597 = ~(l1 ? tmp39513 : tmp39402);
  assign tmp42594 = s1 ? tmp42595 : tmp42597;
  assign tmp42599 = l1 ? tmp39630 : 1;
  assign tmp42600 = ~(l1 ? 1 : tmp39480);
  assign tmp42598 = s1 ? tmp42599 : tmp42600;
  assign tmp42593 = s2 ? tmp42594 : tmp42598;
  assign tmp42602 = ~(s1 ? tmp42453 : tmp42600);
  assign tmp42601 = ~(s2 ? tmp41635 : tmp42602);
  assign tmp42592 = s3 ? tmp42593 : tmp42601;
  assign tmp42605 = s1 ? tmp42457 : tmp40693;
  assign tmp42606 = ~(l1 ? tmp39513 : tmp39518);
  assign tmp42604 = s2 ? tmp42605 : tmp42606;
  assign tmp42608 = ~(l1 ? tmp39513 : tmp39459);
  assign tmp42607 = s1 ? tmp42526 : tmp42608;
  assign tmp42603 = s3 ? tmp42604 : tmp42607;
  assign tmp42591 = s4 ? tmp42592 : tmp42603;
  assign tmp42564 = s5 ? tmp42565 : tmp42591;
  assign tmp42530 = s6 ? tmp42531 : tmp42564;
  assign tmp42529 = s7 ? tmp39370 : tmp42530;
  assign tmp42528 = s8 ? tmp42462 : tmp42529;
  assign tmp42380 = s9 ? tmp42381 : tmp42528;
  assign tmp42616 = l1 ? tmp42268 : tmp40729;
  assign tmp42618 = ~(l2 ? tmp39430 : tmp40634);
  assign tmp42617 = ~(s0 ? tmp41847 : tmp42618);
  assign tmp42615 = s1 ? tmp42616 : tmp42617;
  assign tmp42621 = s0 ? tmp41847 : tmp40743;
  assign tmp42623 = l1 ? tmp40779 : tmp39404;
  assign tmp42622 = s0 ? tmp42623 : tmp40743;
  assign tmp42620 = s1 ? tmp42621 : tmp42622;
  assign tmp42625 = s0 ? tmp42623 : tmp39420;
  assign tmp42627 = ~(l1 ? tmp40779 : tmp40743);
  assign tmp42626 = ~(s0 ? tmp40737 : tmp42627);
  assign tmp42624 = s1 ? tmp42625 : tmp42626;
  assign tmp42619 = ~(s2 ? tmp42620 : tmp42624);
  assign tmp42614 = s3 ? tmp42615 : tmp42619;
  assign tmp42632 = l1 ? tmp39587 : tmp40729;
  assign tmp42631 = s0 ? tmp42632 : tmp40024;
  assign tmp42634 = l1 ? tmp40779 : tmp40743;
  assign tmp42633 = ~(s0 ? tmp42634 : tmp40743);
  assign tmp42630 = s1 ? tmp42631 : tmp42633;
  assign tmp42636 = s0 ? tmp42616 : tmp40225;
  assign tmp42635 = s1 ? tmp42636 : tmp41869;
  assign tmp42629 = s2 ? tmp42630 : tmp42635;
  assign tmp42640 = l1 ? tmp40705 : tmp40737;
  assign tmp42639 = s0 ? tmp40737 : tmp42640;
  assign tmp42641 = s0 ? tmp40693 : tmp40737;
  assign tmp42638 = ~(s1 ? tmp42639 : tmp42641);
  assign tmp42637 = ~(s2 ? tmp42559 : tmp42638);
  assign tmp42628 = s3 ? tmp42629 : tmp42637;
  assign tmp42613 = s4 ? tmp42614 : tmp42628;
  assign tmp42647 = s0 ? tmp40729 : tmp40096;
  assign tmp42646 = s1 ? tmp42647 : tmp39401;
  assign tmp42649 = l1 ? tmp40729 : tmp40771;
  assign tmp42650 = s0 ? tmp42640 : tmp39401;
  assign tmp42648 = s1 ? tmp42649 : tmp42650;
  assign tmp42645 = s2 ? tmp42646 : tmp42648;
  assign tmp42652 = s1 ? tmp42623 : tmp42441;
  assign tmp42654 = ~(s0 ? tmp42634 : tmp40779);
  assign tmp42653 = ~(s1 ? tmp42579 : tmp42654);
  assign tmp42651 = ~(s2 ? tmp42652 : tmp42653);
  assign tmp42644 = s3 ? tmp42645 : tmp42651;
  assign tmp42659 = l1 ? tmp40737 : tmp40771;
  assign tmp42658 = s0 ? tmp42435 : tmp42659;
  assign tmp42657 = s1 ? tmp42658 : tmp41898;
  assign tmp42656 = s2 ? tmp42657 : tmp39401;
  assign tmp42663 = l1 ? 1 : tmp39404;
  assign tmp42664 = ~(l1 ? tmp42173 : tmp40771);
  assign tmp42662 = s0 ? tmp42663 : tmp42664;
  assign tmp42661 = s1 ? tmp42662 : tmp42441;
  assign tmp42660 = ~(s2 ? tmp42661 : tmp42442);
  assign tmp42655 = s3 ? tmp42656 : tmp42660;
  assign tmp42643 = s4 ? tmp42644 : tmp42655;
  assign tmp42669 = s0 ? tmp40705 : tmp42078;
  assign tmp42668 = s1 ? tmp42669 : tmp42597;
  assign tmp42671 = l1 ? tmp39630 : tmp39480;
  assign tmp42670 = s1 ? tmp42671 : 0;
  assign tmp42667 = s2 ? tmp42668 : tmp42670;
  assign tmp42666 = s3 ? tmp42667 : tmp42451;
  assign tmp42674 = ~(l1 ? tmp39513 : tmp39404);
  assign tmp42673 = s2 ? tmp42605 : tmp42674;
  assign tmp42672 = s3 ? tmp42673 : tmp42525;
  assign tmp42665 = s4 ? tmp42666 : tmp42672;
  assign tmp42642 = s5 ? tmp42643 : tmp42665;
  assign tmp42612 = s6 ? tmp42613 : tmp42642;
  assign tmp42611 = s7 ? tmp39370 : tmp42612;
  assign tmp42610 = s8 ? tmp42611 : tmp39370;
  assign tmp42679 = s4 ? tmp42444 : tmp42524;
  assign tmp42678 = s5 ? tmp42416 : tmp42679;
  assign tmp42677 = s6 ? tmp42384 : tmp42678;
  assign tmp42676 = s7 ? tmp42677 : tmp42530;
  assign tmp42680 = s7 ? tmp42463 : tmp42612;
  assign tmp42675 = s8 ? tmp42676 : tmp42680;
  assign tmp42609 = s9 ? tmp42610 : tmp42675;
  assign tmp42379 = s10 ? tmp42380 : tmp42609;
  assign tmp42684 = s7 ? tmp42383 : tmp42530;
  assign tmp42683 = s8 ? tmp42684 : tmp42680;
  assign tmp42682 = s9 ? tmp42610 : tmp42683;
  assign tmp42681 = s10 ? tmp42380 : tmp42682;
  assign tmp42378 = s11 ? tmp42379 : tmp42681;
  assign tmp42103 = s12 ? tmp42104 : tmp42378;
  assign tmp42695 = l2 ? 1 : tmp39616;
  assign tmp42694 = l1 ? tmp40419 : tmp42695;
  assign tmp42697 = ~(l1 ? tmp39397 : tmp39385);
  assign tmp42696 = ~(s0 ? tmp39422 : tmp42697);
  assign tmp42693 = s1 ? tmp42694 : tmp42696;
  assign tmp42701 = ~(l1 ? tmp40419 : tmp40632);
  assign tmp42700 = s0 ? tmp41570 : tmp42701;
  assign tmp42702 = s0 ? tmp39414 : tmp42701;
  assign tmp42699 = s1 ? tmp42700 : tmp42702;
  assign tmp42705 = l1 ? tmp40419 : tmp40632;
  assign tmp42707 = l2 ? tmp39376 : tmp39430;
  assign tmp42708 = ~(l2 ? tmp39378 : tmp39616);
  assign tmp42706 = ~(l1 ? tmp42707 : tmp42708);
  assign tmp42704 = ~(s0 ? tmp42705 : tmp42706);
  assign tmp42703 = s1 ? tmp39446 : tmp42704;
  assign tmp42698 = ~(s2 ? tmp42699 : tmp42703);
  assign tmp42692 = s3 ? tmp42693 : tmp42698;
  assign tmp42712 = s0 ? tmp39383 : tmp40024;
  assign tmp42714 = l1 ? tmp42707 : tmp42708;
  assign tmp42713 = ~(s0 ? tmp42714 : tmp42701);
  assign tmp42711 = s1 ? tmp42712 : tmp42713;
  assign tmp42716 = s0 ? tmp42694 : tmp40225;
  assign tmp42715 = s1 ? tmp42716 : tmp41587;
  assign tmp42710 = s2 ? tmp42711 : tmp42715;
  assign tmp42719 = l1 ? tmp39435 : tmp39430;
  assign tmp42718 = s1 ? tmp39422 : tmp42719;
  assign tmp42722 = l1 ? tmp39915 : tmp40632;
  assign tmp42721 = s0 ? tmp42705 : tmp42722;
  assign tmp42723 = s0 ? tmp39378 : tmp42705;
  assign tmp42720 = ~(s1 ? tmp42721 : tmp42723);
  assign tmp42717 = ~(s2 ? tmp42718 : tmp42720);
  assign tmp42709 = s3 ? tmp42710 : tmp42717;
  assign tmp42691 = s4 ? tmp42692 : tmp42709;
  assign tmp42729 = s0 ? tmp39396 : tmp40096;
  assign tmp42728 = s1 ? tmp42729 : tmp41603;
  assign tmp42731 = l1 ? tmp39397 : 1;
  assign tmp42732 = s0 ? tmp42722 : tmp39401;
  assign tmp42730 = s1 ? tmp42731 : tmp42732;
  assign tmp42727 = s2 ? tmp42728 : tmp42730;
  assign tmp42735 = ~(l1 ? tmp39915 : tmp39378);
  assign tmp42734 = s1 ? tmp39414 : tmp42735;
  assign tmp42738 = l1 ? tmp42707 : tmp39376;
  assign tmp42737 = ~(s0 ? tmp42714 : tmp42738);
  assign tmp42736 = ~(s1 ? tmp39378 : tmp42737);
  assign tmp42733 = ~(s2 ? tmp42734 : tmp42736);
  assign tmp42726 = s3 ? tmp42727 : tmp42733;
  assign tmp42743 = l1 ? tmp40419 : tmp39513;
  assign tmp42742 = s0 ? tmp39378 : tmp42743;
  assign tmp42741 = s1 ? tmp42742 : tmp41620;
  assign tmp42744 = ~(l1 ? tmp39375 : tmp42708);
  assign tmp42740 = s2 ? tmp42741 : tmp42744;
  assign tmp42748 = l1 ? tmp39429 : tmp42708;
  assign tmp42749 = ~(l1 ? tmp39915 : tmp39513);
  assign tmp42747 = s0 ? tmp42748 : tmp42749;
  assign tmp42746 = s1 ? tmp42747 : tmp42735;
  assign tmp42750 = s1 ? 1 : tmp42719;
  assign tmp42745 = ~(s2 ? tmp42746 : tmp42750);
  assign tmp42739 = s3 ? tmp42740 : tmp42745;
  assign tmp42725 = s4 ? tmp42726 : tmp42739;
  assign tmp42756 = l1 ? tmp39915 : tmp39378;
  assign tmp42755 = s0 ? tmp42756 : 0;
  assign tmp42754 = s1 ? tmp42755 : tmp39658;
  assign tmp42753 = s2 ? tmp42754 : tmp40275;
  assign tmp42760 = ~(l1 ? tmp39513 : tmp39378);
  assign tmp42759 = s0 ? tmp39526 : tmp42760;
  assign tmp42758 = s1 ? tmp39435 : tmp42759;
  assign tmp42762 = l1 ? tmp39378 : tmp39513;
  assign tmp42763 = ~(l1 ? tmp39429 : tmp40771);
  assign tmp42761 = ~(s1 ? tmp42762 : tmp42763);
  assign tmp42757 = ~(s2 ? tmp42758 : tmp42761);
  assign tmp42752 = s3 ? tmp42753 : tmp42757;
  assign tmp42766 = s1 ? tmp39512 : tmp39378;
  assign tmp42767 = ~(l1 ? tmp39430 : tmp42708);
  assign tmp42765 = s2 ? tmp42766 : tmp42767;
  assign tmp42770 = l1 ? tmp39513 : tmp39378;
  assign tmp42771 = ~(l1 ? tmp39430 : tmp40771);
  assign tmp42769 = s1 ? tmp42770 : tmp42771;
  assign tmp42772 = ~(l1 ? tmp39435 : tmp39527);
  assign tmp42768 = s2 ? tmp42769 : tmp42772;
  assign tmp42764 = s3 ? tmp42765 : tmp42768;
  assign tmp42751 = s4 ? tmp42752 : tmp42764;
  assign tmp42724 = s5 ? tmp42725 : tmp42751;
  assign tmp42690 = s6 ? tmp42691 : tmp42724;
  assign tmp42689 = s7 ? tmp39370 : tmp42690;
  assign tmp42779 = l1 ? tmp40419 : tmp39397;
  assign tmp42781 = ~(l1 ? tmp39397 : tmp39384);
  assign tmp42780 = ~(s0 ? tmp39422 : tmp42781);
  assign tmp42778 = s1 ? tmp42779 : tmp42780;
  assign tmp42785 = ~(l2 ? tmp39378 : tmp39398);
  assign tmp42784 = s0 ? tmp41570 : tmp42785;
  assign tmp42786 = s0 ? tmp39414 : tmp42785;
  assign tmp42783 = s1 ? tmp42784 : tmp42786;
  assign tmp42789 = ~(l1 ? tmp42707 : tmp42785);
  assign tmp42788 = ~(s0 ? tmp40419 : tmp42789);
  assign tmp42787 = s1 ? tmp39446 : tmp42788;
  assign tmp42782 = ~(s2 ? tmp42783 : tmp42787);
  assign tmp42777 = s3 ? tmp42778 : tmp42782;
  assign tmp42793 = s0 ? tmp39384 : tmp40024;
  assign tmp42795 = l1 ? tmp42707 : tmp42785;
  assign tmp42794 = ~(s0 ? tmp42795 : tmp42785);
  assign tmp42792 = s1 ? tmp42793 : tmp42794;
  assign tmp42797 = s0 ? tmp42779 : tmp40225;
  assign tmp42796 = s1 ? tmp42797 : tmp41587;
  assign tmp42791 = s2 ? tmp42792 : tmp42796;
  assign tmp42801 = l1 ? tmp39915 : tmp40419;
  assign tmp42800 = s0 ? tmp40419 : tmp42801;
  assign tmp42802 = s0 ? tmp39378 : tmp40419;
  assign tmp42799 = ~(s1 ? tmp42800 : tmp42802);
  assign tmp42798 = ~(s2 ? tmp42718 : tmp42799);
  assign tmp42790 = s3 ? tmp42791 : tmp42798;
  assign tmp42776 = s4 ? tmp42777 : tmp42790;
  assign tmp42809 = l1 ? tmp39397 : tmp39384;
  assign tmp42808 = s0 ? tmp42809 : tmp40096;
  assign tmp42807 = s1 ? tmp42808 : tmp41603;
  assign tmp42811 = l1 ? tmp39397 : tmp39480;
  assign tmp42812 = s0 ? tmp42801 : tmp39401;
  assign tmp42810 = s1 ? tmp42811 : tmp42812;
  assign tmp42806 = s2 ? tmp42807 : tmp42810;
  assign tmp42815 = ~(l2 ? tmp39378 : tmp39460);
  assign tmp42814 = s1 ? tmp39414 : tmp42815;
  assign tmp42817 = ~(s0 ? tmp42795 : tmp42707);
  assign tmp42816 = ~(s1 ? tmp39378 : tmp42817);
  assign tmp42813 = ~(s2 ? tmp42814 : tmp42816);
  assign tmp42805 = s3 ? tmp42806 : tmp42813;
  assign tmp42822 = l1 ? tmp40419 : tmp39459;
  assign tmp42821 = s0 ? tmp39378 : tmp42822;
  assign tmp42820 = s1 ? tmp42821 : tmp41620;
  assign tmp42823 = ~(l1 ? tmp39375 : tmp42785);
  assign tmp42819 = s2 ? tmp42820 : tmp42823;
  assign tmp42827 = l1 ? tmp39429 : tmp42785;
  assign tmp42828 = ~(l1 ? tmp39915 : tmp39459);
  assign tmp42826 = s0 ? tmp42827 : tmp42828;
  assign tmp42825 = s1 ? tmp42826 : tmp42815;
  assign tmp42824 = ~(s2 ? tmp42825 : tmp42750);
  assign tmp42818 = s3 ? tmp42819 : tmp42824;
  assign tmp42804 = s4 ? tmp42805 : tmp42818;
  assign tmp42833 = s0 ? tmp39915 : 0;
  assign tmp42832 = s1 ? tmp42833 : tmp39658;
  assign tmp42831 = s2 ? tmp42832 : tmp40275;
  assign tmp42836 = ~(l1 ? tmp39429 : tmp39430);
  assign tmp42835 = ~(s1 ? tmp42762 : tmp42836);
  assign tmp42834 = ~(s2 ? tmp42758 : tmp42835);
  assign tmp42830 = s3 ? tmp42831 : tmp42834;
  assign tmp42839 = ~(l1 ? tmp39430 : tmp42785);
  assign tmp42838 = s2 ? tmp42766 : tmp42839;
  assign tmp42841 = s1 ? tmp42770 : tmp39398;
  assign tmp42840 = s2 ? tmp42841 : tmp42772;
  assign tmp42837 = s3 ? tmp42838 : tmp42840;
  assign tmp42829 = s4 ? tmp42830 : tmp42837;
  assign tmp42803 = s5 ? tmp42804 : tmp42829;
  assign tmp42775 = s6 ? tmp42776 : tmp42803;
  assign tmp42774 = s7 ? tmp39370 : tmp42775;
  assign tmp42773 = s8 ? tmp42689 : tmp42774;
  assign tmp42688 = s9 ? tmp42689 : tmp42773;
  assign tmp42843 = s8 ? tmp42689 : tmp39370;
  assign tmp42849 = s3 ? tmp42765 : tmp42769;
  assign tmp42848 = s4 ? tmp42752 : tmp42849;
  assign tmp42847 = s5 ? tmp42725 : tmp42848;
  assign tmp42846 = s6 ? tmp42691 : tmp42847;
  assign tmp42853 = s3 ? tmp42838 : tmp42841;
  assign tmp42852 = s4 ? tmp42830 : tmp42853;
  assign tmp42851 = s5 ? tmp42804 : tmp42852;
  assign tmp42850 = s6 ? tmp42776 : tmp42851;
  assign tmp42845 = s7 ? tmp42846 : tmp42850;
  assign tmp42844 = s8 ? tmp42845 : tmp42846;
  assign tmp42842 = s9 ? tmp42843 : tmp42844;
  assign tmp42687 = s10 ? tmp42688 : tmp42842;
  assign tmp42857 = s7 ? tmp42690 : tmp42775;
  assign tmp42856 = s8 ? tmp42857 : tmp42690;
  assign tmp42855 = s9 ? tmp42843 : tmp42856;
  assign tmp42854 = s10 ? tmp42688 : tmp42855;
  assign tmp42686 = s11 ? tmp42687 : tmp42854;
  assign tmp42867 = l1 ? tmp42119 : tmp39384;
  assign tmp42869 = l1 ? 1 : tmp39423;
  assign tmp42870 = ~(l1 ? tmp39575 : tmp39384);
  assign tmp42868 = ~(s0 ? tmp42869 : tmp42870);
  assign tmp42866 = s1 ? tmp42867 : tmp42868;
  assign tmp42874 = ~(l1 ? tmp42119 : tmp42017);
  assign tmp42873 = s0 ? tmp39786 : tmp42874;
  assign tmp42876 = l1 ? tmp39513 : tmp39423;
  assign tmp42875 = s0 ? tmp42876 : tmp42874;
  assign tmp42872 = s1 ? tmp42873 : tmp42875;
  assign tmp42878 = s0 ? tmp42876 : tmp39420;
  assign tmp42880 = l1 ? tmp42119 : tmp42017;
  assign tmp42882 = ~(l2 ? tmp39378 : tmp39381);
  assign tmp42881 = ~(l1 ? tmp39527 : tmp42882);
  assign tmp42879 = ~(s0 ? tmp42880 : tmp42881);
  assign tmp42877 = s1 ? tmp42878 : tmp42879;
  assign tmp42871 = ~(s2 ? tmp42872 : tmp42877);
  assign tmp42865 = s3 ? tmp42866 : tmp42871;
  assign tmp42887 = l1 ? tmp39575 : tmp39384;
  assign tmp42886 = s0 ? tmp42887 : tmp40024;
  assign tmp42889 = l1 ? tmp39527 : tmp42882;
  assign tmp42888 = ~(s0 ? tmp42889 : tmp42874);
  assign tmp42885 = s1 ? tmp42886 : tmp42888;
  assign tmp42891 = s0 ? tmp42867 : tmp40225;
  assign tmp42890 = s1 ? tmp42891 : tmp41587;
  assign tmp42884 = s2 ? tmp42885 : tmp42890;
  assign tmp42894 = l1 ? tmp39527 : tmp40982;
  assign tmp42893 = s1 ? tmp39422 : tmp42894;
  assign tmp42897 = l1 ? tmp42155 : tmp42017;
  assign tmp42896 = s0 ? tmp42880 : tmp42897;
  assign tmp42899 = l1 ? tmp41738 : tmp39501;
  assign tmp42898 = s0 ? tmp42899 : tmp42880;
  assign tmp42895 = ~(s1 ? tmp42896 : tmp42898);
  assign tmp42892 = ~(s2 ? tmp42893 : tmp42895);
  assign tmp42883 = s3 ? tmp42884 : tmp42892;
  assign tmp42864 = s4 ? tmp42865 : tmp42883;
  assign tmp42905 = s0 ? tmp42887 : tmp40096;
  assign tmp42904 = s1 ? tmp42905 : tmp40096;
  assign tmp42907 = l1 ? tmp39575 : tmp39480;
  assign tmp42908 = s0 ? tmp42897 : tmp39401;
  assign tmp42906 = s1 ? tmp42907 : tmp42908;
  assign tmp42903 = s2 ? tmp42904 : tmp42906;
  assign tmp42911 = ~(l1 ? tmp42173 : tmp42043);
  assign tmp42910 = s1 ? tmp42876 : tmp42911;
  assign tmp42913 = s0 ? tmp42899 : tmp39501;
  assign tmp42915 = l1 ? tmp39527 : tmp42029;
  assign tmp42914 = ~(s0 ? tmp42889 : tmp42915);
  assign tmp42912 = ~(s1 ? tmp42913 : tmp42914);
  assign tmp42909 = ~(s2 ? tmp42910 : tmp42912);
  assign tmp42902 = s3 ? tmp42903 : tmp42909;
  assign tmp42920 = l1 ? tmp42119 : tmp39480;
  assign tmp42919 = s0 ? tmp39501 : tmp42920;
  assign tmp42918 = s1 ? tmp42919 : tmp41620;
  assign tmp42921 = ~(l1 ? 1 : tmp42785);
  assign tmp42917 = s2 ? tmp42918 : tmp42921;
  assign tmp42925 = l1 ? 1 : tmp42785;
  assign tmp42926 = ~(l1 ? tmp42155 : tmp39480);
  assign tmp42924 = s0 ? tmp42925 : tmp42926;
  assign tmp42923 = s1 ? tmp42924 : tmp42911;
  assign tmp42927 = s1 ? tmp39651 : tmp42894;
  assign tmp42922 = ~(s2 ? tmp42923 : tmp42927);
  assign tmp42916 = s3 ? tmp42917 : tmp42922;
  assign tmp42901 = s4 ? tmp42902 : tmp42916;
  assign tmp42933 = l1 ? tmp42173 : tmp42043;
  assign tmp42932 = s0 ? tmp42933 : tmp42078;
  assign tmp42934 = ~(l1 ? tmp39513 : tmp39375);
  assign tmp42931 = s1 ? tmp42932 : tmp42934;
  assign tmp42930 = s2 ? tmp42931 : tmp42670;
  assign tmp42937 = ~(l1 ? 1 : tmp39501);
  assign tmp42936 = s1 ? tmp39526 : tmp42937;
  assign tmp42939 = ~(l1 ? 1 : tmp39430);
  assign tmp42938 = ~(s1 ? tmp39500 : tmp42939);
  assign tmp42935 = ~(s2 ? tmp42936 : tmp42938);
  assign tmp42929 = s3 ? tmp42930 : tmp42935;
  assign tmp42943 = s0 ? tmp39543 : tmp42899;
  assign tmp42942 = s1 ? tmp39549 : tmp42943;
  assign tmp42944 = ~(l1 ? tmp39527 : tmp42785);
  assign tmp42941 = s2 ? tmp42942 : tmp42944;
  assign tmp42947 = l1 ? tmp39429 : tmp39501;
  assign tmp42948 = ~(l1 ? tmp39527 : tmp40982);
  assign tmp42946 = s1 ? tmp42947 : tmp42948;
  assign tmp42945 = s2 ? tmp42946 : tmp39543;
  assign tmp42940 = s3 ? tmp42941 : tmp42945;
  assign tmp42928 = s4 ? tmp42929 : tmp42940;
  assign tmp42900 = s5 ? tmp42901 : tmp42928;
  assign tmp42863 = s6 ? tmp42864 : tmp42900;
  assign tmp42862 = s7 ? tmp39370 : tmp42863;
  assign tmp42954 = l1 ? tmp42268 : tmp39758;
  assign tmp42956 = l1 ? tmp39402 : tmp41327;
  assign tmp42957 = ~(l1 ? tmp39587 : tmp39758);
  assign tmp42955 = ~(s0 ? tmp42956 : tmp42957);
  assign tmp42953 = s1 ? tmp42954 : tmp42955;
  assign tmp42962 = l2 ? tmp39460 : tmp39381;
  assign tmp42961 = ~(l1 ? tmp42268 : tmp42962);
  assign tmp42960 = s0 ? tmp39477 : tmp42961;
  assign tmp42964 = l1 ? tmp40779 : tmp41327;
  assign tmp42963 = s0 ? tmp42964 : tmp42961;
  assign tmp42959 = s1 ? tmp42960 : tmp42963;
  assign tmp42966 = s0 ? tmp42964 : tmp41336;
  assign tmp42968 = l1 ? tmp42268 : tmp42962;
  assign tmp42970 = ~(l2 ? tmp39460 : tmp39381);
  assign tmp42969 = ~(l1 ? tmp39684 : tmp42970);
  assign tmp42967 = ~(s0 ? tmp42968 : tmp42969);
  assign tmp42965 = s1 ? tmp42966 : tmp42967;
  assign tmp42958 = ~(s2 ? tmp42959 : tmp42965);
  assign tmp42952 = s3 ? tmp42953 : tmp42958;
  assign tmp42975 = l1 ? tmp39587 : tmp39758;
  assign tmp42974 = s0 ? tmp42975 : tmp40024;
  assign tmp42977 = l1 ? tmp39684 : tmp42970;
  assign tmp42976 = ~(s0 ? tmp42977 : tmp42961);
  assign tmp42973 = s1 ? tmp42974 : tmp42976;
  assign tmp42979 = s0 ? tmp42954 : tmp40225;
  assign tmp42980 = l1 ? tmp39384 : tmp39402;
  assign tmp42978 = s1 ? tmp42979 : tmp42980;
  assign tmp42972 = s2 ? tmp42973 : tmp42978;
  assign tmp42982 = s1 ? tmp42956 : tmp42894;
  assign tmp42985 = l1 ? tmp42173 : tmp42962;
  assign tmp42984 = s0 ? tmp42968 : tmp42985;
  assign tmp42988 = l2 ? tmp39460 : 1;
  assign tmp42987 = l1 ? tmp41738 : tmp42988;
  assign tmp42986 = s0 ? tmp42987 : tmp42968;
  assign tmp42983 = ~(s1 ? tmp42984 : tmp42986);
  assign tmp42981 = ~(s2 ? tmp42982 : tmp42983);
  assign tmp42971 = s3 ? tmp42972 : tmp42981;
  assign tmp42951 = s4 ? tmp42952 : tmp42971;
  assign tmp42994 = s0 ? tmp42975 : tmp40096;
  assign tmp42993 = s1 ? tmp42994 : tmp40024;
  assign tmp42996 = l1 ? tmp39587 : tmp39403;
  assign tmp42997 = s0 ? tmp42985 : tmp40024;
  assign tmp42995 = s1 ? tmp42996 : tmp42997;
  assign tmp42992 = s2 ? tmp42993 : tmp42995;
  assign tmp43001 = l2 ? tmp39460 : tmp39403;
  assign tmp43000 = ~(l1 ? tmp42173 : tmp43001);
  assign tmp42999 = s1 ? tmp42964 : tmp43000;
  assign tmp43003 = s0 ? tmp42987 : tmp39501;
  assign tmp43005 = l1 ? tmp39684 : tmp40982;
  assign tmp43004 = ~(s0 ? tmp42977 : tmp43005);
  assign tmp43002 = ~(s1 ? tmp43003 : tmp43004);
  assign tmp42998 = ~(s2 ? tmp42999 : tmp43002);
  assign tmp42991 = s3 ? tmp42992 : tmp42998;
  assign tmp43010 = l1 ? tmp42268 : tmp39403;
  assign tmp43009 = s0 ? tmp39501 : tmp43010;
  assign tmp43011 = s0 ? tmp41587 : tmp40527;
  assign tmp43008 = s1 ? tmp43009 : tmp43011;
  assign tmp43013 = ~(l2 ? tmp39460 : tmp39398);
  assign tmp43012 = ~(l1 ? tmp39402 : tmp43013);
  assign tmp43007 = s2 ? tmp43008 : tmp43012;
  assign tmp43017 = l1 ? 1 : tmp43013;
  assign tmp43018 = ~(l1 ? tmp42173 : tmp39403);
  assign tmp43016 = s0 ? tmp43017 : tmp43018;
  assign tmp43015 = s1 ? tmp43016 : tmp42911;
  assign tmp43014 = ~(s2 ? tmp43015 : tmp42927);
  assign tmp43006 = s3 ? tmp43007 : tmp43014;
  assign tmp42990 = s4 ? tmp42991 : tmp43006;
  assign tmp43024 = l1 ? tmp42173 : tmp43001;
  assign tmp43023 = s0 ? tmp43024 : tmp42078;
  assign tmp43025 = ~(l1 ? tmp39513 : tmp39429);
  assign tmp43022 = s1 ? tmp43023 : tmp43025;
  assign tmp43021 = s2 ? tmp43022 : tmp42522;
  assign tmp43020 = s3 ? tmp43021 : tmp42935;
  assign tmp43029 = s0 ? tmp39543 : tmp42987;
  assign tmp43028 = s1 ? tmp39549 : tmp43029;
  assign tmp43030 = ~(l1 ? tmp39527 : tmp43013);
  assign tmp43027 = s2 ? tmp43028 : tmp43030;
  assign tmp43026 = s3 ? tmp43027 : tmp42945;
  assign tmp43019 = s4 ? tmp43020 : tmp43026;
  assign tmp42989 = s5 ? tmp42990 : tmp43019;
  assign tmp42950 = s6 ? tmp42951 : tmp42989;
  assign tmp42949 = s7 ? tmp39370 : tmp42950;
  assign tmp42861 = s8 ? tmp42862 : tmp42949;
  assign tmp43037 = l1 ? tmp42268 : tmp39384;
  assign tmp43039 = ~(l1 ? tmp39587 : tmp39384);
  assign tmp43038 = ~(s0 ? tmp39422 : tmp43039);
  assign tmp43036 = s1 ? tmp43037 : tmp43038;
  assign tmp43043 = ~(l1 ? tmp42268 : tmp42017);
  assign tmp43042 = s0 ? tmp42540 : tmp43043;
  assign tmp43045 = l1 ? tmp40779 : tmp39388;
  assign tmp43044 = s0 ? tmp43045 : tmp43043;
  assign tmp43041 = s1 ? tmp43042 : tmp43044;
  assign tmp43047 = s0 ? tmp43045 : tmp39420;
  assign tmp43049 = l1 ? tmp42268 : tmp42017;
  assign tmp43050 = ~(l1 ? tmp39684 : tmp42882);
  assign tmp43048 = ~(s0 ? tmp43049 : tmp43050);
  assign tmp43046 = s1 ? tmp43047 : tmp43048;
  assign tmp43040 = ~(s2 ? tmp43041 : tmp43046);
  assign tmp43035 = s3 ? tmp43036 : tmp43040;
  assign tmp43055 = l1 ? tmp39587 : tmp39384;
  assign tmp43054 = s0 ? tmp43055 : tmp40024;
  assign tmp43057 = l1 ? tmp39684 : tmp42882;
  assign tmp43056 = ~(s0 ? tmp43057 : tmp43043);
  assign tmp43053 = s1 ? tmp43054 : tmp43056;
  assign tmp43059 = s0 ? tmp43037 : tmp40225;
  assign tmp43058 = s1 ? tmp43059 : tmp41587;
  assign tmp43052 = s2 ? tmp43053 : tmp43058;
  assign tmp43063 = l1 ? tmp42173 : tmp42017;
  assign tmp43062 = s0 ? tmp43049 : tmp43063;
  assign tmp43064 = s0 ? tmp42899 : tmp43049;
  assign tmp43061 = ~(s1 ? tmp43062 : tmp43064);
  assign tmp43060 = ~(s2 ? tmp42893 : tmp43061);
  assign tmp43051 = s3 ? tmp43052 : tmp43060;
  assign tmp43034 = s4 ? tmp43035 : tmp43051;
  assign tmp43070 = s0 ? tmp43055 : tmp40096;
  assign tmp43069 = s1 ? tmp43070 : tmp42571;
  assign tmp43072 = l1 ? tmp39587 : tmp39480;
  assign tmp43073 = s0 ? tmp43063 : tmp39401;
  assign tmp43071 = s1 ? tmp43072 : tmp43073;
  assign tmp43068 = s2 ? tmp43069 : tmp43071;
  assign tmp43075 = s1 ? tmp43045 : tmp42911;
  assign tmp43078 = l1 ? tmp39684 : tmp42029;
  assign tmp43077 = ~(s0 ? tmp43057 : tmp43078);
  assign tmp43076 = ~(s1 ? tmp42913 : tmp43077);
  assign tmp43074 = ~(s2 ? tmp43075 : tmp43076);
  assign tmp43067 = s3 ? tmp43068 : tmp43074;
  assign tmp43083 = l1 ? tmp42268 : tmp39480;
  assign tmp43082 = s0 ? tmp39501 : tmp43083;
  assign tmp43081 = s1 ? tmp43082 : tmp41620;
  assign tmp43084 = ~(l1 ? tmp39402 : tmp42785);
  assign tmp43080 = s2 ? tmp43081 : tmp43084;
  assign tmp43088 = ~(l1 ? tmp42173 : tmp39480);
  assign tmp43087 = s0 ? tmp42925 : tmp43088;
  assign tmp43086 = s1 ? tmp43087 : tmp42911;
  assign tmp43085 = ~(s2 ? tmp43086 : tmp42927);
  assign tmp43079 = s3 ? tmp43080 : tmp43085;
  assign tmp43066 = s4 ? tmp43067 : tmp43079;
  assign tmp43091 = s2 ? tmp42931 : tmp42598;
  assign tmp43090 = s3 ? tmp43091 : tmp42935;
  assign tmp43089 = s4 ? tmp43090 : tmp42940;
  assign tmp43065 = s5 ? tmp43066 : tmp43089;
  assign tmp43033 = s6 ? tmp43034 : tmp43065;
  assign tmp43032 = s7 ? tmp39370 : tmp43033;
  assign tmp43031 = s8 ? tmp42949 : tmp43032;
  assign tmp42860 = s9 ? tmp42861 : tmp43031;
  assign tmp43100 = s0 ? tmp41847 : tmp43043;
  assign tmp43102 = l1 ? tmp40779 : tmp39423;
  assign tmp43101 = s0 ? tmp43102 : tmp43043;
  assign tmp43099 = s1 ? tmp43100 : tmp43101;
  assign tmp43104 = s0 ? tmp43102 : tmp39420;
  assign tmp43103 = s1 ? tmp43104 : tmp43048;
  assign tmp43098 = ~(s2 ? tmp43099 : tmp43103);
  assign tmp43097 = s3 ? tmp43036 : tmp43098;
  assign tmp43096 = s4 ? tmp43097 : tmp43051;
  assign tmp43109 = s1 ? tmp43070 : tmp39401;
  assign tmp43108 = s2 ? tmp43109 : tmp43071;
  assign tmp43111 = s1 ? tmp43102 : tmp42911;
  assign tmp43110 = ~(s2 ? tmp43111 : tmp43076);
  assign tmp43107 = s3 ? tmp43108 : tmp43110;
  assign tmp43106 = s4 ? tmp43107 : tmp43079;
  assign tmp43105 = s5 ? tmp43106 : tmp42928;
  assign tmp43095 = s6 ? tmp43096 : tmp43105;
  assign tmp43094 = s7 ? tmp39370 : tmp43095;
  assign tmp43093 = s8 ? tmp43094 : tmp39370;
  assign tmp43117 = s3 ? tmp42941 : tmp42946;
  assign tmp43116 = s4 ? tmp42929 : tmp43117;
  assign tmp43115 = s5 ? tmp42901 : tmp43116;
  assign tmp43114 = s6 ? tmp42864 : tmp43115;
  assign tmp43120 = s4 ? tmp43090 : tmp43117;
  assign tmp43119 = s5 ? tmp43066 : tmp43120;
  assign tmp43118 = s6 ? tmp43034 : tmp43119;
  assign tmp43113 = s7 ? tmp43114 : tmp43118;
  assign tmp43125 = s3 ? tmp43027 : tmp42946;
  assign tmp43124 = s4 ? tmp43020 : tmp43125;
  assign tmp43123 = s5 ? tmp42990 : tmp43124;
  assign tmp43122 = s6 ? tmp42951 : tmp43123;
  assign tmp43127 = s5 ? tmp43106 : tmp43116;
  assign tmp43126 = s6 ? tmp43096 : tmp43127;
  assign tmp43121 = s7 ? tmp43122 : tmp43126;
  assign tmp43112 = s8 ? tmp43113 : tmp43121;
  assign tmp43092 = s9 ? tmp43093 : tmp43112;
  assign tmp42859 = s10 ? tmp42860 : tmp43092;
  assign tmp43131 = s7 ? tmp42863 : tmp43033;
  assign tmp43132 = s7 ? tmp42950 : tmp43095;
  assign tmp43130 = s8 ? tmp43131 : tmp43132;
  assign tmp43129 = s9 ? tmp43093 : tmp43130;
  assign tmp43128 = s10 ? tmp42860 : tmp43129;
  assign tmp42858 = s11 ? tmp42859 : tmp43128;
  assign tmp42685 = s12 ? tmp42686 : tmp42858;
  assign tmp42102 = s13 ? tmp42103 : tmp42685;
  assign tmp41554 = s14 ? tmp41555 : tmp42102;
  assign tmp39362 = s15 ? tmp39363 : tmp41554;
  assign tmp43147 = ~(s0 ? tmp39692 : tmp39487);
  assign tmp43146 = s1 ? tmp39483 : tmp43147;
  assign tmp43145 = s2 ? tmp39633 : tmp43146;
  assign tmp43144 = s3 ? tmp43145 : tmp39732;
  assign tmp43143 = s4 ? tmp39711 : tmp43144;
  assign tmp43142 = s5 ? tmp43143 : tmp39736;
  assign tmp43141 = s6 ? tmp39677 : tmp43142;
  assign tmp43140 = s7 ? tmp39370 : tmp43141;
  assign tmp43139 = s8 ? tmp39369 : tmp43140;
  assign tmp43138 = s9 ? tmp43139 : tmp43140;
  assign tmp43149 = s8 ? tmp43140 : tmp39370;
  assign tmp43156 = l1 ? tmp39681 : tmp39755;
  assign tmp43158 = ~(l1 ? tmp39684 : tmp39755);
  assign tmp43157 = ~(s0 ? tmp39569 : tmp43158);
  assign tmp43155 = s1 ? tmp43156 : tmp43157;
  assign tmp43162 = ~(l1 ? tmp39577 : tmp39765);
  assign tmp43161 = s0 ? tmp42996 : tmp43162;
  assign tmp43164 = l1 ? tmp39587 : tmp39621;
  assign tmp43163 = s0 ? tmp43164 : tmp43162;
  assign tmp43160 = s1 ? tmp43161 : tmp43163;
  assign tmp43166 = s0 ? tmp43164 : tmp39695;
  assign tmp43168 = l1 ? tmp39577 : tmp39765;
  assign tmp43169 = ~(l1 ? tmp39587 : tmp39493);
  assign tmp43167 = ~(s0 ? tmp43168 : tmp43169);
  assign tmp43165 = s1 ? tmp43166 : tmp43167;
  assign tmp43159 = ~(s2 ? tmp43160 : tmp43165);
  assign tmp43154 = s3 ? tmp43155 : tmp43159;
  assign tmp43174 = l1 ? tmp39402 : tmp39755;
  assign tmp43173 = s0 ? tmp43174 : tmp39594;
  assign tmp43176 = l1 ? tmp39587 : tmp39493;
  assign tmp43175 = ~(s0 ? tmp43176 : tmp43162);
  assign tmp43172 = s1 ? tmp43173 : tmp43175;
  assign tmp43178 = s0 ? tmp43156 : tmp39487;
  assign tmp43177 = s1 ? tmp43178 : tmp39477;
  assign tmp43171 = s2 ? tmp43172 : tmp43177;
  assign tmp43181 = s0 ? tmp39603 : tmp43168;
  assign tmp43180 = ~(s1 ? tmp43168 : tmp43181);
  assign tmp43179 = ~(s2 ? tmp39600 : tmp43180);
  assign tmp43170 = s3 ? tmp43171 : tmp43179;
  assign tmp43153 = s4 ? tmp43154 : tmp43170;
  assign tmp43188 = l1 ? tmp39684 : tmp39755;
  assign tmp43187 = s0 ? tmp43188 : tmp39487;
  assign tmp43189 = ~(l1 ? tmp39587 : tmp39403);
  assign tmp43186 = s1 ? tmp43187 : tmp43189;
  assign tmp43191 = l1 ? tmp39684 : tmp39801;
  assign tmp43192 = s0 ? tmp43168 : tmp39720;
  assign tmp43190 = s1 ? tmp43191 : tmp43192;
  assign tmp43185 = s2 ? tmp43186 : tmp43190;
  assign tmp43194 = s1 ? tmp39823 : tmp39806;
  assign tmp43197 = l1 ? tmp39630 : tmp39493;
  assign tmp43196 = ~(s0 ? tmp43176 : tmp43197);
  assign tmp43195 = ~(s1 ? tmp39625 : tmp43196);
  assign tmp43193 = ~(s2 ? tmp43194 : tmp43195);
  assign tmp43184 = s3 ? tmp43185 : tmp43193;
  assign tmp43202 = l1 ? tmp39577 : tmp39801;
  assign tmp43201 = s0 ? tmp39635 : tmp43202;
  assign tmp43200 = s1 ? tmp43201 : tmp39638;
  assign tmp43204 = ~(l1 ? tmp39587 : tmp39621);
  assign tmp43203 = s1 ? tmp39483 : tmp43204;
  assign tmp43199 = s2 ? tmp43200 : tmp43203;
  assign tmp43208 = ~(l1 ? tmp39681 : tmp39435);
  assign tmp43207 = s0 ? tmp39823 : tmp43208;
  assign tmp43206 = s1 ? tmp43207 : tmp39648;
  assign tmp43205 = ~(s2 ? tmp43206 : tmp39650);
  assign tmp43198 = s3 ? tmp43199 : tmp43205;
  assign tmp43183 = s4 ? tmp43184 : tmp43198;
  assign tmp43182 = s5 ? tmp43183 : tmp39825;
  assign tmp43152 = s6 ? tmp43153 : tmp43182;
  assign tmp43151 = s7 ? tmp39892 : tmp43152;
  assign tmp43214 = s1 ? tmp39483 : tmp39731;
  assign tmp43213 = s2 ? tmp39633 : tmp43214;
  assign tmp43212 = s3 ? tmp43213 : tmp39732;
  assign tmp43211 = s4 ? tmp39711 : tmp43212;
  assign tmp43210 = s5 ? tmp43211 : tmp39736;
  assign tmp43209 = s6 ? tmp39677 : tmp43210;
  assign tmp43150 = s8 ? tmp43151 : tmp43209;
  assign tmp43148 = s9 ? tmp43149 : tmp43150;
  assign tmp43137 = s10 ? tmp43138 : tmp43148;
  assign tmp43225 = ~(s0 ? tmp43164 : tmp39487);
  assign tmp43224 = s1 ? tmp39483 : tmp43225;
  assign tmp43223 = s2 ? tmp43200 : tmp43224;
  assign tmp43222 = s3 ? tmp43223 : tmp43205;
  assign tmp43221 = s4 ? tmp43184 : tmp43222;
  assign tmp43220 = s5 ? tmp43221 : tmp39825;
  assign tmp43219 = s6 ? tmp43153 : tmp43220;
  assign tmp43218 = s7 ? tmp39562 : tmp43219;
  assign tmp43217 = s8 ? tmp43218 : tmp43141;
  assign tmp43216 = s9 ? tmp43149 : tmp43217;
  assign tmp43215 = s10 ? tmp43138 : tmp43216;
  assign tmp43136 = s11 ? tmp43137 : tmp43215;
  assign tmp43237 = s0 ? tmp40309 : tmp39424;
  assign tmp43236 = s1 ? tmp40308 : tmp43237;
  assign tmp43235 = s2 ? tmp40302 : tmp43236;
  assign tmp43239 = s1 ? tmp40286 : tmp39949;
  assign tmp43238 = ~(s2 ? tmp43239 : tmp40312);
  assign tmp43234 = s3 ? tmp43235 : tmp43238;
  assign tmp43233 = s4 ? tmp40282 : tmp43234;
  assign tmp43232 = s6 ? tmp43233 : tmp40314;
  assign tmp43231 = s7 ? tmp39370 : tmp43232;
  assign tmp43230 = s8 ? tmp40206 : tmp43231;
  assign tmp43246 = l1 ? tmp39460 : tmp39541;
  assign tmp43245 = s1 ? tmp43246 : tmp40285;
  assign tmp43250 = l1 ? tmp39972 : tmp39457;
  assign tmp43251 = ~(l1 ? tmp39925 : tmp39649);
  assign tmp43249 = s0 ? tmp43250 : tmp43251;
  assign tmp43253 = l1 ? tmp39972 : tmp40214;
  assign tmp43252 = s0 ? tmp43253 : tmp43251;
  assign tmp43248 = s1 ? tmp43249 : tmp43252;
  assign tmp43255 = s0 ? tmp43253 : tmp40225;
  assign tmp43257 = l1 ? tmp39925 : tmp39649;
  assign tmp43258 = ~(l1 ? tmp39972 : tmp40360);
  assign tmp43256 = ~(s0 ? tmp43257 : tmp43258);
  assign tmp43254 = s1 ? tmp43255 : tmp43256;
  assign tmp43247 = ~(s2 ? tmp43248 : tmp43254);
  assign tmp43244 = s3 ? tmp43245 : tmp43247;
  assign tmp43263 = l1 ? tmp39972 : tmp40360;
  assign tmp43262 = ~(s0 ? tmp43263 : tmp43251);
  assign tmp43261 = s1 ? tmp40303 : tmp43262;
  assign tmp43265 = s0 ? tmp43246 : tmp39420;
  assign tmp43264 = s1 ? tmp43265 : tmp43237;
  assign tmp43260 = s2 ? tmp43261 : tmp43264;
  assign tmp43268 = s0 ? tmp39603 : tmp43257;
  assign tmp43267 = ~(s1 ? tmp43257 : tmp43268);
  assign tmp43266 = ~(s2 ? tmp43239 : tmp43267);
  assign tmp43259 = s3 ? tmp43260 : tmp43266;
  assign tmp43243 = s4 ? tmp43244 : tmp43259;
  assign tmp43274 = ~(l1 ? tmp39972 : tmp39457);
  assign tmp43273 = s1 ? tmp40319 : tmp43274;
  assign tmp43276 = s0 ? tmp43257 : tmp40324;
  assign tmp43275 = s1 ? tmp40320 : tmp43276;
  assign tmp43272 = s2 ? tmp43273 : tmp43275;
  assign tmp43279 = l1 ? tmp39429 : tmp40214;
  assign tmp43278 = s1 ? tmp43279 : tmp39987;
  assign tmp43277 = ~(s2 ? tmp43278 : tmp40328);
  assign tmp43271 = s3 ? tmp43272 : tmp43277;
  assign tmp43270 = s4 ? tmp43271 : tmp40331;
  assign tmp43269 = s5 ? tmp43270 : tmp40270;
  assign tmp43242 = s6 ? tmp43243 : tmp43269;
  assign tmp43241 = s7 ? tmp39370 : tmp43242;
  assign tmp43240 = s8 ? tmp43231 : tmp43241;
  assign tmp43229 = s9 ? tmp43230 : tmp43240;
  assign tmp43281 = s8 ? tmp43231 : tmp39370;
  assign tmp43287 = ~(s2 ? tmp40311 : tmp43267);
  assign tmp43286 = s3 ? tmp43260 : tmp43287;
  assign tmp43285 = s4 ? tmp43244 : tmp43286;
  assign tmp43284 = s6 ? tmp43285 : tmp43269;
  assign tmp43283 = s7 ? tmp40399 : tmp43284;
  assign tmp43290 = s3 ? tmp43235 : tmp40310;
  assign tmp43289 = s4 ? tmp40282 : tmp43290;
  assign tmp43288 = s6 ? tmp43289 : tmp40314;
  assign tmp43282 = s8 ? tmp43283 : tmp43288;
  assign tmp43280 = s9 ? tmp43281 : tmp43282;
  assign tmp43228 = s10 ? tmp43229 : tmp43280;
  assign tmp43294 = s7 ? tmp40207 : tmp43242;
  assign tmp43293 = s8 ? tmp43294 : tmp43232;
  assign tmp43292 = s9 ? tmp43281 : tmp43293;
  assign tmp43291 = s10 ? tmp43229 : tmp43292;
  assign tmp43227 = s11 ? tmp43228 : tmp43291;
  assign tmp43226 = s12 ? tmp39905 : tmp43227;
  assign tmp43135 = s13 ? tmp43136 : tmp43226;
  assign tmp43306 = l2 ? tmp39460 : tmp39398;
  assign tmp43305 = l1 ? tmp43306 : tmp40477;
  assign tmp43308 = l1 ? 1 : tmp39972;
  assign tmp43310 = l2 ? tmp39403 : 0;
  assign tmp43309 = ~(l1 ? tmp43310 : tmp40477);
  assign tmp43307 = ~(s0 ? tmp43308 : tmp43309);
  assign tmp43304 = s1 ? tmp43305 : tmp43307;
  assign tmp43314 = l1 ? tmp39429 : tmp39384;
  assign tmp43316 = l2 ? tmp39460 : 0;
  assign tmp43315 = ~(l1 ? tmp43316 : tmp39926);
  assign tmp43313 = s0 ? tmp43314 : tmp43315;
  assign tmp43318 = l1 ? tmp39429 : tmp39587;
  assign tmp43317 = s0 ? tmp43318 : tmp43315;
  assign tmp43312 = s1 ? tmp43313 : tmp43317;
  assign tmp43321 = ~(l1 ? tmp39785 : tmp39404);
  assign tmp43320 = s0 ? tmp43318 : tmp43321;
  assign tmp43323 = l1 ? tmp43316 : tmp39926;
  assign tmp43324 = ~(l1 ? tmp39429 : tmp40489);
  assign tmp43322 = ~(s0 ? tmp43323 : tmp43324);
  assign tmp43319 = s1 ? tmp43320 : tmp43322;
  assign tmp43311 = ~(s2 ? tmp43312 : tmp43319);
  assign tmp43303 = s3 ? tmp43304 : tmp43311;
  assign tmp43329 = l1 ? tmp39758 : tmp40477;
  assign tmp43328 = s0 ? tmp43329 : tmp39452;
  assign tmp43331 = l1 ? tmp39429 : tmp40489;
  assign tmp43330 = ~(s0 ? tmp43331 : tmp43315);
  assign tmp43327 = s1 ? tmp43328 : tmp43330;
  assign tmp43333 = s0 ? tmp43305 : tmp39452;
  assign tmp43334 = l1 ? tmp39758 : tmp39404;
  assign tmp43332 = s1 ? tmp43333 : tmp43334;
  assign tmp43326 = s2 ? tmp43327 : tmp43332;
  assign tmp43336 = s1 ? tmp43308 : tmp39531;
  assign tmp43338 = s0 ? tmp43323 : tmp39932;
  assign tmp43339 = s0 ? tmp40505 : tmp43323;
  assign tmp43337 = ~(s1 ? tmp43338 : tmp43339);
  assign tmp43335 = ~(s2 ? tmp43336 : tmp43337);
  assign tmp43325 = s3 ? tmp43326 : tmp43335;
  assign tmp43302 = s4 ? tmp43303 : tmp43325;
  assign tmp43346 = l1 ? tmp43310 : tmp40477;
  assign tmp43345 = s0 ? tmp43346 : tmp39452;
  assign tmp43347 = ~(l1 ? tmp39429 : tmp39384);
  assign tmp43344 = s1 ? tmp43345 : tmp43347;
  assign tmp43348 = s1 ? tmp43346 : tmp40172;
  assign tmp43343 = s2 ? tmp43344 : tmp43348;
  assign tmp43351 = s0 ? tmp39456 : tmp43318;
  assign tmp43350 = s1 ? tmp43351 : tmp39967;
  assign tmp43352 = ~(s1 ? tmp40519 : tmp40004);
  assign tmp43349 = ~(s2 ? tmp43350 : tmp43352);
  assign tmp43342 = s3 ? tmp43343 : tmp43349;
  assign tmp43357 = l1 ? tmp43316 : tmp40477;
  assign tmp43356 = s0 ? tmp39635 : tmp43357;
  assign tmp43359 = l1 ? tmp39758 : tmp39478;
  assign tmp43358 = s0 ? tmp43359 : tmp41059;
  assign tmp43355 = s1 ? tmp43356 : tmp43358;
  assign tmp43354 = s2 ? tmp43355 : tmp39999;
  assign tmp43363 = ~(l1 ? tmp39460 : tmp40534);
  assign tmp43362 = s0 ? tmp40532 : tmp43363;
  assign tmp43361 = s1 ? tmp43362 : tmp39987;
  assign tmp43360 = ~(s2 ? tmp43361 : tmp39650);
  assign tmp43353 = s3 ? tmp43354 : tmp43360;
  assign tmp43341 = s4 ? tmp43342 : tmp43353;
  assign tmp43340 = s5 ? tmp43341 : tmp40535;
  assign tmp43301 = s6 ? tmp43302 : tmp43340;
  assign tmp43300 = s7 ? tmp39370 : tmp43301;
  assign tmp43370 = l1 ? tmp43306 : tmp39615;
  assign tmp43372 = ~(l1 ? tmp43310 : tmp39615);
  assign tmp43371 = ~(s0 ? tmp43308 : tmp43372);
  assign tmp43369 = s1 ? tmp43370 : tmp43371;
  assign tmp43376 = l1 ? tmp39429 : tmp39385;
  assign tmp43377 = ~(l1 ? tmp43316 : tmp39623);
  assign tmp43375 = s0 ? tmp43376 : tmp43377;
  assign tmp43379 = l1 ? tmp39429 : tmp39972;
  assign tmp43378 = s0 ? tmp43379 : tmp43377;
  assign tmp43374 = s1 ? tmp43375 : tmp43378;
  assign tmp43381 = s0 ? tmp43379 : tmp43321;
  assign tmp43383 = l1 ? tmp43316 : tmp39623;
  assign tmp43384 = ~(l1 ? tmp39429 : tmp40564);
  assign tmp43382 = ~(s0 ? tmp43383 : tmp43384);
  assign tmp43380 = s1 ? tmp43381 : tmp43382;
  assign tmp43373 = ~(s2 ? tmp43374 : tmp43380);
  assign tmp43368 = s3 ? tmp43369 : tmp43373;
  assign tmp43389 = l1 ? tmp39758 : tmp39615;
  assign tmp43388 = s0 ? tmp43389 : tmp39452;
  assign tmp43391 = l1 ? tmp39429 : tmp40564;
  assign tmp43390 = ~(s0 ? tmp43391 : tmp43377);
  assign tmp43387 = s1 ? tmp43388 : tmp43390;
  assign tmp43393 = s0 ? tmp43370 : tmp39452;
  assign tmp43392 = s1 ? tmp43393 : tmp43334;
  assign tmp43386 = s2 ? tmp43387 : tmp43392;
  assign tmp43397 = l1 ? tmp39925 : tmp39623;
  assign tmp43396 = s0 ? tmp43383 : tmp43397;
  assign tmp43398 = s0 ? tmp40505 : tmp43383;
  assign tmp43395 = ~(s1 ? tmp43396 : tmp43398);
  assign tmp43394 = ~(s2 ? tmp43336 : tmp43395);
  assign tmp43385 = s3 ? tmp43386 : tmp43394;
  assign tmp43367 = s4 ? tmp43368 : tmp43385;
  assign tmp43405 = l1 ? tmp43310 : tmp39615;
  assign tmp43404 = s0 ? tmp43405 : tmp39452;
  assign tmp43406 = ~(l1 ? tmp39429 : tmp39385);
  assign tmp43403 = s1 ? tmp43404 : tmp43406;
  assign tmp43408 = s0 ? tmp43397 : tmp39452;
  assign tmp43407 = s1 ? tmp43405 : tmp43408;
  assign tmp43402 = s2 ? tmp43403 : tmp43407;
  assign tmp43411 = s0 ? tmp39456 : tmp43379;
  assign tmp43412 = s0 ? tmp39456 : tmp40591;
  assign tmp43410 = s1 ? tmp43411 : tmp43412;
  assign tmp43414 = ~(l1 ? tmp39429 : tmp39532);
  assign tmp43413 = ~(s1 ? tmp40519 : tmp43414);
  assign tmp43409 = ~(s2 ? tmp43410 : tmp43413);
  assign tmp43401 = s3 ? tmp43402 : tmp43409;
  assign tmp43416 = s2 ? tmp43355 : tmp40539;
  assign tmp43419 = s0 ? tmp39429 : tmp43363;
  assign tmp43418 = s1 ? tmp43419 : tmp39987;
  assign tmp43417 = ~(s2 ? tmp43418 : tmp39650);
  assign tmp43415 = s3 ? tmp43416 : tmp43417;
  assign tmp43400 = s4 ? tmp43401 : tmp43415;
  assign tmp43399 = s5 ? tmp43400 : tmp40600;
  assign tmp43366 = s6 ? tmp43367 : tmp43399;
  assign tmp43365 = s7 ? tmp39370 : tmp43366;
  assign tmp43364 = s8 ? tmp43300 : tmp43365;
  assign tmp43299 = s9 ? tmp43300 : tmp43364;
  assign tmp43421 = s8 ? tmp43300 : tmp39370;
  assign tmp43429 = s1 ? tmp43411 : tmp40591;
  assign tmp43428 = ~(s2 ? tmp43429 : tmp43413);
  assign tmp43427 = s3 ? tmp43402 : tmp43428;
  assign tmp43426 = s4 ? tmp43427 : tmp43415;
  assign tmp43425 = s5 ? tmp43426 : tmp40600;
  assign tmp43424 = s6 ? tmp43367 : tmp43425;
  assign tmp43423 = s7 ? tmp40613 : tmp43424;
  assign tmp43435 = s1 ? tmp43351 : tmp39968;
  assign tmp43434 = ~(s2 ? tmp43435 : tmp43352);
  assign tmp43433 = s3 ? tmp43343 : tmp43434;
  assign tmp43432 = s4 ? tmp43433 : tmp43353;
  assign tmp43431 = s5 ? tmp43432 : tmp40535;
  assign tmp43430 = s6 ? tmp43302 : tmp43431;
  assign tmp43422 = s8 ? tmp43423 : tmp43430;
  assign tmp43420 = s9 ? tmp43421 : tmp43422;
  assign tmp43298 = s10 ? tmp43299 : tmp43420;
  assign tmp43439 = s7 ? tmp40414 : tmp43366;
  assign tmp43438 = s8 ? tmp43439 : tmp43301;
  assign tmp43437 = s9 ? tmp43421 : tmp43438;
  assign tmp43436 = s10 ? tmp43299 : tmp43437;
  assign tmp43297 = s11 ? tmp43298 : tmp43436;
  assign tmp43448 = l2 ? tmp39460 : tmp39616;
  assign tmp43447 = l1 ? tmp43448 : tmp40633;
  assign tmp43451 = l2 ? tmp39403 : tmp39389;
  assign tmp43450 = ~(l1 ? tmp43451 : tmp40633);
  assign tmp43449 = ~(s0 ? tmp39946 : tmp43450);
  assign tmp43446 = s1 ? tmp43447 : tmp43449;
  assign tmp43455 = l2 ? tmp39460 : tmp39389;
  assign tmp43454 = ~(l1 ? tmp43455 : tmp40643);
  assign tmp43453 = s0 ? tmp40701 : tmp43454;
  assign tmp43458 = ~(l2 ? tmp39403 : tmp39386);
  assign tmp43457 = s0 ? tmp40701 : tmp43458;
  assign tmp43460 = l1 ? tmp43455 : tmp40643;
  assign tmp43461 = ~(l1 ? tmp39630 : tmp40649);
  assign tmp43459 = ~(s0 ? tmp43460 : tmp43461);
  assign tmp43456 = s1 ? tmp43457 : tmp43459;
  assign tmp43452 = ~(s2 ? tmp43453 : tmp43456);
  assign tmp43445 = s3 ? tmp43446 : tmp43452;
  assign tmp43466 = l1 ? tmp39785 : tmp40633;
  assign tmp43465 = s0 ? tmp43466 : tmp40655;
  assign tmp43468 = l1 ? tmp39630 : tmp40649;
  assign tmp43467 = ~(s0 ? tmp43468 : tmp43454);
  assign tmp43464 = s1 ? tmp43465 : tmp43467;
  assign tmp43470 = s0 ? tmp43447 : 0;
  assign tmp43469 = s1 ? tmp43470 : tmp40660;
  assign tmp43463 = s2 ? tmp43464 : tmp43469;
  assign tmp43473 = s0 ? tmp43460 : tmp40665;
  assign tmp43474 = s0 ? tmp40667 : tmp43460;
  assign tmp43472 = ~(s1 ? tmp43473 : tmp43474);
  assign tmp43471 = ~(s2 ? tmp40662 : tmp43472);
  assign tmp43462 = s3 ? tmp43463 : tmp43471;
  assign tmp43444 = s4 ? tmp43445 : tmp43462;
  assign tmp43481 = l1 ? tmp43451 : tmp40633;
  assign tmp43480 = s0 ? tmp43481 : tmp40096;
  assign tmp43479 = s1 ? tmp43480 : tmp40720;
  assign tmp43483 = l1 ? tmp43451 : tmp39376;
  assign tmp43484 = s0 ? tmp40665 : tmp40096;
  assign tmp43482 = s1 ? tmp43483 : tmp43484;
  assign tmp43478 = s2 ? tmp43479 : tmp43482;
  assign tmp43486 = s1 ? tmp40701 : tmp40682;
  assign tmp43488 = ~(s0 ? tmp43468 : tmp40687);
  assign tmp43487 = ~(s1 ? tmp40685 : tmp43488);
  assign tmp43485 = ~(s2 ? tmp43486 : tmp43487);
  assign tmp43477 = s3 ? tmp43478 : tmp43485;
  assign tmp43493 = l1 ? tmp43455 : tmp39376;
  assign tmp43492 = s0 ? tmp40692 : tmp43493;
  assign tmp43491 = s1 ? tmp43492 : tmp40695;
  assign tmp43494 = ~(s1 ? tmp39495 : tmp40701);
  assign tmp43490 = s2 ? tmp43491 : tmp43494;
  assign tmp43498 = ~(l1 ? tmp39681 : tmp39376);
  assign tmp43497 = s0 ? tmp40701 : tmp43498;
  assign tmp43496 = s1 ? tmp43497 : tmp40703;
  assign tmp43495 = ~(s2 ? tmp43496 : tmp39651);
  assign tmp43489 = s3 ? tmp43490 : tmp43495;
  assign tmp43476 = s4 ? tmp43477 : tmp43489;
  assign tmp43503 = l1 ? 1 : tmp39403;
  assign tmp43502 = s1 ? tmp43503 : tmp39661;
  assign tmp43501 = s2 ? tmp40709 : tmp43502;
  assign tmp43500 = s3 ? tmp43501 : tmp40714;
  assign tmp43499 = s4 ? tmp43500 : tmp40717;
  assign tmp43475 = s5 ? tmp43476 : tmp43499;
  assign tmp43443 = s6 ? tmp43444 : tmp43475;
  assign tmp43442 = s7 ? tmp39370 : tmp43443;
  assign tmp43505 = s8 ? tmp43442 : tmp39370;
  assign tmp43511 = s1 ? tmp43497 : tmp40704;
  assign tmp43510 = ~(s2 ? tmp43511 : tmp39651);
  assign tmp43509 = s3 ? tmp43490 : tmp43510;
  assign tmp43508 = s4 ? tmp43477 : tmp43509;
  assign tmp43507 = s5 ? tmp43508 : tmp43499;
  assign tmp43506 = s6 ? tmp43444 : tmp43507;
  assign tmp43504 = s9 ? tmp43505 : tmp43506;
  assign tmp43441 = s10 ? tmp43442 : tmp43504;
  assign tmp43513 = s9 ? tmp43505 : tmp43443;
  assign tmp43512 = s10 ? tmp43442 : tmp43513;
  assign tmp43440 = s11 ? tmp43441 : tmp43512;
  assign tmp43296 = s12 ? tmp43297 : tmp43440;
  assign tmp43524 = s2 ? tmp40968 : tmp41060;
  assign tmp43525 = ~(s2 ? tmp39663 : tmp40977);
  assign tmp43523 = s3 ? tmp43524 : tmp43525;
  assign tmp43522 = s4 ? tmp43523 : tmp41217;
  assign tmp43521 = s5 ? tmp40937 : tmp43522;
  assign tmp43520 = s6 ? tmp40897 : tmp43521;
  assign tmp43519 = s7 ? tmp39370 : tmp43520;
  assign tmp43530 = s3 ? tmp41057 : tmp43525;
  assign tmp43529 = s4 ? tmp43530 : tmp41229;
  assign tmp43528 = s5 ? tmp41029 : tmp43529;
  assign tmp43527 = s6 ? tmp40988 : tmp43528;
  assign tmp43526 = s7 ? tmp39370 : tmp43527;
  assign tmp43518 = s8 ? tmp43519 : tmp43526;
  assign tmp43537 = s2 ? tmp41058 : tmp40971;
  assign tmp43536 = s3 ? tmp43537 : tmp40974;
  assign tmp43539 = s2 ? tmp41063 : tmp40983;
  assign tmp43538 = s3 ? tmp43539 : tmp40984;
  assign tmp43535 = s4 ? tmp43536 : tmp43538;
  assign tmp43534 = s5 ? tmp41029 : tmp43535;
  assign tmp43533 = s6 ? tmp40988 : tmp43534;
  assign tmp43532 = s7 ? tmp39370 : tmp43533;
  assign tmp43531 = s8 ? tmp43526 : tmp43532;
  assign tmp43517 = s9 ? tmp43518 : tmp43531;
  assign tmp43541 = s8 ? tmp43526 : tmp39370;
  assign tmp43549 = ~(l2 ? tmp39379 : tmp39460);
  assign tmp43548 = l1 ? tmp40992 : tmp43549;
  assign tmp43551 = ~(l1 ? tmp40997 : tmp43549);
  assign tmp43550 = ~(s0 ? tmp40995 : tmp43551);
  assign tmp43547 = s1 ? tmp43548 : tmp43550;
  assign tmp43555 = l1 ? tmp39403 : tmp39480;
  assign tmp43557 = ~(l2 ? tmp39430 : tmp39460);
  assign tmp43556 = ~(l1 ? tmp41002 : tmp43557);
  assign tmp43554 = s0 ? tmp43555 : tmp43556;
  assign tmp43559 = l1 ? tmp39403 : tmp39630;
  assign tmp43558 = s0 ? tmp43559 : tmp43556;
  assign tmp43553 = s1 ? tmp43554 : tmp43558;
  assign tmp43561 = s0 ? tmp43559 : tmp41006;
  assign tmp43563 = l1 ? tmp41002 : tmp43557;
  assign tmp43564 = ~(l1 ? tmp39403 : tmp39840);
  assign tmp43562 = ~(s0 ? tmp43563 : tmp43564);
  assign tmp43560 = s1 ? tmp43561 : tmp43562;
  assign tmp43552 = ~(s2 ? tmp43553 : tmp43560);
  assign tmp43546 = s3 ? tmp43547 : tmp43552;
  assign tmp43569 = l1 ? tmp39972 : tmp43549;
  assign tmp43568 = s0 ? tmp43569 : tmp41015;
  assign tmp43571 = l1 ? tmp39403 : tmp39840;
  assign tmp43570 = ~(s0 ? tmp43571 : tmp43556);
  assign tmp43567 = s1 ? tmp43568 : tmp43570;
  assign tmp43573 = s0 ? tmp43548 : tmp40225;
  assign tmp43572 = s1 ? tmp43573 : tmp41020;
  assign tmp43566 = s2 ? tmp43567 : tmp43572;
  assign tmp43577 = l1 ? tmp39379 : tmp43557;
  assign tmp43576 = s0 ? tmp43563 : tmp43577;
  assign tmp43578 = s0 ? tmp41027 : tmp43563;
  assign tmp43575 = ~(s1 ? tmp43576 : tmp43578);
  assign tmp43574 = ~(s2 ? tmp41022 : tmp43575);
  assign tmp43565 = s3 ? tmp43566 : tmp43574;
  assign tmp43545 = s4 ? tmp43546 : tmp43565;
  assign tmp43585 = l1 ? tmp40997 : tmp43549;
  assign tmp43584 = s0 ? tmp43585 : 0;
  assign tmp43586 = ~(l1 ? tmp39403 : tmp39480);
  assign tmp43583 = s1 ? tmp43584 : tmp43586;
  assign tmp43588 = s0 ? tmp43577 : tmp40225;
  assign tmp43587 = s1 ? tmp41036 : tmp43588;
  assign tmp43582 = s2 ? tmp43583 : tmp43587;
  assign tmp43590 = s1 ? tmp43559 : tmp40948;
  assign tmp43589 = ~(s2 ? tmp43590 : tmp41040);
  assign tmp43581 = s3 ? tmp43582 : tmp43589;
  assign tmp43595 = l1 ? tmp41002 : tmp40477;
  assign tmp43594 = s0 ? tmp39635 : tmp43595;
  assign tmp43593 = s1 ? tmp43594 : tmp41047;
  assign tmp43592 = s2 ? tmp43593 : tmp41049;
  assign tmp43599 = ~(l1 ? tmp39475 : tmp40534);
  assign tmp43598 = s0 ? tmp40962 : tmp43599;
  assign tmp43597 = s1 ? tmp43598 : tmp41127;
  assign tmp43596 = ~(s2 ? tmp43597 : tmp39650);
  assign tmp43591 = s3 ? tmp43592 : tmp43596;
  assign tmp43580 = s4 ? tmp43581 : tmp43591;
  assign tmp43601 = s3 ? tmp43537 : tmp41136;
  assign tmp43602 = s3 ? tmp41230 : tmp41142;
  assign tmp43600 = s4 ? tmp43601 : tmp43602;
  assign tmp43579 = s5 ? tmp43580 : tmp43600;
  assign tmp43544 = s6 ? tmp43545 : tmp43579;
  assign tmp43543 = s7 ? tmp43520 : tmp43544;
  assign tmp43542 = s8 ? tmp43543 : tmp43527;
  assign tmp43540 = s9 ? tmp43541 : tmp43542;
  assign tmp43516 = s10 ? tmp43517 : tmp43540;
  assign tmp43610 = s3 ? tmp43539 : tmp41142;
  assign tmp43609 = s4 ? tmp43601 : tmp43610;
  assign tmp43608 = s5 ? tmp43580 : tmp43609;
  assign tmp43607 = s6 ? tmp43545 : tmp43608;
  assign tmp43606 = s7 ? tmp43520 : tmp43607;
  assign tmp43605 = s8 ? tmp43606 : tmp43527;
  assign tmp43604 = s9 ? tmp43541 : tmp43605;
  assign tmp43603 = s10 ? tmp43517 : tmp43604;
  assign tmp43515 = s11 ? tmp43516 : tmp43603;
  assign tmp43619 = s3 ? tmp41310 : tmp43525;
  assign tmp43618 = s4 ? tmp43619 : tmp41532;
  assign tmp43617 = s5 ? tmp41284 : tmp43618;
  assign tmp43616 = s6 ? tmp41247 : tmp43617;
  assign tmp43615 = s7 ? tmp39370 : tmp43616;
  assign tmp43624 = s3 ? tmp41386 : tmp43525;
  assign tmp43623 = s4 ? tmp43624 : tmp41544;
  assign tmp43622 = s5 ? tmp41358 : tmp43623;
  assign tmp43621 = s6 ? tmp41321 : tmp43622;
  assign tmp43620 = s7 ? tmp39370 : tmp43621;
  assign tmp43614 = s8 ? tmp43615 : tmp43620;
  assign tmp43625 = s8 ? tmp43620 : tmp41396;
  assign tmp43613 = s9 ? tmp43614 : tmp43625;
  assign tmp43630 = s5 ? tmp41504 : tmp43618;
  assign tmp43629 = s6 ? tmp41472 : tmp43630;
  assign tmp43628 = s7 ? tmp39370 : tmp43629;
  assign tmp43627 = s8 ? tmp43628 : tmp39370;
  assign tmp43632 = s7 ? tmp43616 : tmp41534;
  assign tmp43633 = s7 ? tmp43621 : tmp43629;
  assign tmp43631 = s8 ? tmp43632 : tmp43633;
  assign tmp43626 = s9 ? tmp43627 : tmp43631;
  assign tmp43612 = s10 ? tmp43613 : tmp43626;
  assign tmp43637 = s7 ? tmp43616 : tmp41397;
  assign tmp43636 = s8 ? tmp43637 : tmp43633;
  assign tmp43635 = s9 ? tmp43627 : tmp43636;
  assign tmp43634 = s10 ? tmp43613 : tmp43635;
  assign tmp43611 = s11 ? tmp43612 : tmp43634;
  assign tmp43514 = s12 ? tmp43515 : tmp43611;
  assign tmp43295 = s13 ? tmp43296 : tmp43514;
  assign tmp43134 = s14 ? tmp43135 : tmp43295;
  assign tmp43651 = s1 ? tmp42136 : tmp39664;
  assign tmp43650 = ~(s2 ? tmp43651 : tmp42184);
  assign tmp43649 = s3 ? tmp42177 : tmp43650;
  assign tmp43655 = l1 ? tmp40982 : 1;
  assign tmp43654 = s1 ? tmp43655 : tmp42141;
  assign tmp43656 = ~(l1 ? tmp39480 : tmp39801);
  assign tmp43653 = s2 ? tmp43654 : tmp43656;
  assign tmp43652 = s3 ? tmp43653 : tmp42193;
  assign tmp43648 = s4 ? tmp43649 : tmp43652;
  assign tmp43647 = s5 ? tmp42143 : tmp43648;
  assign tmp43646 = s6 ? tmp42110 : tmp43647;
  assign tmp43645 = s7 ? tmp39370 : tmp43646;
  assign tmp43661 = s3 ? tmp42255 : tmp43650;
  assign tmp43660 = s4 ? tmp43661 : tmp43652;
  assign tmp43659 = s5 ? tmp42228 : tmp43660;
  assign tmp43658 = s6 ? tmp42198 : tmp43659;
  assign tmp43657 = s7 ? tmp39370 : tmp43658;
  assign tmp43644 = s8 ? tmp43645 : tmp43657;
  assign tmp43662 = s8 ? tmp43657 : tmp42257;
  assign tmp43643 = s9 ? tmp43644 : tmp43662;
  assign tmp43669 = s3 ? tmp42348 : tmp43650;
  assign tmp43672 = s1 ? tmp43655 : tmp42290;
  assign tmp43673 = ~(l1 ? tmp39480 : tmp40477);
  assign tmp43671 = s2 ? tmp43672 : tmp43673;
  assign tmp43670 = s3 ? tmp43671 : tmp42193;
  assign tmp43668 = s4 ? tmp43669 : tmp43670;
  assign tmp43667 = s5 ? tmp42340 : tmp43668;
  assign tmp43666 = s6 ? tmp42333 : tmp43667;
  assign tmp43665 = s7 ? tmp39370 : tmp43666;
  assign tmp43664 = s8 ? tmp43665 : tmp39370;
  assign tmp43677 = s5 ? tmp42353 : tmp43648;
  assign tmp43676 = s6 ? tmp42110 : tmp43677;
  assign tmp43675 = s7 ? tmp43676 : tmp42361;
  assign tmp43678 = s7 ? tmp43658 : tmp43666;
  assign tmp43674 = s8 ? tmp43675 : tmp43678;
  assign tmp43663 = s9 ? tmp43664 : tmp43674;
  assign tmp43642 = s10 ? tmp43643 : tmp43663;
  assign tmp43682 = s7 ? tmp43646 : tmp42258;
  assign tmp43681 = s8 ? tmp43682 : tmp43678;
  assign tmp43680 = s9 ? tmp43664 : tmp43681;
  assign tmp43679 = s10 ? tmp43643 : tmp43680;
  assign tmp43641 = s11 ? tmp43642 : tmp43679;
  assign tmp43695 = ~(l1 ? tmp39630 : tmp39403);
  assign tmp43694 = s0 ? tmp39516 : tmp43695;
  assign tmp43693 = ~(s1 ? tmp43694 : 1);
  assign tmp43692 = s2 ? tmp42446 : tmp43693;
  assign tmp43691 = s3 ? tmp43692 : tmp42451;
  assign tmp43690 = s4 ? tmp43691 : tmp42454;
  assign tmp43689 = s5 ? tmp42496 : tmp43690;
  assign tmp43688 = s6 ? tmp42464 : tmp43689;
  assign tmp43687 = s7 ? tmp39370 : tmp43688;
  assign tmp43686 = s8 ? tmp42382 : tmp43687;
  assign tmp43685 = s9 ? tmp43686 : tmp43687;
  assign tmp43697 = s8 ? tmp43687 : tmp39370;
  assign tmp43705 = l2 ? tmp39376 : tmp39380;
  assign tmp43704 = l1 ? tmp42268 : tmp43705;
  assign tmp43707 = ~(l1 ? tmp40729 : tmp43705);
  assign tmp43706 = ~(s0 ? tmp39477 : tmp43707);
  assign tmp43703 = s1 ? tmp43704 : tmp43706;
  assign tmp43712 = l2 ? tmp39440 : tmp39380;
  assign tmp43711 = ~(l1 ? tmp40737 : tmp43712);
  assign tmp43710 = s0 ? tmp39477 : tmp43711;
  assign tmp43713 = s0 ? tmp42475 : tmp43711;
  assign tmp43709 = s1 ? tmp43710 : tmp43713;
  assign tmp43716 = l1 ? tmp40737 : tmp43712;
  assign tmp43718 = ~(l2 ? tmp39440 : tmp39380);
  assign tmp43717 = ~(l1 ? tmp40779 : tmp43718);
  assign tmp43715 = ~(s0 ? tmp43716 : tmp43717);
  assign tmp43714 = s1 ? tmp42477 : tmp43715;
  assign tmp43708 = ~(s2 ? tmp43709 : tmp43714);
  assign tmp43702 = s3 ? tmp43703 : tmp43708;
  assign tmp43723 = l1 ? tmp39587 : tmp43705;
  assign tmp43722 = s0 ? tmp43723 : tmp40024;
  assign tmp43725 = l1 ? tmp40779 : tmp43718;
  assign tmp43724 = ~(s0 ? tmp43725 : tmp43711);
  assign tmp43721 = s1 ? tmp43722 : tmp43724;
  assign tmp43727 = s0 ? tmp43704 : tmp40225;
  assign tmp43726 = s1 ? tmp43727 : tmp39569;
  assign tmp43720 = s2 ? tmp43721 : tmp43726;
  assign tmp43731 = l1 ? tmp40705 : tmp43712;
  assign tmp43730 = s0 ? tmp43716 : tmp43731;
  assign tmp43732 = s0 ? tmp42414 : tmp43716;
  assign tmp43729 = ~(s1 ? tmp43730 : tmp43732);
  assign tmp43728 = ~(s2 ? tmp42409 : tmp43729);
  assign tmp43719 = s3 ? tmp43720 : tmp43728;
  assign tmp43701 = s4 ? tmp43702 : tmp43719;
  assign tmp43739 = l1 ? tmp40729 : tmp43705;
  assign tmp43738 = s0 ? tmp43739 : tmp40096;
  assign tmp43737 = s1 ? tmp43738 : tmp40024;
  assign tmp43741 = l1 ? tmp40729 : tmp42707;
  assign tmp43742 = s0 ? tmp43731 : tmp40024;
  assign tmp43740 = s1 ? tmp43741 : tmp43742;
  assign tmp43736 = s2 ? tmp43737 : tmp43740;
  assign tmp43745 = ~(l1 ? tmp40705 : tmp40668);
  assign tmp43744 = s1 ? tmp42475 : tmp43745;
  assign tmp43748 = l1 ? tmp40779 : tmp39459;
  assign tmp43747 = ~(s0 ? tmp43725 : tmp43748);
  assign tmp43746 = ~(s1 ? tmp42428 : tmp43747);
  assign tmp43743 = ~(s2 ? tmp43744 : tmp43746);
  assign tmp43735 = s3 ? tmp43736 : tmp43743;
  assign tmp43753 = l1 ? tmp40737 : tmp42707;
  assign tmp43752 = s0 ? tmp42435 : tmp43753;
  assign tmp43751 = s1 ? tmp43752 : tmp41813;
  assign tmp43754 = ~(l1 ? tmp39402 : tmp39744);
  assign tmp43750 = s2 ? tmp43751 : tmp43754;
  assign tmp43758 = ~(l1 ? tmp42173 : tmp42707);
  assign tmp43757 = s0 ? tmp39743 : tmp43758;
  assign tmp43756 = s1 ? tmp43757 : tmp42577;
  assign tmp43755 = ~(s2 ? tmp43756 : tmp42442);
  assign tmp43749 = s3 ? tmp43750 : tmp43755;
  assign tmp43734 = s4 ? tmp43735 : tmp43749;
  assign tmp43764 = l1 ? tmp40705 : tmp40668;
  assign tmp43763 = s0 ? tmp43764 : tmp42078;
  assign tmp43762 = s1 ? tmp43763 : tmp42078;
  assign tmp43765 = ~(s1 ? tmp43694 : tmp40713);
  assign tmp43761 = s2 ? tmp43762 : tmp43765;
  assign tmp43760 = s3 ? tmp43761 : tmp42601;
  assign tmp43768 = ~(l1 ? tmp39513 : tmp39744);
  assign tmp43767 = s2 ? tmp42456 : tmp43768;
  assign tmp43766 = s3 ? tmp43767 : tmp42607;
  assign tmp43759 = s4 ? tmp43760 : tmp43766;
  assign tmp43733 = s5 ? tmp43734 : tmp43759;
  assign tmp43700 = s6 ? tmp43701 : tmp43733;
  assign tmp43699 = s7 ? tmp42677 : tmp43700;
  assign tmp43771 = s4 ? tmp43691 : tmp42524;
  assign tmp43770 = s5 ? tmp42496 : tmp43771;
  assign tmp43769 = s6 ? tmp42464 : tmp43770;
  assign tmp43698 = s8 ? tmp43699 : tmp43769;
  assign tmp43696 = s9 ? tmp43697 : tmp43698;
  assign tmp43684 = s10 ? tmp43685 : tmp43696;
  assign tmp43781 = l1 ? tmp39513 : tmp39459;
  assign tmp43780 = ~(s1 ? tmp42460 : tmp43781);
  assign tmp43779 = s3 ? tmp43767 : tmp43780;
  assign tmp43778 = s4 ? tmp43760 : tmp43779;
  assign tmp43777 = s5 ? tmp43734 : tmp43778;
  assign tmp43776 = s6 ? tmp43701 : tmp43777;
  assign tmp43775 = s7 ? tmp42383 : tmp43776;
  assign tmp43774 = s8 ? tmp43775 : tmp43688;
  assign tmp43773 = s9 ? tmp43697 : tmp43774;
  assign tmp43772 = s10 ? tmp43685 : tmp43773;
  assign tmp43683 = s11 ? tmp43684 : tmp43772;
  assign tmp43640 = s12 ? tmp43641 : tmp43683;
  assign tmp43639 = s13 ? tmp43640 : tmp42685;
  assign tmp43638 = s14 ? tmp41555 : tmp43639;
  assign tmp43133 = s15 ? tmp43134 : tmp43638;
  assign tmp39361 = s16 ? tmp39362 : tmp43133;
  assign tmp43789 = s8 ? tmp43140 : tmp39749;
  assign tmp43788 = s9 ? tmp43139 : tmp43789;
  assign tmp43792 = s7 ? tmp43209 : tmp39844;
  assign tmp43791 = s8 ? tmp39891 : tmp43792;
  assign tmp43790 = s9 ? tmp39842 : tmp43791;
  assign tmp43787 = s10 ? tmp43788 : tmp43790;
  assign tmp43796 = s7 ? tmp43141 : tmp39844;
  assign tmp43795 = s8 ? tmp39903 : tmp43796;
  assign tmp43794 = s9 ? tmp39842 : tmp43795;
  assign tmp43793 = s10 ? tmp43788 : tmp43794;
  assign tmp43786 = s11 ? tmp43787 : tmp43793;
  assign tmp43801 = s8 ? tmp43231 : tmp40342;
  assign tmp43800 = s9 ? tmp43230 : tmp43801;
  assign tmp43804 = s7 ? tmp43288 : tmp40386;
  assign tmp43803 = s8 ? tmp40398 : tmp43804;
  assign tmp43802 = s9 ? tmp40384 : tmp43803;
  assign tmp43799 = s10 ? tmp43800 : tmp43802;
  assign tmp43808 = s7 ? tmp43232 : tmp40386;
  assign tmp43807 = s8 ? tmp40406 : tmp43808;
  assign tmp43806 = s9 ? tmp40384 : tmp43807;
  assign tmp43805 = s10 ? tmp43800 : tmp43806;
  assign tmp43798 = s11 ? tmp43799 : tmp43805;
  assign tmp43797 = s12 ? tmp39905 : tmp43798;
  assign tmp43785 = s13 ? tmp43786 : tmp43797;
  assign tmp43814 = s8 ? tmp43300 : tmp40544;
  assign tmp43813 = s9 ? tmp43300 : tmp43814;
  assign tmp43817 = s7 ? tmp43430 : tmp40472;
  assign tmp43816 = s8 ? tmp40612 : tmp43817;
  assign tmp43815 = s9 ? tmp40610 : tmp43816;
  assign tmp43812 = s10 ? tmp43813 : tmp43815;
  assign tmp43821 = s7 ? tmp43301 : tmp40472;
  assign tmp43820 = s8 ? tmp40621 : tmp43821;
  assign tmp43819 = s9 ? tmp40610 : tmp43820;
  assign tmp43818 = s10 ? tmp43813 : tmp43819;
  assign tmp43811 = s11 ? tmp43812 : tmp43818;
  assign tmp43826 = s7 ? tmp39370 : tmp40811;
  assign tmp43825 = s8 ? tmp43442 : tmp43826;
  assign tmp43824 = s9 ? tmp43442 : tmp43825;
  assign tmp43828 = s7 ? tmp43506 : tmp40724;
  assign tmp43827 = s9 ? tmp40802 : tmp43828;
  assign tmp43823 = s10 ? tmp43824 : tmp43827;
  assign tmp43831 = s7 ? tmp43443 : tmp40724;
  assign tmp43830 = s9 ? tmp40802 : tmp43831;
  assign tmp43829 = s10 ? tmp43824 : tmp43830;
  assign tmp43822 = s11 ? tmp43823 : tmp43829;
  assign tmp43810 = s12 ? tmp43811 : tmp43822;
  assign tmp43836 = s8 ? tmp40895 : tmp43532;
  assign tmp43837 = s8 ? tmp43532 : tmp41066;
  assign tmp43835 = s9 ? tmp43836 : tmp43837;
  assign tmp43843 = s4 ? tmp43536 : tmp41229;
  assign tmp43842 = s5 ? tmp41029 : tmp43843;
  assign tmp43841 = s6 ? tmp40988 : tmp43842;
  assign tmp43840 = s7 ? tmp43841 : tmp41231;
  assign tmp43839 = s8 ? tmp41213 : tmp43840;
  assign tmp43838 = s9 ? tmp41145 : tmp43839;
  assign tmp43834 = s10 ? tmp43835 : tmp43838;
  assign tmp43847 = s7 ? tmp43533 : tmp41147;
  assign tmp43846 = s8 ? tmp41239 : tmp43847;
  assign tmp43845 = s9 ? tmp41145 : tmp43846;
  assign tmp43844 = s10 ? tmp43835 : tmp43845;
  assign tmp43833 = s11 ? tmp43834 : tmp43844;
  assign tmp43832 = s12 ? tmp43833 : tmp41241;
  assign tmp43809 = s13 ? tmp43810 : tmp43832;
  assign tmp43784 = s14 ? tmp43785 : tmp43809;
  assign tmp43854 = s8 ? tmp43687 : tmp42529;
  assign tmp43853 = s9 ? tmp43686 : tmp43854;
  assign tmp43857 = s7 ? tmp43769 : tmp42612;
  assign tmp43856 = s8 ? tmp42676 : tmp43857;
  assign tmp43855 = s9 ? tmp42610 : tmp43856;
  assign tmp43852 = s10 ? tmp43853 : tmp43855;
  assign tmp43861 = s7 ? tmp43688 : tmp42612;
  assign tmp43860 = s8 ? tmp42684 : tmp43861;
  assign tmp43859 = s9 ? tmp42610 : tmp43860;
  assign tmp43858 = s10 ? tmp43853 : tmp43859;
  assign tmp43851 = s11 ? tmp43852 : tmp43858;
  assign tmp43850 = s12 ? tmp42104 : tmp43851;
  assign tmp43849 = s13 ? tmp43850 : tmp42685;
  assign tmp43848 = s14 ? tmp41555 : tmp43849;
  assign tmp43783 = s15 ? tmp43784 : tmp43848;
  assign tmp43868 = s9 ? tmp43836 : tmp43532;
  assign tmp43870 = s8 ? tmp43532 : tmp39370;
  assign tmp43872 = s7 ? tmp41214 : tmp43544;
  assign tmp43871 = s8 ? tmp43872 : tmp43841;
  assign tmp43869 = s9 ? tmp43870 : tmp43871;
  assign tmp43867 = s10 ? tmp43868 : tmp43869;
  assign tmp43876 = s7 ? tmp40896 : tmp43607;
  assign tmp43875 = s8 ? tmp43876 : tmp43533;
  assign tmp43874 = s9 ? tmp43870 : tmp43875;
  assign tmp43873 = s10 ? tmp43868 : tmp43874;
  assign tmp43866 = s11 ? tmp43867 : tmp43873;
  assign tmp43865 = s12 ? tmp43866 : tmp41241;
  assign tmp43864 = s13 ? tmp43296 : tmp43865;
  assign tmp43863 = s14 ? tmp43135 : tmp43864;
  assign tmp43879 = s12 ? tmp42104 : tmp43683;
  assign tmp43878 = s13 ? tmp43879 : tmp42685;
  assign tmp43877 = s14 ? tmp41555 : tmp43878;
  assign tmp43862 = s15 ? tmp43863 : tmp43877;
  assign tmp43782 = s16 ? tmp43783 : tmp43862;
  assign tmp39360 = ~(s17 ? tmp39361 : tmp43782);
  assign s1n = tmp39360;

  assign tmp43897 = l4 ? 1 : 0;
  assign tmp43896 = l3 ? tmp43897 : 0;
  assign tmp43898 = ~(l3 ? 1 : 0);
  assign tmp43895 = l2 ? tmp43896 : tmp43898;
  assign tmp43901 = ~(l4 ? 1 : 0);
  assign tmp43900 = l3 ? tmp43897 : tmp43901;
  assign tmp43902 = ~(l3 ? tmp43897 : 0);
  assign tmp43899 = ~(l2 ? tmp43900 : tmp43902);
  assign tmp43894 = l1 ? tmp43895 : tmp43899;
  assign tmp43906 = l3 ? 1 : tmp43901;
  assign tmp43905 = l2 ? 1 : tmp43906;
  assign tmp43907 = l2 ? tmp43906 : tmp43902;
  assign tmp43904 = l1 ? tmp43905 : tmp43907;
  assign tmp43910 = l3 ? 1 : 0;
  assign tmp43911 = ~(l3 ? 1 : tmp43901);
  assign tmp43909 = l2 ? tmp43910 : tmp43911;
  assign tmp43912 = ~(l2 ? tmp43900 : tmp43898);
  assign tmp43908 = ~(l1 ? tmp43909 : tmp43912);
  assign tmp43903 = ~(s0 ? tmp43904 : tmp43908);
  assign tmp43893 = s1 ? tmp43894 : tmp43903;
  assign tmp43917 = l2 ? tmp43900 : tmp43902;
  assign tmp43916 = l1 ? tmp43905 : tmp43917;
  assign tmp43915 = s0 ? tmp43904 : tmp43916;
  assign tmp43920 = l2 ? tmp43910 : tmp43898;
  assign tmp43921 = ~(l2 ? tmp43900 : tmp43911);
  assign tmp43919 = l1 ? tmp43920 : tmp43921;
  assign tmp43922 = ~(l1 ? tmp43905 : tmp43917);
  assign tmp43918 = ~(s0 ? tmp43919 : tmp43922);
  assign tmp43914 = s1 ? tmp43915 : tmp43918;
  assign tmp43925 = ~(l1 ? 1 : tmp43907);
  assign tmp43924 = s0 ? tmp43919 : tmp43925;
  assign tmp43928 = l2 ? tmp43896 : tmp43911;
  assign tmp43927 = ~(l1 ? tmp43928 : tmp43899);
  assign tmp43926 = ~(s0 ? tmp43916 : tmp43927);
  assign tmp43923 = ~(s1 ? tmp43924 : tmp43926);
  assign tmp43913 = ~(s2 ? tmp43914 : tmp43923);
  assign tmp43892 = s3 ? tmp43893 : tmp43913;
  assign tmp43934 = l2 ? tmp43910 : tmp43902;
  assign tmp43933 = l1 ? tmp43934 : tmp43912;
  assign tmp43936 = l2 ? 1 : tmp43902;
  assign tmp43935 = ~(l1 ? tmp43905 : tmp43936);
  assign tmp43932 = s0 ? tmp43933 : tmp43935;
  assign tmp43938 = l1 ? tmp43928 : tmp43899;
  assign tmp43937 = s0 ? tmp43938 : tmp43922;
  assign tmp43931 = s1 ? tmp43932 : tmp43937;
  assign tmp43941 = l1 ? tmp43907 : 1;
  assign tmp43940 = s0 ? tmp43894 : tmp43941;
  assign tmp43944 = l2 ? tmp43906 : 1;
  assign tmp43943 = l1 ? tmp43905 : tmp43944;
  assign tmp43945 = ~(l1 ? tmp43907 : tmp43936);
  assign tmp43942 = ~(s0 ? tmp43943 : tmp43945);
  assign tmp43939 = s1 ? tmp43940 : tmp43942;
  assign tmp43930 = s2 ? tmp43931 : tmp43939;
  assign tmp43950 = ~(l2 ? tmp43896 : 0);
  assign tmp43949 = l1 ? 1 : tmp43950;
  assign tmp43948 = s0 ? tmp43949 : tmp43904;
  assign tmp43952 = l1 ? tmp43907 : tmp43936;
  assign tmp43955 = l3 ? tmp43897 : 1;
  assign tmp43954 = l2 ? tmp43955 : 1;
  assign tmp43953 = ~(l1 ? 1 : tmp43954);
  assign tmp43951 = ~(s0 ? tmp43952 : tmp43953);
  assign tmp43947 = s1 ? tmp43948 : tmp43951;
  assign tmp43959 = l2 ? tmp43896 : tmp43897;
  assign tmp43958 = ~(l1 ? tmp43959 : tmp43899);
  assign tmp43957 = s0 ? tmp43916 : tmp43958;
  assign tmp43963 = l3 ? 1 : tmp43897;
  assign tmp43962 = l2 ? tmp43963 : tmp43897;
  assign tmp43961 = l1 ? tmp43897 : tmp43962;
  assign tmp43960 = ~(s0 ? tmp43961 : tmp43922);
  assign tmp43956 = s1 ? tmp43957 : tmp43960;
  assign tmp43946 = ~(s2 ? tmp43947 : tmp43956);
  assign tmp43929 = s3 ? tmp43930 : tmp43946;
  assign tmp43891 = s4 ? tmp43892 : tmp43929;
  assign tmp43970 = l1 ? tmp43909 : tmp43912;
  assign tmp43971 = l1 ? tmp43936 : tmp43950;
  assign tmp43969 = s0 ? tmp43970 : tmp43971;
  assign tmp43973 = ~(l1 ? tmp43905 : tmp43907);
  assign tmp43972 = s0 ? tmp43936 : tmp43973;
  assign tmp43968 = s1 ? tmp43969 : tmp43972;
  assign tmp43976 = ~(l1 ? tmp43905 : tmp43944);
  assign tmp43975 = s0 ? tmp43936 : tmp43976;
  assign tmp43978 = l1 ? tmp43959 : tmp43899;
  assign tmp43979 = l1 ? tmp43944 : 1;
  assign tmp43977 = s0 ? tmp43978 : tmp43979;
  assign tmp43974 = s1 ? tmp43975 : tmp43977;
  assign tmp43967 = s2 ? tmp43968 : tmp43974;
  assign tmp43984 = ~(l2 ? tmp43897 : tmp43896);
  assign tmp43983 = l1 ? tmp43944 : tmp43984;
  assign tmp43982 = s0 ? tmp43983 : tmp43973;
  assign tmp43987 = l2 ? tmp43900 : 1;
  assign tmp43986 = ~(l1 ? tmp43905 : tmp43987);
  assign tmp43985 = s0 ? tmp43983 : tmp43986;
  assign tmp43981 = s1 ? tmp43982 : tmp43985;
  assign tmp43991 = l2 ? tmp43955 : tmp43897;
  assign tmp43992 = l2 ? 1 : tmp43955;
  assign tmp43990 = l1 ? tmp43991 : tmp43992;
  assign tmp43989 = s0 ? tmp43961 : tmp43990;
  assign tmp43994 = l1 ? tmp43905 : tmp43987;
  assign tmp43996 = l2 ? tmp43963 : tmp43896;
  assign tmp43995 = ~(l1 ? tmp43959 : tmp43996);
  assign tmp43993 = ~(s0 ? tmp43994 : tmp43995);
  assign tmp43988 = s1 ? tmp43989 : tmp43993;
  assign tmp43980 = s2 ? tmp43981 : tmp43988;
  assign tmp43966 = s3 ? tmp43967 : tmp43980;
  assign tmp44001 = l1 ? 1 : tmp43954;
  assign tmp44000 = s0 ? tmp44001 : tmp43927;
  assign tmp44003 = l1 ? tmp43907 : tmp43950;
  assign tmp44005 = l2 ? tmp43963 : 1;
  assign tmp44004 = l1 ? tmp43944 : tmp44005;
  assign tmp44002 = ~(s0 ? tmp44003 : tmp44004);
  assign tmp43999 = s1 ? tmp44000 : tmp44002;
  assign tmp44009 = l2 ? tmp43906 : tmp43901;
  assign tmp44008 = l1 ? tmp44009 : 1;
  assign tmp44011 = l2 ? tmp43910 : 1;
  assign tmp44010 = l1 ? tmp43906 : tmp44011;
  assign tmp44007 = s0 ? tmp44008 : tmp44010;
  assign tmp44013 = ~(l1 ? tmp44009 : 1);
  assign tmp44012 = ~(s0 ? tmp43943 : tmp44013);
  assign tmp44006 = ~(s1 ? tmp44007 : tmp44012);
  assign tmp43998 = s2 ? tmp43999 : tmp44006;
  assign tmp44017 = l1 ? tmp44005 : tmp43912;
  assign tmp44016 = s0 ? tmp44017 : tmp43976;
  assign tmp44019 = l1 ? tmp43897 : tmp43996;
  assign tmp44018 = s0 ? tmp44010 : tmp44019;
  assign tmp44015 = s1 ? tmp44016 : tmp44018;
  assign tmp44021 = l1 ? tmp43954 : tmp43992;
  assign tmp44023 = ~(l1 ? tmp43954 : tmp43992);
  assign tmp44022 = ~(s0 ? tmp44001 : tmp44023);
  assign tmp44020 = s1 ? tmp44021 : tmp44022;
  assign tmp44014 = ~(s2 ? tmp44015 : tmp44020);
  assign tmp43997 = ~(s3 ? tmp43998 : tmp44014);
  assign tmp43965 = s4 ? tmp43966 : tmp43997;
  assign tmp44028 = s0 ? tmp43994 : tmp44001;
  assign tmp44031 = l2 ? tmp43963 : tmp43955;
  assign tmp44030 = ~(l1 ? tmp44031 : tmp44005);
  assign tmp44029 = s0 ? tmp44001 : tmp44030;
  assign tmp44027 = s1 ? tmp44028 : tmp44029;
  assign tmp44034 = l1 ? tmp43992 : tmp44011;
  assign tmp44033 = s0 ? tmp44034 : tmp43976;
  assign tmp44036 = l1 ? tmp43905 : 1;
  assign tmp44038 = ~(l2 ? tmp43896 : tmp43911);
  assign tmp44037 = l1 ? tmp44005 : tmp44038;
  assign tmp44035 = ~(s0 ? tmp44036 : tmp44037);
  assign tmp44032 = ~(s1 ? tmp44033 : tmp44035);
  assign tmp44026 = s2 ? tmp44027 : tmp44032;
  assign tmp44042 = l1 ? tmp44005 : tmp43905;
  assign tmp44044 = l2 ? 1 : tmp43963;
  assign tmp44045 = l2 ? 1 : tmp43897;
  assign tmp44043 = ~(l1 ? tmp44044 : tmp44045);
  assign tmp44041 = s0 ? tmp44042 : tmp44043;
  assign tmp44047 = l1 ? tmp44044 : tmp43992;
  assign tmp44046 = ~(s0 ? tmp44047 : tmp43953);
  assign tmp44040 = s1 ? tmp44041 : tmp44046;
  assign tmp44050 = ~(l1 ? tmp43955 : tmp43962);
  assign tmp44049 = s0 ? tmp44001 : tmp44050;
  assign tmp44052 = l1 ? tmp43955 : tmp44031;
  assign tmp44054 = l2 ? tmp43963 : tmp43910;
  assign tmp44053 = l1 ? tmp44005 : tmp44054;
  assign tmp44051 = ~(s0 ? tmp44052 : tmp44053);
  assign tmp44048 = s1 ? tmp44049 : tmp44051;
  assign tmp44039 = s2 ? tmp44040 : tmp44048;
  assign tmp44025 = s3 ? tmp44026 : tmp44039;
  assign tmp44059 = l1 ? tmp43905 : tmp44005;
  assign tmp44060 = l1 ? tmp43962 : tmp44044;
  assign tmp44058 = s0 ? tmp44059 : tmp44060;
  assign tmp44062 = l1 ? tmp44045 : 1;
  assign tmp44061 = s0 ? tmp44062 : tmp43961;
  assign tmp44057 = s1 ? tmp44058 : tmp44061;
  assign tmp44065 = ~(l1 ? tmp43962 : tmp43912);
  assign tmp44064 = s0 ? tmp44001 : tmp44065;
  assign tmp44066 = s0 ? tmp44037 : tmp44042;
  assign tmp44063 = ~(s1 ? tmp44064 : tmp44066);
  assign tmp44056 = s2 ? tmp44057 : tmp44063;
  assign tmp44070 = l1 ? tmp43962 : tmp44045;
  assign tmp44069 = s0 ? tmp44034 : tmp44070;
  assign tmp44071 = ~(s0 ? tmp44001 : tmp44036);
  assign tmp44068 = s1 ? tmp44069 : tmp44071;
  assign tmp44073 = s0 ? tmp44052 : tmp44059;
  assign tmp44074 = s0 ? tmp44047 : tmp44062;
  assign tmp44072 = s1 ? tmp44073 : tmp44074;
  assign tmp44067 = s2 ? tmp44068 : tmp44072;
  assign tmp44055 = ~(s3 ? tmp44056 : tmp44067);
  assign tmp44024 = ~(s4 ? tmp44025 : tmp44055);
  assign tmp43964 = s5 ? tmp43965 : tmp44024;
  assign tmp43890 = s6 ? tmp43891 : tmp43964;
  assign tmp44079 = l1 ? tmp43936 : tmp44038;
  assign tmp44081 = l1 ? tmp43905 : tmp43934;
  assign tmp44082 = ~(l1 ? tmp43936 : tmp44038);
  assign tmp44080 = ~(s0 ? tmp44081 : tmp44082);
  assign tmp44078 = s1 ? tmp44079 : tmp44080;
  assign tmp44087 = l2 ? tmp43910 : tmp43906;
  assign tmp44086 = l1 ? tmp44087 : tmp43907;
  assign tmp44089 = l2 ? tmp43897 : tmp43896;
  assign tmp44088 = l1 ? tmp44089 : tmp43909;
  assign tmp44085 = s0 ? tmp44086 : tmp44088;
  assign tmp44091 = ~(l1 ? tmp44089 : tmp43909);
  assign tmp44090 = ~(s0 ? tmp44079 : tmp44091);
  assign tmp44084 = s1 ? tmp44085 : tmp44090;
  assign tmp44093 = s0 ? tmp44079 : tmp43925;
  assign tmp44095 = ~(l1 ? tmp43907 : tmp44038);
  assign tmp44094 = ~(s0 ? tmp44088 : tmp44095);
  assign tmp44092 = ~(s1 ? tmp44093 : tmp44094);
  assign tmp44083 = ~(s2 ? tmp44084 : tmp44092);
  assign tmp44077 = s3 ? tmp44078 : tmp44083;
  assign tmp44099 = s0 ? tmp44079 : tmp43935;
  assign tmp44101 = l1 ? tmp43907 : tmp44038;
  assign tmp44100 = s0 ? tmp44101 : tmp44091;
  assign tmp44098 = s1 ? tmp44099 : tmp44100;
  assign tmp44103 = s0 ? tmp44079 : tmp43941;
  assign tmp44104 = ~(l1 ? tmp43905 : tmp44011);
  assign tmp44102 = s1 ? tmp44103 : tmp44104;
  assign tmp44097 = s2 ? tmp44098 : tmp44102;
  assign tmp44107 = l1 ? tmp43991 : tmp43962;
  assign tmp44106 = s1 ? tmp44081 : tmp44107;
  assign tmp44111 = ~(l2 ? tmp43910 : tmp43911);
  assign tmp44110 = ~(l1 ? tmp43944 : tmp44111);
  assign tmp44109 = s0 ? tmp44088 : tmp44110;
  assign tmp44112 = ~(s0 ? tmp44001 : tmp44091);
  assign tmp44108 = s1 ? tmp44109 : tmp44112;
  assign tmp44105 = ~(s2 ? tmp44106 : tmp44108);
  assign tmp44096 = s3 ? tmp44097 : tmp44105;
  assign tmp44076 = s4 ? tmp44077 : tmp44096;
  assign tmp44118 = s0 ? tmp44079 : tmp43971;
  assign tmp44119 = ~(l1 ? tmp44087 : tmp43907);
  assign tmp44117 = s1 ? tmp44118 : tmp44119;
  assign tmp44122 = l2 ? tmp43910 : tmp43896;
  assign tmp44123 = l2 ? tmp43910 : tmp43963;
  assign tmp44121 = l1 ? tmp44122 : tmp44123;
  assign tmp44125 = l1 ? tmp43944 : tmp44111;
  assign tmp44124 = ~(s0 ? tmp44125 : tmp43979);
  assign tmp44120 = ~(s1 ? tmp44121 : tmp44124);
  assign tmp44116 = s2 ? tmp44117 : tmp44120;
  assign tmp44129 = l2 ? tmp43910 : tmp43900;
  assign tmp44128 = l1 ? tmp44129 : tmp43934;
  assign tmp44131 = l2 ? tmp43910 : tmp43897;
  assign tmp44130 = l1 ? tmp44089 : tmp44131;
  assign tmp44127 = s1 ? tmp44128 : tmp44130;
  assign tmp44135 = l2 ? tmp43955 : tmp43906;
  assign tmp44134 = ~(l1 ? tmp43944 : tmp44135);
  assign tmp44133 = ~(s0 ? tmp44130 : tmp44134);
  assign tmp44132 = ~(s1 ? tmp44001 : tmp44133);
  assign tmp44126 = ~(s2 ? tmp44127 : tmp44132);
  assign tmp44115 = s3 ? tmp44116 : tmp44126;
  assign tmp44140 = l1 ? tmp43955 : tmp43962;
  assign tmp44139 = s0 ? tmp44140 : tmp44095;
  assign tmp44141 = ~(s0 ? tmp44003 : tmp43979);
  assign tmp44138 = s1 ? tmp44139 : tmp44141;
  assign tmp44144 = l1 ? tmp44087 : tmp44123;
  assign tmp44143 = ~(s0 ? tmp44144 : tmp44013);
  assign tmp44142 = ~(s1 ? tmp44008 : tmp44143);
  assign tmp44137 = s2 ? tmp44138 : tmp44142;
  assign tmp44148 = l1 ? 1 : tmp44038;
  assign tmp44150 = l2 ? tmp43896 : tmp43900;
  assign tmp44149 = ~(l1 ? tmp44150 : tmp44131);
  assign tmp44147 = s0 ? tmp44148 : tmp44149;
  assign tmp44151 = l1 ? 1 : tmp44135;
  assign tmp44146 = s1 ? tmp44147 : tmp44151;
  assign tmp44153 = ~(l1 ? tmp43991 : tmp43962);
  assign tmp44152 = s1 ? tmp44001 : tmp44153;
  assign tmp44145 = ~(s2 ? tmp44146 : tmp44152);
  assign tmp44136 = ~(s3 ? tmp44137 : tmp44145);
  assign tmp44114 = s4 ? tmp44115 : tmp44136;
  assign tmp44159 = l1 ? tmp43955 : 1;
  assign tmp44158 = s0 ? tmp44130 : tmp44159;
  assign tmp44157 = s1 ? tmp44158 : 0;
  assign tmp44162 = l2 ? tmp43963 : tmp43906;
  assign tmp44161 = l1 ? tmp44162 : tmp43944;
  assign tmp44163 = l1 ? tmp44162 : 1;
  assign tmp44160 = s1 ? tmp44161 : tmp44163;
  assign tmp44156 = s2 ? tmp44157 : tmp44160;
  assign tmp44166 = ~(l1 ? tmp44045 : tmp43992);
  assign tmp44165 = s1 ? 1 : tmp44166;
  assign tmp44168 = l1 ? 1 : tmp43905;
  assign tmp44167 = s1 ? 1 : tmp44168;
  assign tmp44164 = ~(s2 ? tmp44165 : tmp44167);
  assign tmp44155 = s3 ? tmp44156 : tmp44164;
  assign tmp44171 = s1 ? 1 : tmp44001;
  assign tmp44170 = s2 ? tmp44171 : tmp44148;
  assign tmp44173 = ~(l1 ? tmp44089 : tmp43962);
  assign tmp44172 = s1 ? tmp44001 : tmp44173;
  assign tmp44169 = ~(s3 ? tmp44170 : tmp44172);
  assign tmp44154 = ~(s4 ? tmp44155 : tmp44169);
  assign tmp44113 = s5 ? tmp44114 : tmp44154;
  assign tmp44075 = s6 ? tmp44076 : tmp44113;
  assign tmp43889 = s7 ? tmp43890 : tmp44075;
  assign tmp44179 = ~(s0 ? tmp44081 : tmp44095);
  assign tmp44178 = s1 ? tmp44101 : tmp44179;
  assign tmp44183 = l1 ? tmp44162 : tmp43907;
  assign tmp44182 = s0 ? tmp44183 : tmp44088;
  assign tmp44184 = ~(s0 ? tmp44101 : tmp44091);
  assign tmp44181 = s1 ? tmp44182 : tmp44184;
  assign tmp44186 = s0 ? tmp44101 : tmp43925;
  assign tmp44185 = ~(s1 ? tmp44186 : tmp44094);
  assign tmp44180 = ~(s2 ? tmp44181 : tmp44185);
  assign tmp44177 = s3 ? tmp44178 : tmp44180;
  assign tmp44190 = s0 ? tmp44101 : tmp43935;
  assign tmp44189 = s1 ? tmp44190 : tmp44100;
  assign tmp44192 = s0 ? tmp44101 : tmp43941;
  assign tmp44191 = s1 ? tmp44192 : tmp44104;
  assign tmp44188 = s2 ? tmp44189 : tmp44191;
  assign tmp44187 = s3 ? tmp44188 : tmp44105;
  assign tmp44176 = s4 ? tmp44177 : tmp44187;
  assign tmp44198 = s0 ? tmp44101 : tmp43971;
  assign tmp44199 = ~(l1 ? tmp44162 : tmp43907);
  assign tmp44197 = s1 ? tmp44198 : tmp44199;
  assign tmp44201 = l1 ? tmp43996 : tmp44123;
  assign tmp44200 = ~(s1 ? tmp44201 : tmp44124);
  assign tmp44196 = s2 ? tmp44197 : tmp44200;
  assign tmp44205 = l2 ? tmp43963 : tmp43900;
  assign tmp44204 = l1 ? tmp44205 : tmp43934;
  assign tmp44203 = s1 ? tmp44204 : tmp44130;
  assign tmp44202 = ~(s2 ? tmp44203 : tmp44132);
  assign tmp44195 = s3 ? tmp44196 : tmp44202;
  assign tmp44208 = l1 ? tmp44162 : tmp44123;
  assign tmp44207 = s2 ? tmp44138 : tmp44208;
  assign tmp44213 = l2 ? tmp43897 : tmp43900;
  assign tmp44212 = ~(l1 ? tmp44213 : tmp44131);
  assign tmp44211 = s0 ? tmp44148 : tmp44212;
  assign tmp44210 = s1 ? tmp44211 : tmp44151;
  assign tmp44209 = ~(s2 ? tmp44210 : tmp44152);
  assign tmp44206 = ~(s3 ? tmp44207 : tmp44209);
  assign tmp44194 = s4 ? tmp44195 : tmp44206;
  assign tmp44193 = s5 ? tmp44194 : tmp44154;
  assign tmp44175 = s6 ? tmp44176 : tmp44193;
  assign tmp44174 = s7 ? tmp43890 : tmp44175;
  assign tmp43888 = s8 ? tmp43889 : tmp44174;
  assign tmp44221 = l1 ? tmp43906 : tmp43934;
  assign tmp44220 = ~(s0 ? tmp44221 : tmp44082);
  assign tmp44219 = s1 ? tmp44079 : tmp44220;
  assign tmp44225 = l1 ? tmp43896 : tmp43909;
  assign tmp44224 = s0 ? tmp44086 : tmp44225;
  assign tmp44227 = ~(l1 ? tmp43896 : tmp43909);
  assign tmp44226 = ~(s0 ? tmp44079 : tmp44227);
  assign tmp44223 = s1 ? tmp44224 : tmp44226;
  assign tmp44230 = ~(l1 ? tmp43944 : tmp43907);
  assign tmp44229 = s0 ? tmp44079 : tmp44230;
  assign tmp44231 = ~(s0 ? tmp44225 : tmp44082);
  assign tmp44228 = ~(s1 ? tmp44229 : tmp44231);
  assign tmp44222 = ~(s2 ? tmp44223 : tmp44228);
  assign tmp44218 = s3 ? tmp44219 : tmp44222;
  assign tmp44236 = ~(l1 ? tmp43906 : tmp43936);
  assign tmp44235 = s0 ? tmp44079 : tmp44236;
  assign tmp44237 = s0 ? tmp44079 : tmp44227;
  assign tmp44234 = s1 ? tmp44235 : tmp44237;
  assign tmp44240 = l1 ? tmp43936 : 1;
  assign tmp44239 = s0 ? tmp44079 : tmp44240;
  assign tmp44241 = ~(l1 ? tmp43906 : tmp44011);
  assign tmp44238 = s1 ? tmp44239 : tmp44241;
  assign tmp44233 = s2 ? tmp44234 : tmp44238;
  assign tmp44243 = s1 ? tmp44221 : tmp44107;
  assign tmp44246 = ~(l1 ? 1 : tmp44111);
  assign tmp44245 = s0 ? tmp44225 : tmp44246;
  assign tmp44247 = ~(s0 ? tmp44001 : tmp44227);
  assign tmp44244 = s1 ? tmp44245 : tmp44247;
  assign tmp44242 = ~(s2 ? tmp44243 : tmp44244);
  assign tmp44232 = s3 ? tmp44233 : tmp44242;
  assign tmp44217 = s4 ? tmp44218 : tmp44232;
  assign tmp44254 = l1 ? 1 : tmp44111;
  assign tmp44253 = ~(s0 ? tmp44254 : 1);
  assign tmp44252 = ~(s1 ? tmp44121 : tmp44253);
  assign tmp44251 = s2 ? tmp44117 : tmp44252;
  assign tmp44258 = l1 ? tmp43896 : tmp44131;
  assign tmp44259 = ~(l1 ? 1 : tmp44135);
  assign tmp44257 = ~(s0 ? tmp44258 : tmp44259);
  assign tmp44256 = ~(s1 ? tmp44001 : tmp44257);
  assign tmp44255 = ~(s2 ? tmp44127 : tmp44256);
  assign tmp44250 = s3 ? tmp44251 : tmp44255;
  assign tmp44263 = s0 ? tmp44140 : tmp44082;
  assign tmp44264 = ~(s0 ? tmp43971 : 1);
  assign tmp44262 = s1 ? tmp44263 : tmp44264;
  assign tmp44261 = s2 ? tmp44262 : tmp44144;
  assign tmp44260 = ~(s3 ? tmp44261 : tmp44145);
  assign tmp44249 = s4 ? tmp44250 : tmp44260;
  assign tmp44248 = s5 ? tmp44249 : tmp44154;
  assign tmp44216 = s6 ? tmp44217 : tmp44248;
  assign tmp44215 = s7 ? tmp43890 : tmp44216;
  assign tmp44214 = s8 ? tmp44174 : tmp44215;
  assign tmp43887 = s9 ? tmp43888 : tmp44214;
  assign tmp44266 = s8 ? tmp44215 : tmp43890;
  assign tmp44275 = ~(l1 ? tmp44087 : tmp44123);
  assign tmp44274 = ~(s1 ? tmp44008 : tmp44275);
  assign tmp44273 = s2 ? tmp44138 : tmp44274;
  assign tmp44272 = ~(s3 ? tmp44273 : tmp44145);
  assign tmp44271 = s4 ? tmp44115 : tmp44272;
  assign tmp44270 = s5 ? tmp44271 : tmp44154;
  assign tmp44269 = s6 ? tmp44076 : tmp44270;
  assign tmp44268 = s7 ? tmp44269 : tmp44216;
  assign tmp44276 = s7 ? tmp44175 : tmp44216;
  assign tmp44267 = s8 ? tmp44268 : tmp44276;
  assign tmp44265 = s9 ? tmp44266 : tmp44267;
  assign tmp43886 = s10 ? tmp43887 : tmp44265;
  assign tmp44280 = s7 ? tmp44075 : tmp44216;
  assign tmp44279 = s8 ? tmp44280 : tmp44276;
  assign tmp44278 = s9 ? tmp44266 : tmp44279;
  assign tmp44277 = s10 ? tmp43887 : tmp44278;
  assign tmp43885 = s11 ? tmp43886 : tmp44277;
  assign tmp44292 = ~(s0 ? tmp44088 : tmp44082);
  assign tmp44291 = ~(s1 ? tmp44093 : tmp44292);
  assign tmp44290 = ~(s2 ? tmp44084 : tmp44291);
  assign tmp44289 = s3 ? tmp44219 : tmp44290;
  assign tmp44296 = s0 ? tmp44079 : tmp44091;
  assign tmp44295 = s1 ? tmp44235 : tmp44296;
  assign tmp44298 = ~(s0 ? tmp44010 : tmp43945);
  assign tmp44297 = s1 ? tmp44103 : tmp44298;
  assign tmp44294 = s2 ? tmp44295 : tmp44297;
  assign tmp44301 = ~(s0 ? tmp43952 : tmp44153);
  assign tmp44300 = s1 ? tmp44221 : tmp44301;
  assign tmp44299 = ~(s2 ? tmp44300 : tmp44108);
  assign tmp44293 = s3 ? tmp44294 : tmp44299;
  assign tmp44288 = s4 ? tmp44289 : tmp44293;
  assign tmp44307 = s0 ? tmp43936 : tmp44119;
  assign tmp44306 = s1 ? tmp44118 : tmp44307;
  assign tmp44310 = ~(l1 ? tmp44122 : tmp44123);
  assign tmp44309 = s0 ? tmp43936 : tmp44310;
  assign tmp44311 = s0 ? tmp44125 : tmp43979;
  assign tmp44308 = s1 ? tmp44309 : tmp44311;
  assign tmp44305 = s2 ? tmp44306 : tmp44308;
  assign tmp44315 = ~(l1 ? tmp44129 : tmp43934);
  assign tmp44314 = s0 ? tmp43983 : tmp44315;
  assign tmp44317 = ~(l1 ? tmp44089 : tmp44131);
  assign tmp44316 = s0 ? tmp43983 : tmp44317;
  assign tmp44313 = s1 ? tmp44314 : tmp44316;
  assign tmp44318 = s1 ? tmp44001 : tmp44133;
  assign tmp44312 = s2 ? tmp44313 : tmp44318;
  assign tmp44304 = s3 ? tmp44305 : tmp44312;
  assign tmp44303 = s4 ? tmp44304 : tmp44260;
  assign tmp44302 = s5 ? tmp44303 : tmp44154;
  assign tmp44287 = s6 ? tmp44288 : tmp44302;
  assign tmp44286 = s7 ? tmp43890 : tmp44287;
  assign tmp44326 = s0 ? tmp43936 : tmp44199;
  assign tmp44325 = s1 ? tmp44198 : tmp44326;
  assign tmp44329 = ~(l1 ? tmp43996 : tmp44123);
  assign tmp44328 = s0 ? tmp43936 : tmp44329;
  assign tmp44327 = s1 ? tmp44328 : tmp44311;
  assign tmp44324 = s2 ? tmp44325 : tmp44327;
  assign tmp44323 = s3 ? tmp44324 : tmp44202;
  assign tmp44322 = s4 ? tmp44323 : tmp44206;
  assign tmp44321 = s5 ? tmp44322 : tmp44154;
  assign tmp44320 = s6 ? tmp44176 : tmp44321;
  assign tmp44319 = s7 ? tmp43890 : tmp44320;
  assign tmp44285 = s8 ? tmp44286 : tmp44319;
  assign tmp44338 = s0 ? tmp44254 : 1;
  assign tmp44337 = s1 ? tmp44309 : tmp44338;
  assign tmp44336 = s2 ? tmp44306 : tmp44337;
  assign tmp44335 = s3 ? tmp44336 : tmp44255;
  assign tmp44334 = s4 ? tmp44335 : tmp44260;
  assign tmp44333 = s5 ? tmp44334 : tmp44154;
  assign tmp44332 = s6 ? tmp44217 : tmp44333;
  assign tmp44331 = s7 ? tmp43890 : tmp44332;
  assign tmp44330 = s8 ? tmp44319 : tmp44331;
  assign tmp44284 = s9 ? tmp44285 : tmp44330;
  assign tmp44340 = s8 ? tmp44331 : tmp43890;
  assign tmp44346 = ~(s2 ? tmp44243 : tmp44108);
  assign tmp44345 = s3 ? tmp44294 : tmp44346;
  assign tmp44344 = s4 ? tmp44289 : tmp44345;
  assign tmp44350 = s2 ? tmp44306 : tmp44120;
  assign tmp44352 = s1 ? tmp44314 : tmp44317;
  assign tmp44351 = s2 ? tmp44352 : tmp44318;
  assign tmp44349 = s3 ? tmp44350 : tmp44351;
  assign tmp44348 = s4 ? tmp44349 : tmp44260;
  assign tmp44347 = s5 ? tmp44348 : tmp44154;
  assign tmp44343 = s6 ? tmp44344 : tmp44347;
  assign tmp44357 = s2 ? tmp44306 : tmp44252;
  assign tmp44356 = s3 ? tmp44357 : tmp44255;
  assign tmp44355 = s4 ? tmp44356 : tmp44260;
  assign tmp44354 = s5 ? tmp44355 : tmp44154;
  assign tmp44353 = s6 ? tmp44217 : tmp44354;
  assign tmp44342 = s7 ? tmp44343 : tmp44353;
  assign tmp44363 = s2 ? tmp44325 : tmp44200;
  assign tmp44362 = s3 ? tmp44363 : tmp44202;
  assign tmp44361 = s4 ? tmp44362 : tmp44206;
  assign tmp44360 = s5 ? tmp44361 : tmp44154;
  assign tmp44359 = s6 ? tmp44176 : tmp44360;
  assign tmp44358 = s7 ? tmp44359 : tmp44353;
  assign tmp44341 = s8 ? tmp44342 : tmp44358;
  assign tmp44339 = s9 ? tmp44340 : tmp44341;
  assign tmp44283 = s10 ? tmp44284 : tmp44339;
  assign tmp44367 = s7 ? tmp44287 : tmp44332;
  assign tmp44368 = s7 ? tmp44320 : tmp44332;
  assign tmp44366 = s8 ? tmp44367 : tmp44368;
  assign tmp44365 = s9 ? tmp44340 : tmp44366;
  assign tmp44364 = s10 ? tmp44284 : tmp44365;
  assign tmp44282 = s11 ? tmp44283 : tmp44364;
  assign tmp44378 = ~(s1 ? tmp44093 : tmp44231);
  assign tmp44377 = ~(s2 ? tmp44223 : tmp44378);
  assign tmp44376 = s3 ? tmp44219 : tmp44377;
  assign tmp44380 = s2 ? tmp44234 : tmp44297;
  assign tmp44381 = ~(s2 ? tmp44300 : tmp44244);
  assign tmp44379 = s3 ? tmp44380 : tmp44381;
  assign tmp44375 = s4 ? tmp44376 : tmp44379;
  assign tmp44374 = s6 ? tmp44375 : tmp44248;
  assign tmp44373 = s7 ? tmp43890 : tmp44374;
  assign tmp44372 = s8 ? tmp44373 : tmp44174;
  assign tmp44371 = s9 ? tmp44372 : tmp44214;
  assign tmp44387 = s3 ? tmp44380 : tmp44242;
  assign tmp44386 = s4 ? tmp44376 : tmp44387;
  assign tmp44385 = s6 ? tmp44386 : tmp44248;
  assign tmp44384 = s7 ? tmp44385 : tmp44216;
  assign tmp44383 = s8 ? tmp44384 : tmp44276;
  assign tmp44382 = s9 ? tmp44266 : tmp44383;
  assign tmp44370 = s10 ? tmp44371 : tmp44382;
  assign tmp44391 = s7 ? tmp44374 : tmp44216;
  assign tmp44390 = s8 ? tmp44391 : tmp44276;
  assign tmp44389 = s9 ? tmp44266 : tmp44390;
  assign tmp44388 = s10 ? tmp44371 : tmp44389;
  assign tmp44369 = s11 ? tmp44370 : tmp44388;
  assign tmp44281 = s12 ? tmp44282 : tmp44369;
  assign tmp43884 = s13 ? tmp43885 : tmp44281;
  assign tmp44404 = l1 ? tmp44009 : tmp43934;
  assign tmp44405 = ~(l1 ? 1 : tmp44038);
  assign tmp44403 = ~(s0 ? tmp44404 : tmp44405);
  assign tmp44402 = s1 ? tmp44148 : tmp44403;
  assign tmp44410 = l2 ? tmp43910 : tmp43901;
  assign tmp44409 = l1 ? tmp44410 : tmp43907;
  assign tmp44412 = l2 ? tmp43896 : 0;
  assign tmp44411 = l1 ? tmp44412 : tmp43909;
  assign tmp44408 = s0 ? tmp44409 : tmp44411;
  assign tmp44414 = ~(l1 ? tmp44412 : tmp43909);
  assign tmp44413 = ~(s0 ? tmp44148 : tmp44414);
  assign tmp44407 = s1 ? tmp44408 : tmp44413;
  assign tmp44417 = ~(l2 ? tmp43906 : tmp43902);
  assign tmp44416 = s0 ? tmp44148 : tmp44417;
  assign tmp44418 = ~(s0 ? tmp44411 : tmp44405);
  assign tmp44415 = ~(s1 ? tmp44416 : tmp44418);
  assign tmp44406 = ~(s2 ? tmp44407 : tmp44415);
  assign tmp44401 = s3 ? tmp44402 : tmp44406;
  assign tmp44423 = ~(l1 ? tmp44009 : tmp43936);
  assign tmp44422 = s0 ? tmp44148 : tmp44423;
  assign tmp44424 = s0 ? tmp44148 : tmp44414;
  assign tmp44421 = s1 ? tmp44422 : tmp44424;
  assign tmp44426 = s0 ? tmp44148 : 1;
  assign tmp44427 = ~(l1 ? tmp44009 : tmp44011);
  assign tmp44425 = s1 ? tmp44426 : tmp44427;
  assign tmp44420 = s2 ? tmp44421 : tmp44425;
  assign tmp44429 = s1 ? tmp44404 : tmp44107;
  assign tmp44431 = s0 ? tmp44411 : tmp44110;
  assign tmp44432 = ~(s0 ? tmp44001 : tmp44414);
  assign tmp44430 = s1 ? tmp44431 : tmp44432;
  assign tmp44428 = ~(s2 ? tmp44429 : tmp44430);
  assign tmp44419 = s3 ? tmp44420 : tmp44428;
  assign tmp44400 = s4 ? tmp44401 : tmp44419;
  assign tmp44438 = s0 ? tmp44148 : tmp43949;
  assign tmp44439 = ~(l1 ? tmp44410 : tmp43907);
  assign tmp44437 = s1 ? tmp44438 : tmp44439;
  assign tmp44442 = l2 ? tmp43910 : 0;
  assign tmp44441 = l1 ? tmp44442 : tmp44123;
  assign tmp44440 = ~(s1 ? tmp44441 : tmp44124);
  assign tmp44436 = s2 ? tmp44437 : tmp44440;
  assign tmp44446 = l1 ? tmp44412 : tmp44131;
  assign tmp44445 = ~(s0 ? tmp44446 : tmp44259);
  assign tmp44444 = s1 ? tmp44001 : tmp44445;
  assign tmp44443 = s2 ? tmp44313 : tmp44444;
  assign tmp44435 = s3 ? tmp44436 : tmp44443;
  assign tmp44450 = s0 ? tmp44140 : tmp44405;
  assign tmp44451 = ~(s0 ? tmp43949 : 1);
  assign tmp44449 = s1 ? tmp44450 : tmp44451;
  assign tmp44452 = l1 ? tmp44410 : tmp44123;
  assign tmp44448 = s2 ? tmp44449 : tmp44452;
  assign tmp44447 = ~(s3 ? tmp44448 : tmp44145);
  assign tmp44434 = s4 ? tmp44435 : tmp44447;
  assign tmp44433 = s5 ? tmp44434 : tmp44154;
  assign tmp44399 = s6 ? tmp44400 : tmp44433;
  assign tmp44398 = s7 ? tmp43890 : tmp44399;
  assign tmp44459 = s0 ? tmp44411 : tmp44246;
  assign tmp44458 = s1 ? tmp44459 : tmp44432;
  assign tmp44457 = ~(s2 ? tmp44429 : tmp44458);
  assign tmp44456 = s3 ? tmp44420 : tmp44457;
  assign tmp44455 = s4 ? tmp44401 : tmp44456;
  assign tmp44464 = ~(s1 ? tmp44441 : tmp44253);
  assign tmp44463 = s2 ? tmp44437 : tmp44464;
  assign tmp44466 = ~(s1 ? tmp44001 : tmp44445);
  assign tmp44465 = ~(s2 ? tmp44127 : tmp44466);
  assign tmp44462 = s3 ? tmp44463 : tmp44465;
  assign tmp44461 = s4 ? tmp44462 : tmp44447;
  assign tmp44460 = s5 ? tmp44461 : tmp44154;
  assign tmp44454 = s6 ? tmp44455 : tmp44460;
  assign tmp44453 = s7 ? tmp43890 : tmp44454;
  assign tmp44397 = s8 ? tmp44398 : tmp44453;
  assign tmp44396 = s9 ? tmp44397 : tmp44453;
  assign tmp44468 = s8 ? tmp44453 : tmp43890;
  assign tmp44475 = s2 ? tmp44352 : tmp44444;
  assign tmp44474 = s3 ? tmp44436 : tmp44475;
  assign tmp44473 = s4 ? tmp44474 : tmp44447;
  assign tmp44472 = s5 ? tmp44473 : tmp44154;
  assign tmp44471 = s6 ? tmp44400 : tmp44472;
  assign tmp44470 = s7 ? tmp44471 : tmp44454;
  assign tmp44469 = s8 ? tmp44470 : tmp44454;
  assign tmp44467 = s9 ? tmp44468 : tmp44469;
  assign tmp44395 = s10 ? tmp44396 : tmp44467;
  assign tmp44479 = s7 ? tmp44399 : tmp44454;
  assign tmp44478 = s8 ? tmp44479 : tmp44454;
  assign tmp44477 = s9 ? tmp44468 : tmp44478;
  assign tmp44476 = s10 ? tmp44396 : tmp44477;
  assign tmp44394 = s11 ? tmp44395 : tmp44476;
  assign tmp44489 = l1 ? 1 : tmp43921;
  assign tmp44492 = l2 ? 1 : tmp43901;
  assign tmp44491 = l1 ? tmp44492 : tmp43907;
  assign tmp44493 = ~(l1 ? 1 : tmp43921);
  assign tmp44490 = ~(s0 ? tmp44491 : tmp44493);
  assign tmp44488 = s1 ? tmp44489 : tmp44490;
  assign tmp44498 = l2 ? tmp43906 : tmp43911;
  assign tmp44497 = l1 ? tmp44412 : tmp44498;
  assign tmp44496 = s0 ? tmp44409 : tmp44497;
  assign tmp44500 = ~(l1 ? tmp44412 : tmp44498);
  assign tmp44499 = ~(s0 ? tmp44489 : tmp44500);
  assign tmp44495 = s1 ? tmp44496 : tmp44499;
  assign tmp44502 = s0 ? tmp44489 : tmp44417;
  assign tmp44503 = ~(s0 ? tmp44497 : tmp44493);
  assign tmp44501 = ~(s1 ? tmp44502 : tmp44503);
  assign tmp44494 = ~(s2 ? tmp44495 : tmp44501);
  assign tmp44487 = s3 ? tmp44488 : tmp44494;
  assign tmp44508 = ~(l1 ? tmp44492 : tmp43936);
  assign tmp44507 = s0 ? tmp44489 : tmp44508;
  assign tmp44509 = s0 ? tmp44489 : tmp44500;
  assign tmp44506 = s1 ? tmp44507 : tmp44509;
  assign tmp44511 = s0 ? tmp44489 : 1;
  assign tmp44512 = ~(l1 ? tmp44492 : tmp43944);
  assign tmp44510 = s1 ? tmp44511 : tmp44512;
  assign tmp44505 = s2 ? tmp44506 : tmp44510;
  assign tmp44515 = l1 ? tmp43991 : tmp44045;
  assign tmp44514 = s1 ? tmp44491 : tmp44515;
  assign tmp44519 = ~(l2 ? tmp43906 : tmp43911);
  assign tmp44518 = ~(l1 ? tmp43944 : tmp44519);
  assign tmp44517 = s0 ? tmp44497 : tmp44518;
  assign tmp44522 = l2 ? tmp43897 : 1;
  assign tmp44521 = l1 ? 1 : tmp44522;
  assign tmp44520 = ~(s0 ? tmp44521 : tmp44500);
  assign tmp44516 = s1 ? tmp44517 : tmp44520;
  assign tmp44513 = ~(s2 ? tmp44514 : tmp44516);
  assign tmp44504 = s3 ? tmp44505 : tmp44513;
  assign tmp44486 = s4 ? tmp44487 : tmp44504;
  assign tmp44528 = s0 ? tmp44489 : tmp43949;
  assign tmp44527 = s1 ? tmp44528 : tmp44439;
  assign tmp44531 = l2 ? tmp43906 : tmp43963;
  assign tmp44530 = l1 ? tmp44442 : tmp44531;
  assign tmp44533 = l1 ? tmp43944 : tmp44519;
  assign tmp44532 = ~(s0 ? tmp44533 : 1);
  assign tmp44529 = ~(s1 ? tmp44530 : tmp44532);
  assign tmp44526 = s2 ? tmp44527 : tmp44529;
  assign tmp44536 = l1 ? tmp44129 : tmp43907;
  assign tmp44538 = l2 ? tmp43906 : tmp43897;
  assign tmp44537 = l1 ? tmp44089 : tmp44538;
  assign tmp44535 = s1 ? tmp44536 : tmp44537;
  assign tmp44540 = s0 ? tmp44521 : tmp44001;
  assign tmp44542 = l1 ? tmp44412 : tmp44538;
  assign tmp44544 = l2 ? tmp43897 : tmp43906;
  assign tmp44543 = ~(l1 ? tmp43944 : tmp44544);
  assign tmp44541 = ~(s0 ? tmp44542 : tmp44543);
  assign tmp44539 = ~(s1 ? tmp44540 : tmp44541);
  assign tmp44534 = ~(s2 ? tmp44535 : tmp44539);
  assign tmp44525 = s3 ? tmp44526 : tmp44534;
  assign tmp44549 = l1 ? tmp43955 : tmp44045;
  assign tmp44548 = s0 ? tmp44549 : tmp44493;
  assign tmp44551 = l1 ? tmp43944 : tmp43950;
  assign tmp44550 = ~(s0 ? tmp44551 : tmp44004);
  assign tmp44547 = s1 ? tmp44548 : tmp44550;
  assign tmp44553 = ~(l1 ? tmp44410 : tmp44531);
  assign tmp44552 = ~(s1 ? tmp44010 : tmp44553);
  assign tmp44546 = s2 ? tmp44547 : tmp44552;
  assign tmp44557 = ~(l1 ? tmp44150 : tmp44538);
  assign tmp44556 = s0 ? tmp44489 : tmp44557;
  assign tmp44559 = l1 ? 1 : tmp44544;
  assign tmp44558 = s0 ? tmp44010 : tmp44559;
  assign tmp44555 = s1 ? tmp44556 : tmp44558;
  assign tmp44561 = ~(l1 ? tmp43991 : tmp44045);
  assign tmp44560 = s1 ? tmp44001 : tmp44561;
  assign tmp44554 = ~(s2 ? tmp44555 : tmp44560);
  assign tmp44545 = ~(s3 ? tmp44546 : tmp44554);
  assign tmp44524 = s4 ? tmp44525 : tmp44545;
  assign tmp44566 = s0 ? tmp44537 : tmp44159;
  assign tmp44567 = ~(l1 ? 1 : tmp44005);
  assign tmp44565 = s1 ? tmp44566 : tmp44567;
  assign tmp44564 = s2 ? tmp44565 : tmp44160;
  assign tmp44570 = l1 ? 1 : tmp44005;
  assign tmp44571 = l1 ? 1 : tmp44162;
  assign tmp44569 = s1 ? tmp44570 : tmp44571;
  assign tmp44568 = ~(s2 ? tmp44165 : tmp44569);
  assign tmp44563 = s3 ? tmp44564 : tmp44568;
  assign tmp44574 = s1 ? 1 : tmp44521;
  assign tmp44573 = s2 ? tmp44574 : tmp44489;
  assign tmp44576 = ~(l1 ? tmp44089 : tmp44045);
  assign tmp44575 = s1 ? tmp44001 : tmp44576;
  assign tmp44572 = ~(s3 ? tmp44573 : tmp44575);
  assign tmp44562 = ~(s4 ? tmp44563 : tmp44572);
  assign tmp44523 = s5 ? tmp44524 : tmp44562;
  assign tmp44485 = s6 ? tmp44486 : tmp44523;
  assign tmp44484 = s7 ? tmp43890 : tmp44485;
  assign tmp44583 = l1 ? tmp44009 : tmp43907;
  assign tmp44582 = ~(s0 ? tmp44583 : tmp44493);
  assign tmp44581 = s1 ? tmp44489 : tmp44582;
  assign tmp44580 = s3 ? tmp44581 : tmp44494;
  assign tmp44587 = s0 ? tmp44489 : tmp44423;
  assign tmp44586 = s1 ? tmp44587 : tmp44509;
  assign tmp44589 = ~(l1 ? tmp44009 : tmp43944);
  assign tmp44588 = s1 ? tmp44511 : tmp44589;
  assign tmp44585 = s2 ? tmp44586 : tmp44588;
  assign tmp44591 = s1 ? tmp44583 : tmp44515;
  assign tmp44594 = ~(l1 ? 1 : tmp44519);
  assign tmp44593 = s0 ? tmp44497 : tmp44594;
  assign tmp44592 = s1 ? tmp44593 : tmp44520;
  assign tmp44590 = ~(s2 ? tmp44591 : tmp44592);
  assign tmp44584 = s3 ? tmp44585 : tmp44590;
  assign tmp44579 = s4 ? tmp44580 : tmp44584;
  assign tmp44601 = l1 ? 1 : tmp44519;
  assign tmp44600 = ~(s0 ? tmp44601 : 1);
  assign tmp44599 = ~(s1 ? tmp44530 : tmp44600);
  assign tmp44598 = s2 ? tmp44527 : tmp44599;
  assign tmp44605 = ~(l1 ? 1 : tmp44544);
  assign tmp44604 = ~(s0 ? tmp44542 : tmp44605);
  assign tmp44603 = ~(s1 ? tmp44540 : tmp44604);
  assign tmp44602 = ~(s2 ? tmp44535 : tmp44603);
  assign tmp44597 = s3 ? tmp44598 : tmp44602;
  assign tmp44609 = ~(s0 ? tmp43949 : tmp44570);
  assign tmp44608 = s1 ? tmp44548 : tmp44609;
  assign tmp44610 = l1 ? tmp44410 : tmp44531;
  assign tmp44607 = s2 ? tmp44608 : tmp44610;
  assign tmp44612 = s1 ? tmp44556 : tmp44559;
  assign tmp44611 = ~(s2 ? tmp44612 : tmp44560);
  assign tmp44606 = ~(s3 ? tmp44607 : tmp44611);
  assign tmp44596 = s4 ? tmp44597 : tmp44606;
  assign tmp44595 = s5 ? tmp44596 : tmp44562;
  assign tmp44578 = s6 ? tmp44579 : tmp44595;
  assign tmp44577 = s7 ? tmp43890 : tmp44578;
  assign tmp44483 = s8 ? tmp44484 : tmp44577;
  assign tmp44482 = s9 ? tmp44483 : tmp44577;
  assign tmp44614 = s8 ? tmp44577 : tmp43890;
  assign tmp44620 = ~(s3 ? tmp44546 : tmp44611);
  assign tmp44619 = s4 ? tmp44525 : tmp44620;
  assign tmp44618 = s5 ? tmp44619 : tmp44562;
  assign tmp44617 = s6 ? tmp44486 : tmp44618;
  assign tmp44616 = s7 ? tmp44617 : tmp44578;
  assign tmp44615 = s8 ? tmp44616 : tmp44578;
  assign tmp44613 = s9 ? tmp44614 : tmp44615;
  assign tmp44481 = s10 ? tmp44482 : tmp44613;
  assign tmp44624 = s7 ? tmp44485 : tmp44578;
  assign tmp44623 = s8 ? tmp44624 : tmp44578;
  assign tmp44622 = s9 ? tmp44614 : tmp44623;
  assign tmp44621 = s10 ? tmp44482 : tmp44622;
  assign tmp44480 = s11 ? tmp44481 : tmp44621;
  assign tmp44393 = s12 ? tmp44394 : tmp44480;
  assign tmp44635 = l1 ? tmp44011 : tmp44038;
  assign tmp44637 = l1 ? tmp44492 : tmp43934;
  assign tmp44638 = ~(l1 ? tmp44011 : tmp44038);
  assign tmp44636 = ~(s0 ? tmp44637 : tmp44638);
  assign tmp44634 = s1 ? tmp44635 : tmp44636;
  assign tmp44643 = l2 ? tmp43955 : 0;
  assign tmp44642 = l1 ? tmp44643 : tmp43909;
  assign tmp44641 = s0 ? tmp44491 : tmp44642;
  assign tmp44645 = ~(l1 ? tmp44643 : tmp43909);
  assign tmp44644 = ~(s0 ? tmp44635 : tmp44645);
  assign tmp44640 = s1 ? tmp44641 : tmp44644;
  assign tmp44648 = ~(l1 ? tmp43936 : tmp43907);
  assign tmp44647 = s0 ? tmp44635 : tmp44648;
  assign tmp44649 = ~(s0 ? tmp44642 : tmp44638);
  assign tmp44646 = ~(s1 ? tmp44647 : tmp44649);
  assign tmp44639 = ~(s2 ? tmp44640 : tmp44646);
  assign tmp44633 = s3 ? tmp44634 : tmp44639;
  assign tmp44653 = s0 ? tmp44635 : tmp44508;
  assign tmp44654 = s0 ? tmp44635 : tmp44645;
  assign tmp44652 = s1 ? tmp44653 : tmp44654;
  assign tmp44656 = s0 ? tmp44635 : 1;
  assign tmp44657 = ~(l1 ? tmp44492 : tmp44011);
  assign tmp44655 = s1 ? tmp44656 : tmp44657;
  assign tmp44651 = s2 ? tmp44652 : tmp44655;
  assign tmp44659 = s1 ? tmp44637 : tmp44107;
  assign tmp44662 = ~(l1 ? tmp44011 : tmp44111);
  assign tmp44661 = s0 ? tmp44642 : tmp44662;
  assign tmp44664 = l1 ? tmp44005 : tmp43954;
  assign tmp44663 = ~(s0 ? tmp44664 : tmp44645);
  assign tmp44660 = s1 ? tmp44661 : tmp44663;
  assign tmp44658 = ~(s2 ? tmp44659 : tmp44660);
  assign tmp44650 = s3 ? tmp44651 : tmp44658;
  assign tmp44632 = s4 ? tmp44633 : tmp44650;
  assign tmp44670 = s0 ? tmp44635 : tmp43949;
  assign tmp44671 = ~(l1 ? tmp44492 : tmp43907);
  assign tmp44669 = s1 ? tmp44670 : tmp44671;
  assign tmp44674 = l2 ? 1 : 0;
  assign tmp44673 = l1 ? tmp44674 : tmp44123;
  assign tmp44676 = l1 ? tmp44011 : tmp44111;
  assign tmp44675 = ~(s0 ? tmp44676 : tmp43979);
  assign tmp44672 = ~(s1 ? tmp44673 : tmp44675);
  assign tmp44668 = s2 ? tmp44669 : tmp44672;
  assign tmp44680 = l2 ? 1 : tmp43900;
  assign tmp44679 = l1 ? tmp44680 : tmp43934;
  assign tmp44682 = l2 ? tmp43955 : tmp43896;
  assign tmp44681 = l1 ? tmp44682 : tmp44131;
  assign tmp44678 = s1 ? tmp44679 : tmp44681;
  assign tmp44684 = s0 ? tmp44664 : tmp44001;
  assign tmp44686 = l1 ? tmp44643 : tmp44131;
  assign tmp44687 = ~(l1 ? tmp44011 : tmp44135);
  assign tmp44685 = ~(s0 ? tmp44686 : tmp44687);
  assign tmp44683 = ~(s1 ? tmp44684 : tmp44685);
  assign tmp44677 = ~(s2 ? tmp44678 : tmp44683);
  assign tmp44667 = s3 ? tmp44668 : tmp44677;
  assign tmp44691 = s0 ? tmp44140 : tmp44638;
  assign tmp44692 = ~(s0 ? tmp44551 : tmp43979);
  assign tmp44690 = s1 ? tmp44691 : tmp44692;
  assign tmp44693 = l1 ? tmp44492 : tmp44123;
  assign tmp44689 = s2 ? tmp44690 : tmp44693;
  assign tmp44698 = l2 ? tmp43955 : tmp43900;
  assign tmp44697 = ~(l1 ? tmp44698 : tmp44131);
  assign tmp44696 = s0 ? tmp44037 : tmp44697;
  assign tmp44699 = l1 ? tmp44005 : tmp44135;
  assign tmp44695 = s1 ? tmp44696 : tmp44699;
  assign tmp44694 = ~(s2 ? tmp44695 : tmp44152);
  assign tmp44688 = ~(s3 ? tmp44689 : tmp44694);
  assign tmp44666 = s4 ? tmp44667 : tmp44688;
  assign tmp44704 = s0 ? tmp44681 : tmp44159;
  assign tmp44705 = ~(l1 ? tmp44005 : 1);
  assign tmp44703 = s1 ? tmp44704 : tmp44705;
  assign tmp44707 = s0 ? tmp44036 : tmp44037;
  assign tmp44706 = s1 ? tmp43943 : tmp44707;
  assign tmp44702 = s2 ? tmp44703 : tmp44706;
  assign tmp44710 = s0 ? tmp44042 : 0;
  assign tmp44711 = l1 ? tmp44045 : tmp43992;
  assign tmp44709 = s1 ? tmp44710 : tmp44711;
  assign tmp44712 = ~(s1 ? 1 : tmp44042);
  assign tmp44708 = s2 ? tmp44709 : tmp44712;
  assign tmp44701 = s3 ? tmp44702 : tmp44708;
  assign tmp44716 = l1 ? tmp44005 : 1;
  assign tmp44715 = s1 ? tmp44716 : tmp44664;
  assign tmp44718 = ~(s0 ? tmp44037 : tmp44042);
  assign tmp44717 = s1 ? tmp44037 : tmp44718;
  assign tmp44714 = s2 ? tmp44715 : tmp44717;
  assign tmp44720 = ~(l1 ? tmp44682 : tmp43962);
  assign tmp44719 = s1 ? tmp44664 : tmp44720;
  assign tmp44713 = ~(s3 ? tmp44714 : tmp44719);
  assign tmp44700 = ~(s4 ? tmp44701 : tmp44713);
  assign tmp44665 = s5 ? tmp44666 : tmp44700;
  assign tmp44631 = s6 ? tmp44632 : tmp44665;
  assign tmp44630 = s7 ? tmp43890 : tmp44631;
  assign tmp44727 = ~(l1 ? tmp44005 : tmp44038);
  assign tmp44726 = ~(s0 ? tmp44404 : tmp44727);
  assign tmp44725 = s1 ? tmp44037 : tmp44726;
  assign tmp44732 = l2 ? tmp43900 : 0;
  assign tmp44731 = l1 ? tmp44732 : tmp43909;
  assign tmp44730 = s0 ? tmp44583 : tmp44731;
  assign tmp44734 = ~(l1 ? tmp44732 : tmp43909);
  assign tmp44733 = ~(s0 ? tmp44037 : tmp44734);
  assign tmp44729 = s1 ? tmp44730 : tmp44733;
  assign tmp44736 = s0 ? tmp44037 : tmp44417;
  assign tmp44737 = ~(s0 ? tmp44731 : tmp44727);
  assign tmp44735 = ~(s1 ? tmp44736 : tmp44737);
  assign tmp44728 = ~(s2 ? tmp44729 : tmp44735);
  assign tmp44724 = s3 ? tmp44725 : tmp44728;
  assign tmp44741 = s0 ? tmp44037 : tmp44423;
  assign tmp44742 = s0 ? tmp44037 : tmp44734;
  assign tmp44740 = s1 ? tmp44741 : tmp44742;
  assign tmp44744 = s0 ? tmp44037 : 1;
  assign tmp44743 = s1 ? tmp44744 : tmp44427;
  assign tmp44739 = s2 ? tmp44740 : tmp44743;
  assign tmp44748 = ~(l1 ? tmp44005 : tmp44111);
  assign tmp44747 = s0 ? tmp44731 : tmp44748;
  assign tmp44749 = ~(s0 ? tmp44664 : tmp44734);
  assign tmp44746 = s1 ? tmp44747 : tmp44749;
  assign tmp44745 = ~(s2 ? tmp44429 : tmp44746);
  assign tmp44738 = s3 ? tmp44739 : tmp44745;
  assign tmp44723 = s4 ? tmp44724 : tmp44738;
  assign tmp44755 = s0 ? tmp44037 : tmp43949;
  assign tmp44756 = ~(l1 ? tmp44009 : tmp43907);
  assign tmp44754 = s1 ? tmp44755 : tmp44756;
  assign tmp44759 = l2 ? tmp43906 : 0;
  assign tmp44758 = l1 ? tmp44759 : tmp44123;
  assign tmp44761 = l1 ? tmp44005 : tmp44111;
  assign tmp44760 = ~(s0 ? tmp44761 : 1);
  assign tmp44757 = ~(s1 ? tmp44758 : tmp44760);
  assign tmp44753 = s2 ? tmp44754 : tmp44757;
  assign tmp44765 = l2 ? tmp43906 : tmp43900;
  assign tmp44764 = l1 ? tmp44765 : tmp43934;
  assign tmp44763 = s1 ? tmp44764 : tmp44681;
  assign tmp44768 = l1 ? tmp44732 : tmp44131;
  assign tmp44769 = ~(l1 ? tmp44005 : tmp44135);
  assign tmp44767 = ~(s0 ? tmp44768 : tmp44769);
  assign tmp44766 = ~(s1 ? tmp44684 : tmp44767);
  assign tmp44762 = ~(s2 ? tmp44763 : tmp44766);
  assign tmp44752 = s3 ? tmp44753 : tmp44762;
  assign tmp44773 = s0 ? tmp44140 : tmp44727;
  assign tmp44772 = s1 ? tmp44773 : tmp44451;
  assign tmp44774 = l1 ? tmp44009 : tmp44123;
  assign tmp44771 = s2 ? tmp44772 : tmp44774;
  assign tmp44778 = ~(l1 ? tmp43900 : tmp44131);
  assign tmp44777 = s0 ? tmp44037 : tmp44778;
  assign tmp44776 = s1 ? tmp44777 : tmp44699;
  assign tmp44775 = ~(s2 ? tmp44776 : tmp44152);
  assign tmp44770 = ~(s3 ? tmp44771 : tmp44775);
  assign tmp44751 = s4 ? tmp44752 : tmp44770;
  assign tmp44782 = s1 ? tmp43943 : tmp44036;
  assign tmp44781 = s2 ? tmp44703 : tmp44782;
  assign tmp44780 = s3 ? tmp44781 : tmp44708;
  assign tmp44786 = ~(l1 ? tmp44005 : tmp43905);
  assign tmp44785 = s1 ? tmp44037 : tmp44786;
  assign tmp44784 = s2 ? tmp44715 : tmp44785;
  assign tmp44783 = ~(s3 ? tmp44784 : tmp44719);
  assign tmp44779 = ~(s4 ? tmp44780 : tmp44783);
  assign tmp44750 = s5 ? tmp44751 : tmp44779;
  assign tmp44722 = s6 ? tmp44723 : tmp44750;
  assign tmp44721 = s7 ? tmp43890 : tmp44722;
  assign tmp44629 = s8 ? tmp44630 : tmp44721;
  assign tmp44628 = s9 ? tmp44629 : tmp44721;
  assign tmp44788 = s8 ? tmp44721 : tmp43890;
  assign tmp44795 = s2 ? tmp44715 : tmp44037;
  assign tmp44794 = ~(s3 ? tmp44795 : tmp44719);
  assign tmp44793 = ~(s4 ? tmp44701 : tmp44794);
  assign tmp44792 = s5 ? tmp44666 : tmp44793;
  assign tmp44791 = s6 ? tmp44632 : tmp44792;
  assign tmp44798 = ~(s4 ? tmp44780 : tmp44794);
  assign tmp44797 = s5 ? tmp44751 : tmp44798;
  assign tmp44796 = s6 ? tmp44723 : tmp44797;
  assign tmp44790 = s7 ? tmp44791 : tmp44796;
  assign tmp44789 = s8 ? tmp44790 : tmp44796;
  assign tmp44787 = s9 ? tmp44788 : tmp44789;
  assign tmp44627 = s10 ? tmp44628 : tmp44787;
  assign tmp44802 = s7 ? tmp44631 : tmp44722;
  assign tmp44801 = s8 ? tmp44802 : tmp44722;
  assign tmp44800 = s9 ? tmp44788 : tmp44801;
  assign tmp44799 = s10 ? tmp44628 : tmp44800;
  assign tmp44626 = s11 ? tmp44627 : tmp44799;
  assign tmp44813 = s0 ? tmp44635 : tmp44417;
  assign tmp44812 = ~(s1 ? tmp44813 : tmp44649);
  assign tmp44811 = ~(s2 ? tmp44640 : tmp44812);
  assign tmp44810 = s3 ? tmp44634 : tmp44811;
  assign tmp44809 = s4 ? tmp44810 : tmp44650;
  assign tmp44819 = ~(s0 ? tmp44676 : 1);
  assign tmp44818 = ~(s1 ? tmp44673 : tmp44819);
  assign tmp44817 = s2 ? tmp44669 : tmp44818;
  assign tmp44816 = s3 ? tmp44817 : tmp44677;
  assign tmp44815 = s4 ? tmp44816 : tmp44688;
  assign tmp44814 = s5 ? tmp44815 : tmp44779;
  assign tmp44808 = s6 ? tmp44809 : tmp44814;
  assign tmp44807 = s7 ? tmp43890 : tmp44808;
  assign tmp44806 = s8 ? tmp44807 : tmp44721;
  assign tmp44805 = s9 ? tmp44806 : tmp44721;
  assign tmp44824 = s5 ? tmp44815 : tmp44798;
  assign tmp44823 = s6 ? tmp44809 : tmp44824;
  assign tmp44822 = s7 ? tmp44823 : tmp44796;
  assign tmp44821 = s8 ? tmp44822 : tmp44796;
  assign tmp44820 = s9 ? tmp44788 : tmp44821;
  assign tmp44804 = s10 ? tmp44805 : tmp44820;
  assign tmp44828 = s7 ? tmp44808 : tmp44722;
  assign tmp44827 = s8 ? tmp44828 : tmp44722;
  assign tmp44826 = s9 ? tmp44788 : tmp44827;
  assign tmp44825 = s10 ? tmp44805 : tmp44826;
  assign tmp44803 = s11 ? tmp44804 : tmp44825;
  assign tmp44625 = s12 ? tmp44626 : tmp44803;
  assign tmp44392 = s13 ? tmp44393 : tmp44625;
  assign tmp43883 = s14 ? tmp43884 : tmp44392;
  assign tmp44839 = l1 ? tmp43955 : tmp44038;
  assign tmp44841 = ~(l1 ? tmp43992 : tmp44038);
  assign tmp44840 = ~(s0 ? tmp44404 : tmp44841);
  assign tmp44838 = s1 ? tmp44839 : tmp44840;
  assign tmp44847 = ~(l3 ? tmp43897 : 1);
  assign tmp44846 = l2 ? tmp43910 : tmp44847;
  assign tmp44845 = l1 ? tmp44846 : tmp43928;
  assign tmp44844 = s0 ? tmp44409 : tmp44845;
  assign tmp44849 = l1 ? tmp43992 : tmp44038;
  assign tmp44850 = ~(l1 ? tmp44846 : tmp43928);
  assign tmp44848 = ~(s0 ? tmp44849 : tmp44850);
  assign tmp44843 = s1 ? tmp44844 : tmp44848;
  assign tmp44852 = s0 ? tmp44849 : tmp44417;
  assign tmp44854 = ~(l1 ? tmp43955 : tmp44038);
  assign tmp44853 = ~(s0 ? tmp44845 : tmp44854);
  assign tmp44851 = ~(s1 ? tmp44852 : tmp44853);
  assign tmp44842 = ~(s2 ? tmp44843 : tmp44851);
  assign tmp44837 = s3 ? tmp44838 : tmp44842;
  assign tmp44858 = s0 ? tmp44839 : tmp44850;
  assign tmp44857 = s1 ? tmp44422 : tmp44858;
  assign tmp44860 = s0 ? tmp44839 : 1;
  assign tmp44859 = s1 ? tmp44860 : tmp44427;
  assign tmp44856 = s2 ? tmp44857 : tmp44859;
  assign tmp44863 = l1 ? tmp44044 : tmp43897;
  assign tmp44862 = s1 ? tmp44404 : tmp44863;
  assign tmp44865 = s0 ? tmp44845 : tmp44854;
  assign tmp44866 = ~(s0 ? tmp44159 : tmp44850);
  assign tmp44864 = s1 ? tmp44865 : tmp44866;
  assign tmp44861 = ~(s2 ? tmp44862 : tmp44864);
  assign tmp44855 = s3 ? tmp44856 : tmp44861;
  assign tmp44836 = s4 ? tmp44837 : tmp44855;
  assign tmp44872 = s0 ? tmp44849 : tmp43949;
  assign tmp44871 = s1 ? tmp44872 : tmp44439;
  assign tmp44874 = l1 ? tmp44846 : tmp44123;
  assign tmp44875 = ~(s0 ? tmp44839 : 1);
  assign tmp44873 = ~(s1 ? tmp44874 : tmp44875);
  assign tmp44870 = s2 ? tmp44871 : tmp44873;
  assign tmp44878 = l1 ? tmp44087 : tmp43934;
  assign tmp44879 = l1 ? tmp44054 : tmp43959;
  assign tmp44877 = s1 ? tmp44878 : tmp44879;
  assign tmp44882 = l1 ? tmp44846 : tmp43959;
  assign tmp44883 = ~(l1 ? tmp43955 : tmp43905);
  assign tmp44881 = ~(s0 ? tmp44882 : tmp44883);
  assign tmp44880 = ~(s1 ? tmp44159 : tmp44881);
  assign tmp44876 = ~(s2 ? tmp44877 : tmp44880);
  assign tmp44869 = s3 ? tmp44870 : tmp44876;
  assign tmp44888 = l1 ? 1 : tmp43897;
  assign tmp44887 = s0 ? tmp44888 : tmp44854;
  assign tmp44886 = s1 ? tmp44887 : tmp44451;
  assign tmp44885 = s2 ? tmp44886 : tmp44452;
  assign tmp44892 = ~(l1 ? tmp44087 : tmp44131);
  assign tmp44891 = s0 ? tmp44148 : tmp44892;
  assign tmp44893 = l1 ? tmp43955 : tmp43905;
  assign tmp44890 = s1 ? tmp44891 : tmp44893;
  assign tmp44895 = l1 ? tmp43954 : 1;
  assign tmp44896 = ~(l1 ? tmp44044 : tmp43897);
  assign tmp44894 = s1 ? tmp44895 : tmp44896;
  assign tmp44889 = ~(s2 ? tmp44890 : tmp44894);
  assign tmp44884 = ~(s3 ? tmp44885 : tmp44889);
  assign tmp44868 = s4 ? tmp44869 : tmp44884;
  assign tmp44901 = s0 ? tmp44879 : tmp44001;
  assign tmp44903 = ~(l1 ? tmp43992 : 1);
  assign tmp44902 = s0 ? tmp44001 : tmp44903;
  assign tmp44900 = s1 ? tmp44901 : tmp44902;
  assign tmp44899 = s2 ? tmp44900 : tmp44160;
  assign tmp44906 = ~(l1 ? tmp44044 : tmp43955);
  assign tmp44905 = s1 ? 1 : tmp44906;
  assign tmp44907 = s1 ? tmp44159 : tmp44168;
  assign tmp44904 = ~(s2 ? tmp44905 : tmp44907);
  assign tmp44898 = s3 ? tmp44899 : tmp44904;
  assign tmp44911 = l1 ? tmp43992 : 1;
  assign tmp44910 = s1 ? tmp44911 : tmp44159;
  assign tmp44912 = ~(s0 ? tmp44001 : tmp44841);
  assign tmp44909 = s2 ? tmp44910 : tmp44912;
  assign tmp44914 = ~(l1 ? tmp44054 : tmp43962);
  assign tmp44913 = s1 ? tmp44911 : tmp44914;
  assign tmp44908 = ~(s3 ? tmp44909 : tmp44913);
  assign tmp44897 = ~(s4 ? tmp44898 : tmp44908);
  assign tmp44867 = s5 ? tmp44868 : tmp44897;
  assign tmp44835 = s6 ? tmp44836 : tmp44867;
  assign tmp44834 = s7 ? tmp43890 : tmp44835;
  assign tmp44916 = s8 ? tmp44834 : tmp43890;
  assign tmp44921 = s2 ? tmp44910 : tmp44849;
  assign tmp44920 = ~(s3 ? tmp44921 : tmp44913);
  assign tmp44919 = ~(s4 ? tmp44898 : tmp44920);
  assign tmp44918 = s5 ? tmp44868 : tmp44919;
  assign tmp44917 = s6 ? tmp44836 : tmp44918;
  assign tmp44915 = s9 ? tmp44916 : tmp44917;
  assign tmp44833 = s10 ? tmp44834 : tmp44915;
  assign tmp44923 = s9 ? tmp44916 : tmp44835;
  assign tmp44922 = s10 ? tmp44834 : tmp44923;
  assign tmp44832 = s11 ? tmp44833 : tmp44922;
  assign tmp44933 = ~(l3 ? tmp43897 : tmp43901);
  assign tmp44932 = ~(l2 ? tmp43896 : tmp44933);
  assign tmp44931 = l1 ? tmp43954 : tmp44932;
  assign tmp44930 = s1 ? tmp44931 : tmp44403;
  assign tmp44938 = l2 ? tmp43896 : tmp44933;
  assign tmp44937 = l1 ? tmp44442 : tmp44938;
  assign tmp44936 = s0 ? tmp44409 : tmp44937;
  assign tmp44940 = ~(l1 ? tmp44442 : tmp44938);
  assign tmp44939 = ~(s0 ? tmp44148 : tmp44940);
  assign tmp44935 = s1 ? tmp44936 : tmp44939;
  assign tmp44943 = ~(l1 ? tmp43954 : tmp44932);
  assign tmp44942 = ~(s0 ? tmp44937 : tmp44943);
  assign tmp44941 = ~(s1 ? tmp44416 : tmp44942);
  assign tmp44934 = ~(s2 ? tmp44935 : tmp44941);
  assign tmp44929 = s3 ? tmp44930 : tmp44934;
  assign tmp44947 = s0 ? tmp44931 : tmp44940;
  assign tmp44946 = s1 ? tmp44422 : tmp44947;
  assign tmp44949 = s0 ? tmp44931 : 1;
  assign tmp44948 = s1 ? tmp44949 : tmp44427;
  assign tmp44945 = s2 ? tmp44946 : tmp44948;
  assign tmp44953 = l2 ? tmp43897 : tmp43963;
  assign tmp44952 = l1 ? tmp44045 : tmp44953;
  assign tmp44951 = s1 ? tmp44404 : tmp44952;
  assign tmp44955 = s0 ? tmp44937 : tmp44943;
  assign tmp44956 = ~(s0 ? tmp44021 : tmp44940);
  assign tmp44954 = s1 ? tmp44955 : tmp44956;
  assign tmp44950 = ~(s2 ? tmp44951 : tmp44954);
  assign tmp44944 = s3 ? tmp44945 : tmp44950;
  assign tmp44928 = s4 ? tmp44929 : tmp44944;
  assign tmp44962 = ~(s0 ? tmp44931 : 1);
  assign tmp44961 = ~(s1 ? tmp44441 : tmp44962);
  assign tmp44960 = s2 ? tmp44437 : tmp44961;
  assign tmp44966 = l2 ? tmp43896 : tmp43963;
  assign tmp44965 = l1 ? tmp43996 : tmp44966;
  assign tmp44964 = s1 ? tmp44128 : tmp44965;
  assign tmp44969 = l1 ? tmp44442 : tmp44966;
  assign tmp44970 = ~(l1 ? tmp43954 : tmp44680);
  assign tmp44968 = ~(s0 ? tmp44969 : tmp44970);
  assign tmp44967 = ~(s1 ? tmp44021 : tmp44968);
  assign tmp44963 = ~(s2 ? tmp44964 : tmp44967);
  assign tmp44959 = s3 ? tmp44960 : tmp44963;
  assign tmp44975 = l1 ? tmp43992 : tmp44953;
  assign tmp44974 = s0 ? tmp44975 : tmp44943;
  assign tmp44973 = s1 ? tmp44974 : tmp44451;
  assign tmp44972 = s2 ? tmp44973 : tmp44452;
  assign tmp44979 = ~(l1 ? tmp44129 : tmp44123);
  assign tmp44978 = s0 ? tmp44148 : tmp44979;
  assign tmp44980 = l1 ? tmp43954 : tmp44680;
  assign tmp44977 = s1 ? tmp44978 : tmp44980;
  assign tmp44982 = ~(s0 ? tmp44952 : tmp44023);
  assign tmp44981 = s1 ? tmp44021 : tmp44982;
  assign tmp44976 = ~(s2 ? tmp44977 : tmp44981);
  assign tmp44971 = ~(s3 ? tmp44972 : tmp44976);
  assign tmp44958 = s4 ? tmp44959 : tmp44971;
  assign tmp44988 = l1 ? tmp43992 : tmp43954;
  assign tmp44987 = s0 ? tmp44965 : tmp44988;
  assign tmp44986 = s1 ? tmp44987 : 0;
  assign tmp44985 = s2 ? tmp44986 : tmp44160;
  assign tmp44991 = l1 ? 1 : tmp43992;
  assign tmp44992 = ~(l1 ? tmp44045 : tmp43954);
  assign tmp44990 = s1 ? tmp44991 : tmp44992;
  assign tmp44993 = s1 ? tmp44021 : tmp44168;
  assign tmp44989 = ~(s2 ? tmp44990 : tmp44993);
  assign tmp44984 = s3 ? tmp44985 : tmp44989;
  assign tmp44996 = s1 ? 1 : tmp44021;
  assign tmp44995 = s2 ? tmp44996 : tmp44148;
  assign tmp44998 = ~(l1 ? tmp43996 : tmp43963);
  assign tmp44997 = s1 ? tmp44991 : tmp44998;
  assign tmp44994 = ~(s3 ? tmp44995 : tmp44997);
  assign tmp44983 = ~(s4 ? tmp44984 : tmp44994);
  assign tmp44957 = s5 ? tmp44958 : tmp44983;
  assign tmp44927 = s6 ? tmp44928 : tmp44957;
  assign tmp44926 = s7 ? tmp43890 : tmp44927;
  assign tmp45000 = s8 ? tmp44926 : tmp43890;
  assign tmp45007 = ~(l1 ? tmp44045 : tmp44953);
  assign tmp45006 = s1 ? tmp44021 : tmp45007;
  assign tmp45005 = ~(s2 ? tmp44977 : tmp45006);
  assign tmp45004 = ~(s3 ? tmp44972 : tmp45005);
  assign tmp45003 = s4 ? tmp44959 : tmp45004;
  assign tmp45002 = s5 ? tmp45003 : tmp44983;
  assign tmp45001 = s6 ? tmp44928 : tmp45002;
  assign tmp44999 = s9 ? tmp45000 : tmp45001;
  assign tmp44925 = s10 ? tmp44926 : tmp44999;
  assign tmp45009 = s9 ? tmp45000 : tmp44927;
  assign tmp45008 = s10 ? tmp44926 : tmp45009;
  assign tmp44924 = s11 ? tmp44925 : tmp45008;
  assign tmp44831 = s12 ? tmp44832 : tmp44924;
  assign tmp45018 = l1 ? tmp43955 : tmp43899;
  assign tmp45020 = ~(l1 ? tmp43992 : tmp43912);
  assign tmp45019 = ~(s0 ? tmp44583 : tmp45020);
  assign tmp45017 = s1 ? tmp45018 : tmp45019;
  assign tmp45024 = l1 ? tmp44846 : tmp43907;
  assign tmp45023 = s0 ? tmp44409 : tmp45024;
  assign tmp45026 = l1 ? tmp43992 : tmp43921;
  assign tmp45027 = ~(l1 ? tmp44846 : tmp43907);
  assign tmp45025 = ~(s0 ? tmp45026 : tmp45027);
  assign tmp45022 = s1 ? tmp45023 : tmp45025;
  assign tmp45029 = s0 ? tmp45026 : tmp44417;
  assign tmp45031 = ~(l1 ? tmp43955 : tmp43899);
  assign tmp45030 = ~(s0 ? tmp45024 : tmp45031);
  assign tmp45028 = ~(s1 ? tmp45029 : tmp45030);
  assign tmp45021 = ~(s2 ? tmp45022 : tmp45028);
  assign tmp45016 = s3 ? tmp45017 : tmp45021;
  assign tmp45036 = l1 ? 1 : tmp43912;
  assign tmp45035 = s0 ? tmp45036 : tmp44423;
  assign tmp45037 = s0 ? tmp45018 : tmp45027;
  assign tmp45034 = s1 ? tmp45035 : tmp45037;
  assign tmp45039 = s0 ? tmp45018 : 1;
  assign tmp45038 = s1 ? tmp45039 : tmp44589;
  assign tmp45033 = s2 ? tmp45034 : tmp45038;
  assign tmp45042 = l1 ? tmp44044 : 1;
  assign tmp45041 = s1 ? tmp44583 : tmp45042;
  assign tmp45045 = ~(l1 ? tmp43955 : tmp44417);
  assign tmp45044 = s0 ? tmp45024 : tmp45045;
  assign tmp45047 = l1 ? tmp43955 : tmp43897;
  assign tmp45046 = ~(s0 ? tmp45047 : tmp45027);
  assign tmp45043 = s1 ? tmp45044 : tmp45046;
  assign tmp45040 = ~(s2 ? tmp45041 : tmp45043);
  assign tmp45032 = s3 ? tmp45033 : tmp45040;
  assign tmp45015 = s4 ? tmp45016 : tmp45032;
  assign tmp45054 = l1 ? tmp43992 : tmp43912;
  assign tmp45053 = s0 ? tmp45054 : tmp43949;
  assign tmp45052 = s1 ? tmp45053 : tmp44439;
  assign tmp45056 = l1 ? tmp44846 : tmp43944;
  assign tmp45058 = l1 ? tmp43955 : tmp44417;
  assign tmp45057 = ~(s0 ? tmp45058 : 1);
  assign tmp45055 = ~(s1 ? tmp45056 : tmp45057);
  assign tmp45051 = s2 ? tmp45052 : tmp45055;
  assign tmp45061 = l1 ? tmp44054 : tmp43944;
  assign tmp45060 = s1 ? tmp44086 : tmp45061;
  assign tmp45063 = s0 ? tmp45047 : tmp43955;
  assign tmp45065 = ~(l1 ? tmp43955 : tmp44089);
  assign tmp45064 = ~(s0 ? tmp45056 : tmp45065);
  assign tmp45062 = ~(s1 ? tmp45063 : tmp45064);
  assign tmp45059 = ~(s2 ? tmp45060 : tmp45062);
  assign tmp45050 = s3 ? tmp45051 : tmp45059;
  assign tmp45069 = s0 ? 1 : tmp45031;
  assign tmp45068 = s1 ? tmp45069 : tmp44609;
  assign tmp45070 = l1 ? tmp44410 : tmp43944;
  assign tmp45067 = s2 ? tmp45068 : tmp45070;
  assign tmp45074 = ~(l1 ? tmp44087 : tmp43944);
  assign tmp45073 = s0 ? tmp45036 : tmp45074;
  assign tmp45075 = l1 ? tmp43955 : tmp44089;
  assign tmp45072 = s1 ? tmp45073 : tmp45075;
  assign tmp45077 = l1 ? tmp43954 : tmp43955;
  assign tmp45078 = ~(l1 ? tmp44044 : 1);
  assign tmp45076 = s1 ? tmp45077 : tmp45078;
  assign tmp45071 = ~(s2 ? tmp45072 : tmp45076);
  assign tmp45066 = ~(s3 ? tmp45067 : tmp45071);
  assign tmp45049 = s4 ? tmp45050 : tmp45066;
  assign tmp45083 = s0 ? tmp45061 : 1;
  assign tmp45084 = ~(l1 ? tmp43992 : tmp44005);
  assign tmp45082 = s1 ? tmp45083 : tmp45084;
  assign tmp45081 = s2 ? tmp45082 : tmp44160;
  assign tmp45087 = l1 ? 1 : tmp44045;
  assign tmp45086 = s1 ? tmp45087 : tmp45078;
  assign tmp45090 = l1 ? 1 : tmp44054;
  assign tmp45089 = s0 ? tmp44052 : tmp45090;
  assign tmp45088 = s1 ? tmp44140 : tmp45089;
  assign tmp45085 = ~(s2 ? tmp45086 : tmp45088);
  assign tmp45080 = s3 ? tmp45081 : tmp45085;
  assign tmp45094 = l1 ? tmp43992 : tmp44044;
  assign tmp45093 = s1 ? tmp45094 : tmp45047;
  assign tmp45092 = s2 ? tmp45093 : tmp45054;
  assign tmp45097 = l1 ? tmp43992 : tmp43991;
  assign tmp45098 = ~(l1 ? tmp44054 : 1);
  assign tmp45096 = s1 ? tmp45097 : tmp45098;
  assign tmp45095 = s2 ? tmp45096 : tmp44052;
  assign tmp45091 = ~(s3 ? tmp45092 : tmp45095);
  assign tmp45079 = ~(s4 ? tmp45080 : tmp45091);
  assign tmp45048 = s5 ? tmp45049 : tmp45079;
  assign tmp45014 = s6 ? tmp45015 : tmp45048;
  assign tmp45013 = s7 ? tmp43890 : tmp45014;
  assign tmp45100 = s8 ? tmp45013 : tmp43890;
  assign tmp45104 = ~(s3 ? tmp45092 : tmp45096);
  assign tmp45103 = ~(s4 ? tmp45080 : tmp45104);
  assign tmp45102 = s5 ? tmp45049 : tmp45103;
  assign tmp45101 = s6 ? tmp45015 : tmp45102;
  assign tmp45099 = s9 ? tmp45100 : tmp45101;
  assign tmp45012 = s10 ? tmp45013 : tmp45099;
  assign tmp45106 = s9 ? tmp45100 : tmp45014;
  assign tmp45105 = s10 ? tmp45013 : tmp45106;
  assign tmp45011 = s11 ? tmp45012 : tmp45105;
  assign tmp45114 = l1 ? tmp43992 : tmp44932;
  assign tmp45116 = ~(l1 ? tmp44045 : tmp44038);
  assign tmp45115 = ~(s0 ? tmp44404 : tmp45116);
  assign tmp45113 = s1 ? tmp45114 : tmp45115;
  assign tmp45121 = l2 ? tmp43896 : tmp43901;
  assign tmp45120 = l1 ? tmp45121 : tmp44938;
  assign tmp45119 = s0 ? tmp44409 : tmp45120;
  assign tmp45123 = ~(l1 ? tmp45121 : tmp44938);
  assign tmp45122 = ~(s0 ? tmp44849 : tmp45123);
  assign tmp45118 = s1 ? tmp45119 : tmp45122;
  assign tmp45126 = ~(l1 ? tmp44045 : tmp44932);
  assign tmp45125 = ~(s0 ? tmp45120 : tmp45126);
  assign tmp45124 = ~(s1 ? tmp44852 : tmp45125);
  assign tmp45117 = ~(s2 ? tmp45118 : tmp45124);
  assign tmp45112 = s3 ? tmp45113 : tmp45117;
  assign tmp45131 = l1 ? tmp44045 : tmp44932;
  assign tmp45130 = s0 ? tmp45131 : tmp45123;
  assign tmp45129 = s1 ? tmp44422 : tmp45130;
  assign tmp45133 = s0 ? tmp45114 : 1;
  assign tmp45132 = s1 ? tmp45133 : tmp44427;
  assign tmp45128 = s2 ? tmp45129 : tmp45132;
  assign tmp45136 = l1 ? tmp43954 : tmp44953;
  assign tmp45135 = s1 ? tmp44404 : tmp45136;
  assign tmp45138 = s0 ? tmp45120 : tmp45126;
  assign tmp45139 = ~(s0 ? tmp44711 : tmp45123);
  assign tmp45137 = s1 ? tmp45138 : tmp45139;
  assign tmp45134 = ~(s2 ? tmp45135 : tmp45137);
  assign tmp45127 = s3 ? tmp45128 : tmp45134;
  assign tmp45111 = s4 ? tmp45112 : tmp45127;
  assign tmp45146 = l1 ? tmp44045 : tmp44038;
  assign tmp45145 = s0 ? tmp45146 : tmp43949;
  assign tmp45144 = s1 ? tmp45145 : tmp44439;
  assign tmp45148 = ~(s0 ? tmp45131 : 1);
  assign tmp45147 = ~(s1 ? tmp44452 : tmp45148);
  assign tmp45143 = s2 ? tmp45144 : tmp45147;
  assign tmp45151 = l1 ? tmp44544 : tmp44966;
  assign tmp45150 = s1 ? tmp44878 : tmp45151;
  assign tmp45154 = l1 ? tmp45121 : tmp44966;
  assign tmp45155 = ~(l1 ? tmp44045 : tmp44680);
  assign tmp45153 = ~(s0 ? tmp45154 : tmp45155);
  assign tmp45152 = ~(s1 ? tmp44711 : tmp45153);
  assign tmp45149 = ~(s2 ? tmp45150 : tmp45152);
  assign tmp45142 = s3 ? tmp45143 : tmp45149;
  assign tmp45159 = s0 ? tmp45136 : tmp45126;
  assign tmp45158 = s1 ? tmp45159 : tmp44451;
  assign tmp45157 = s2 ? tmp45158 : tmp44452;
  assign tmp45164 = l2 ? tmp43896 : tmp43906;
  assign tmp45163 = ~(l1 ? tmp45164 : tmp44123);
  assign tmp45162 = s0 ? tmp44148 : tmp45163;
  assign tmp45165 = l1 ? tmp44045 : tmp44680;
  assign tmp45161 = s1 ? tmp45162 : tmp45165;
  assign tmp45167 = ~(l1 ? tmp43954 : tmp44953);
  assign tmp45166 = s1 ? tmp44991 : tmp45167;
  assign tmp45160 = ~(s2 ? tmp45161 : tmp45166);
  assign tmp45156 = ~(s3 ? tmp45157 : tmp45160);
  assign tmp45141 = s4 ? tmp45142 : tmp45156;
  assign tmp45172 = s0 ? tmp45151 : tmp43954;
  assign tmp45171 = s1 ? tmp45172 : tmp44903;
  assign tmp45170 = s2 ? tmp45171 : tmp44160;
  assign tmp45174 = s1 ? tmp44047 : tmp43953;
  assign tmp45177 = ~(l2 ? 1 : tmp43955);
  assign tmp45176 = s0 ? tmp44001 : tmp45177;
  assign tmp45178 = ~(l1 ? 1 : tmp43905);
  assign tmp45175 = ~(s1 ? tmp45176 : tmp45178);
  assign tmp45173 = ~(s2 ? tmp45174 : tmp45175);
  assign tmp45169 = s3 ? tmp45170 : tmp45173;
  assign tmp45181 = s1 ? tmp44062 : tmp44711;
  assign tmp45180 = s2 ? tmp45181 : tmp45146;
  assign tmp45184 = l1 ? tmp44544 : tmp43963;
  assign tmp45183 = ~(s0 ? tmp44001 : tmp45184);
  assign tmp45182 = s1 ? tmp44711 : tmp45183;
  assign tmp45179 = ~(s3 ? tmp45180 : tmp45182);
  assign tmp45168 = ~(s4 ? tmp45169 : tmp45179);
  assign tmp45140 = s5 ? tmp45141 : tmp45168;
  assign tmp45110 = s6 ? tmp45111 : tmp45140;
  assign tmp45109 = s7 ? tmp43890 : tmp45110;
  assign tmp45186 = s8 ? tmp45109 : tmp43890;
  assign tmp45192 = ~(l1 ? tmp44544 : tmp43963);
  assign tmp45191 = s1 ? tmp44711 : tmp45192;
  assign tmp45190 = ~(s3 ? tmp45180 : tmp45191);
  assign tmp45189 = ~(s4 ? tmp45169 : tmp45190);
  assign tmp45188 = s5 ? tmp45141 : tmp45189;
  assign tmp45187 = s6 ? tmp45111 : tmp45188;
  assign tmp45185 = s9 ? tmp45186 : tmp45187;
  assign tmp45108 = s10 ? tmp45109 : tmp45185;
  assign tmp45194 = s9 ? tmp45186 : tmp45110;
  assign tmp45193 = s10 ? tmp45109 : tmp45194;
  assign tmp45107 = s11 ? tmp45108 : tmp45193;
  assign tmp45010 = s12 ? tmp45011 : tmp45107;
  assign tmp44830 = s13 ? tmp44831 : tmp45010;
  assign tmp45206 = l1 ? tmp44011 : tmp43912;
  assign tmp45208 = ~(l1 ? tmp44011 : tmp43912);
  assign tmp45207 = ~(s0 ? tmp44491 : tmp45208);
  assign tmp45205 = s1 ? tmp45206 : tmp45207;
  assign tmp45213 = l2 ? tmp43906 : tmp43898;
  assign tmp45212 = l1 ? tmp44643 : tmp45213;
  assign tmp45211 = s0 ? tmp44491 : tmp45212;
  assign tmp45215 = l1 ? tmp44011 : tmp43921;
  assign tmp45216 = ~(l1 ? tmp44643 : tmp45213);
  assign tmp45214 = ~(s0 ? tmp45215 : tmp45216);
  assign tmp45210 = s1 ? tmp45211 : tmp45214;
  assign tmp45218 = s0 ? tmp45215 : tmp44417;
  assign tmp45219 = ~(s0 ? tmp45212 : tmp45208);
  assign tmp45217 = ~(s1 ? tmp45218 : tmp45219);
  assign tmp45209 = ~(s2 ? tmp45210 : tmp45217);
  assign tmp45204 = s3 ? tmp45205 : tmp45209;
  assign tmp45223 = s0 ? tmp45206 : tmp44508;
  assign tmp45224 = s0 ? tmp45206 : tmp45216;
  assign tmp45222 = s1 ? tmp45223 : tmp45224;
  assign tmp45226 = s0 ? tmp45206 : 1;
  assign tmp45225 = s1 ? tmp45226 : tmp44512;
  assign tmp45221 = s2 ? tmp45222 : tmp45225;
  assign tmp45228 = s1 ? tmp44491 : tmp43990;
  assign tmp45232 = ~(l2 ? tmp43906 : tmp43898);
  assign tmp45231 = ~(l1 ? tmp44011 : tmp45232);
  assign tmp45230 = s0 ? tmp45212 : tmp45231;
  assign tmp45234 = l1 ? tmp44005 : tmp44953;
  assign tmp45233 = ~(s0 ? tmp45234 : tmp45216);
  assign tmp45229 = s1 ? tmp45230 : tmp45233;
  assign tmp45227 = ~(s2 ? tmp45228 : tmp45229);
  assign tmp45220 = s3 ? tmp45221 : tmp45227;
  assign tmp45203 = s4 ? tmp45204 : tmp45220;
  assign tmp45240 = s0 ? tmp45206 : tmp43949;
  assign tmp45239 = s1 ? tmp45240 : tmp44671;
  assign tmp45242 = l1 ? tmp44674 : tmp43944;
  assign tmp45244 = l1 ? tmp44011 : tmp45232;
  assign tmp45243 = ~(s0 ? tmp45244 : 1);
  assign tmp45241 = ~(s1 ? tmp45242 : tmp45243);
  assign tmp45238 = s2 ? tmp45239 : tmp45241;
  assign tmp45247 = l1 ? tmp44680 : tmp43907;
  assign tmp45249 = l2 ? tmp43906 : tmp43955;
  assign tmp45248 = l1 ? tmp44682 : tmp45249;
  assign tmp45246 = s1 ? tmp45247 : tmp45248;
  assign tmp45251 = s0 ? tmp45234 : tmp44001;
  assign tmp45253 = l1 ? tmp44643 : tmp45249;
  assign tmp45255 = l2 ? tmp43897 : tmp43910;
  assign tmp45254 = ~(l1 ? tmp44011 : tmp45255);
  assign tmp45252 = ~(s0 ? tmp45253 : tmp45254);
  assign tmp45250 = ~(s1 ? tmp45251 : tmp45252);
  assign tmp45245 = ~(s2 ? tmp45246 : tmp45250);
  assign tmp45237 = s3 ? tmp45238 : tmp45245;
  assign tmp45260 = l1 ? tmp43955 : tmp43992;
  assign tmp45259 = s0 ? tmp45260 : tmp45208;
  assign tmp45258 = s1 ? tmp45259 : tmp44550;
  assign tmp45261 = ~(s1 ? tmp44010 : tmp44512);
  assign tmp45257 = s2 ? tmp45258 : tmp45261;
  assign tmp45265 = ~(l1 ? tmp44698 : tmp45249);
  assign tmp45264 = s0 ? tmp44017 : tmp45265;
  assign tmp45267 = l1 ? tmp44005 : tmp45255;
  assign tmp45266 = s0 ? tmp44010 : tmp45267;
  assign tmp45263 = s1 ? tmp45264 : tmp45266;
  assign tmp45269 = ~(l1 ? tmp43991 : tmp43992);
  assign tmp45268 = s1 ? tmp44001 : tmp45269;
  assign tmp45262 = ~(s2 ? tmp45263 : tmp45268);
  assign tmp45256 = ~(s3 ? tmp45257 : tmp45262);
  assign tmp45236 = s4 ? tmp45237 : tmp45256;
  assign tmp45274 = s0 ? tmp45248 : tmp44159;
  assign tmp45275 = ~(l2 ? tmp43963 : 1);
  assign tmp45273 = s1 ? tmp45274 : tmp45275;
  assign tmp45272 = s2 ? tmp45273 : tmp44782;
  assign tmp45279 = ~(l1 ? 1 : tmp44044);
  assign tmp45278 = s0 ? tmp44042 : tmp45279;
  assign tmp45277 = s1 ? tmp45278 : tmp44711;
  assign tmp45281 = l1 ? 1 : tmp43963;
  assign tmp45280 = ~(s1 ? tmp45281 : tmp44053);
  assign tmp45276 = s2 ? tmp45277 : tmp45280;
  assign tmp45271 = s3 ? tmp45272 : tmp45276;
  assign tmp45286 = l1 ? tmp44005 : tmp44044;
  assign tmp45285 = s0 ? tmp44059 : tmp45286;
  assign tmp45284 = s1 ? tmp45285 : tmp45234;
  assign tmp45287 = s1 ? tmp44017 : tmp44786;
  assign tmp45283 = s2 ? tmp45284 : tmp45287;
  assign tmp45291 = l2 ? tmp43955 : tmp43963;
  assign tmp45290 = l1 ? tmp44005 : tmp45291;
  assign tmp45292 = ~(l1 ? tmp44682 : tmp43992);
  assign tmp45289 = s1 ? tmp45290 : tmp45292;
  assign tmp45288 = s2 ? tmp45289 : tmp44059;
  assign tmp45282 = ~(s3 ? tmp45283 : tmp45288);
  assign tmp45270 = ~(s4 ? tmp45271 : tmp45282);
  assign tmp45235 = s5 ? tmp45236 : tmp45270;
  assign tmp45202 = s6 ? tmp45203 : tmp45235;
  assign tmp45201 = s7 ? tmp43890 : tmp45202;
  assign tmp45299 = ~(l1 ? tmp44005 : tmp43912);
  assign tmp45298 = ~(s0 ? tmp44583 : tmp45299);
  assign tmp45297 = s1 ? tmp44017 : tmp45298;
  assign tmp45303 = l1 ? tmp44732 : tmp45213;
  assign tmp45302 = s0 ? tmp44583 : tmp45303;
  assign tmp45305 = l1 ? tmp44005 : tmp43921;
  assign tmp45306 = ~(l1 ? tmp44732 : tmp45213);
  assign tmp45304 = ~(s0 ? tmp45305 : tmp45306);
  assign tmp45301 = s1 ? tmp45302 : tmp45304;
  assign tmp45308 = s0 ? tmp45305 : tmp44417;
  assign tmp45309 = ~(s0 ? tmp45303 : tmp45299);
  assign tmp45307 = ~(s1 ? tmp45308 : tmp45309);
  assign tmp45300 = ~(s2 ? tmp45301 : tmp45307);
  assign tmp45296 = s3 ? tmp45297 : tmp45300;
  assign tmp45313 = s0 ? tmp44017 : tmp44423;
  assign tmp45314 = s0 ? tmp44017 : tmp45306;
  assign tmp45312 = s1 ? tmp45313 : tmp45314;
  assign tmp45316 = s0 ? tmp44017 : 1;
  assign tmp45315 = s1 ? tmp45316 : tmp44589;
  assign tmp45311 = s2 ? tmp45312 : tmp45315;
  assign tmp45318 = s1 ? tmp44583 : tmp43990;
  assign tmp45321 = ~(l1 ? tmp44005 : tmp45232);
  assign tmp45320 = s0 ? tmp45303 : tmp45321;
  assign tmp45322 = ~(s0 ? tmp45234 : tmp45306);
  assign tmp45319 = s1 ? tmp45320 : tmp45322;
  assign tmp45317 = ~(s2 ? tmp45318 : tmp45319);
  assign tmp45310 = s3 ? tmp45311 : tmp45317;
  assign tmp45295 = s4 ? tmp45296 : tmp45310;
  assign tmp45328 = s0 ? tmp44017 : tmp43949;
  assign tmp45327 = s1 ? tmp45328 : tmp44756;
  assign tmp45330 = l1 ? tmp44759 : tmp43944;
  assign tmp45332 = l1 ? tmp44005 : tmp45232;
  assign tmp45331 = ~(s0 ? tmp45332 : 1);
  assign tmp45329 = ~(s1 ? tmp45330 : tmp45331);
  assign tmp45326 = s2 ? tmp45327 : tmp45329;
  assign tmp45335 = l1 ? tmp44765 : tmp43907;
  assign tmp45334 = s1 ? tmp45335 : tmp45248;
  assign tmp45338 = l1 ? tmp44732 : tmp45249;
  assign tmp45339 = ~(l1 ? tmp44005 : tmp45255);
  assign tmp45337 = ~(s0 ? tmp45338 : tmp45339);
  assign tmp45336 = ~(s1 ? tmp45251 : tmp45337);
  assign tmp45333 = ~(s2 ? tmp45334 : tmp45336);
  assign tmp45325 = s3 ? tmp45326 : tmp45333;
  assign tmp45343 = s0 ? tmp45260 : tmp45299;
  assign tmp45342 = s1 ? tmp45343 : tmp44609;
  assign tmp45344 = l1 ? tmp44009 : tmp43944;
  assign tmp45341 = s2 ? tmp45342 : tmp45344;
  assign tmp45348 = ~(l1 ? tmp43900 : tmp45249);
  assign tmp45347 = s0 ? tmp44017 : tmp45348;
  assign tmp45346 = s1 ? tmp45347 : tmp45267;
  assign tmp45345 = ~(s2 ? tmp45346 : tmp45268);
  assign tmp45340 = ~(s3 ? tmp45341 : tmp45345);
  assign tmp45324 = s4 ? tmp45325 : tmp45340;
  assign tmp45323 = s5 ? tmp45324 : tmp45270;
  assign tmp45294 = s6 ? tmp45295 : tmp45323;
  assign tmp45293 = s7 ? tmp43890 : tmp45294;
  assign tmp45200 = s8 ? tmp45201 : tmp45293;
  assign tmp45199 = s9 ? tmp45200 : tmp45293;
  assign tmp45350 = s8 ? tmp45293 : tmp43890;
  assign tmp45358 = s1 ? tmp45264 : tmp45267;
  assign tmp45357 = ~(s2 ? tmp45358 : tmp45268);
  assign tmp45356 = ~(s3 ? tmp45257 : tmp45357);
  assign tmp45355 = s4 ? tmp45237 : tmp45356;
  assign tmp45361 = s2 ? tmp45284 : tmp44017;
  assign tmp45360 = ~(s3 ? tmp45361 : tmp45289);
  assign tmp45359 = ~(s4 ? tmp45271 : tmp45360);
  assign tmp45354 = s5 ? tmp45355 : tmp45359;
  assign tmp45353 = s6 ? tmp45203 : tmp45354;
  assign tmp45363 = s5 ? tmp45324 : tmp45359;
  assign tmp45362 = s6 ? tmp45295 : tmp45363;
  assign tmp45352 = s7 ? tmp45353 : tmp45362;
  assign tmp45351 = s8 ? tmp45352 : tmp45362;
  assign tmp45349 = s9 ? tmp45350 : tmp45351;
  assign tmp45198 = s10 ? tmp45199 : tmp45349;
  assign tmp45367 = s7 ? tmp45202 : tmp45294;
  assign tmp45366 = s8 ? tmp45367 : tmp45294;
  assign tmp45365 = s9 ? tmp45350 : tmp45366;
  assign tmp45364 = s10 ? tmp45199 : tmp45365;
  assign tmp45197 = s11 ? tmp45198 : tmp45364;
  assign tmp45378 = l2 ? tmp43910 : tmp43955;
  assign tmp45377 = l1 ? tmp45378 : tmp43921;
  assign tmp45380 = ~(l1 ? tmp45378 : tmp43921);
  assign tmp45379 = ~(s0 ? tmp44583 : tmp45380);
  assign tmp45376 = s1 ? tmp45377 : tmp45379;
  assign tmp45385 = l2 ? tmp43955 : tmp44847;
  assign tmp45384 = l1 ? tmp45385 : tmp44498;
  assign tmp45383 = s0 ? tmp44491 : tmp45384;
  assign tmp45387 = ~(l1 ? tmp45385 : tmp44498);
  assign tmp45386 = ~(s0 ? tmp45377 : tmp45387);
  assign tmp45382 = s1 ? tmp45383 : tmp45386;
  assign tmp45389 = s0 ? tmp45377 : tmp44417;
  assign tmp45390 = ~(s0 ? tmp45384 : tmp45380);
  assign tmp45388 = ~(s1 ? tmp45389 : tmp45390);
  assign tmp45381 = ~(s2 ? tmp45382 : tmp45388);
  assign tmp45375 = s3 ? tmp45376 : tmp45381;
  assign tmp45394 = s0 ? tmp45215 : tmp44423;
  assign tmp45395 = s0 ? tmp45377 : tmp45387;
  assign tmp45393 = s1 ? tmp45394 : tmp45395;
  assign tmp45397 = s0 ? tmp45377 : 1;
  assign tmp45396 = s1 ? tmp45397 : tmp44589;
  assign tmp45392 = s2 ? tmp45393 : tmp45396;
  assign tmp45400 = l1 ? tmp45291 : tmp44045;
  assign tmp45399 = s1 ? tmp44583 : tmp45400;
  assign tmp45403 = ~(l1 ? tmp45378 : tmp44519);
  assign tmp45402 = s0 ? tmp45384 : tmp45403;
  assign tmp45405 = l1 ? tmp44031 : tmp44522;
  assign tmp45404 = ~(s0 ? tmp45405 : tmp45387);
  assign tmp45401 = s1 ? tmp45402 : tmp45404;
  assign tmp45398 = ~(s2 ? tmp45399 : tmp45401);
  assign tmp45391 = s3 ? tmp45392 : tmp45398;
  assign tmp45374 = s4 ? tmp45375 : tmp45391;
  assign tmp45411 = s0 ? tmp45377 : tmp43949;
  assign tmp45410 = s1 ? tmp45411 : tmp44671;
  assign tmp45414 = l2 ? 1 : tmp44847;
  assign tmp45413 = l1 ? tmp45414 : tmp44531;
  assign tmp45416 = l1 ? tmp45378 : tmp44519;
  assign tmp45415 = ~(s0 ? tmp45416 : 1);
  assign tmp45412 = ~(s1 ? tmp45413 : tmp45415);
  assign tmp45409 = s2 ? tmp45410 : tmp45412;
  assign tmp45420 = l2 ? tmp43955 : tmp43910;
  assign tmp45419 = l1 ? tmp45420 : tmp44538;
  assign tmp45418 = s1 ? tmp43904 : tmp45419;
  assign tmp45422 = s0 ? tmp45405 : tmp44988;
  assign tmp45424 = l1 ? tmp45385 : tmp44538;
  assign tmp45425 = ~(l1 ? tmp45378 : tmp44544);
  assign tmp45423 = ~(s0 ? tmp45424 : tmp45425);
  assign tmp45421 = ~(s1 ? tmp45422 : tmp45423);
  assign tmp45417 = ~(s2 ? tmp45418 : tmp45421);
  assign tmp45408 = s3 ? tmp45409 : tmp45417;
  assign tmp45430 = l1 ? tmp43954 : tmp44045;
  assign tmp45429 = s0 ? tmp45430 : tmp45380;
  assign tmp45428 = s1 ? tmp45429 : tmp44609;
  assign tmp45431 = l1 ? tmp44492 : tmp44531;
  assign tmp45427 = s2 ? tmp45428 : tmp45431;
  assign tmp45435 = ~(l1 ? tmp44135 : tmp44538);
  assign tmp45434 = s0 ? tmp45305 : tmp45435;
  assign tmp45436 = l1 ? tmp44031 : tmp44544;
  assign tmp45433 = s1 ? tmp45434 : tmp45436;
  assign tmp45438 = ~(l1 ? tmp45291 : tmp44045);
  assign tmp45437 = s1 ? tmp44001 : tmp45438;
  assign tmp45432 = ~(s2 ? tmp45433 : tmp45437);
  assign tmp45426 = ~(s3 ? tmp45427 : tmp45432);
  assign tmp45407 = s4 ? tmp45408 : tmp45426;
  assign tmp45443 = s0 ? tmp45419 : tmp44895;
  assign tmp45442 = s1 ? tmp45443 : tmp44030;
  assign tmp45445 = ~(l1 ? tmp43905 : 1);
  assign tmp45444 = ~(s1 ? tmp44033 : tmp45445);
  assign tmp45441 = s2 ? tmp45442 : tmp45444;
  assign tmp45448 = ~(l1 ? tmp44044 : tmp43992);
  assign tmp45447 = s1 ? 1 : tmp45448;
  assign tmp45450 = l1 ? tmp43992 : tmp44005;
  assign tmp45451 = l1 ? tmp44005 : tmp44162;
  assign tmp45449 = s1 ? tmp45450 : tmp45451;
  assign tmp45446 = ~(s2 ? tmp45447 : tmp45449);
  assign tmp45440 = s3 ? tmp45441 : tmp45446;
  assign tmp45455 = l1 ? tmp44031 : 1;
  assign tmp45454 = s1 ? tmp45455 : tmp45405;
  assign tmp45456 = l1 ? tmp44031 : tmp43921;
  assign tmp45453 = s2 ? tmp45454 : tmp45456;
  assign tmp45459 = l1 ? tmp44031 : tmp43954;
  assign tmp45458 = s0 ? tmp44034 : tmp45459;
  assign tmp45460 = ~(l1 ? tmp45420 : tmp44045);
  assign tmp45457 = s1 ? tmp45458 : tmp45460;
  assign tmp45452 = ~(s3 ? tmp45453 : tmp45457);
  assign tmp45439 = ~(s4 ? tmp45440 : tmp45452);
  assign tmp45406 = s5 ? tmp45407 : tmp45439;
  assign tmp45373 = s6 ? tmp45374 : tmp45406;
  assign tmp45372 = s7 ? tmp43890 : tmp45373;
  assign tmp45467 = ~(l1 ? tmp44031 : tmp43921);
  assign tmp45466 = ~(s0 ? tmp44583 : tmp45467);
  assign tmp45465 = s1 ? tmp45456 : tmp45466;
  assign tmp45472 = l2 ? tmp43900 : tmp44847;
  assign tmp45471 = l1 ? tmp45472 : tmp44498;
  assign tmp45470 = s0 ? tmp44583 : tmp45471;
  assign tmp45474 = ~(l1 ? tmp45472 : tmp44498);
  assign tmp45473 = ~(s0 ? tmp45456 : tmp45474);
  assign tmp45469 = s1 ? tmp45470 : tmp45473;
  assign tmp45476 = s0 ? tmp45456 : tmp44417;
  assign tmp45477 = ~(s0 ? tmp45471 : tmp45467);
  assign tmp45475 = ~(s1 ? tmp45476 : tmp45477);
  assign tmp45468 = ~(s2 ? tmp45469 : tmp45475);
  assign tmp45464 = s3 ? tmp45465 : tmp45468;
  assign tmp45481 = s0 ? tmp45305 : tmp44423;
  assign tmp45482 = s0 ? tmp45456 : tmp45474;
  assign tmp45480 = s1 ? tmp45481 : tmp45482;
  assign tmp45484 = s0 ? tmp45456 : 1;
  assign tmp45483 = s1 ? tmp45484 : tmp44589;
  assign tmp45479 = s2 ? tmp45480 : tmp45483;
  assign tmp45488 = ~(l1 ? tmp44031 : tmp44519);
  assign tmp45487 = s0 ? tmp45471 : tmp45488;
  assign tmp45489 = ~(s0 ? tmp45405 : tmp45474);
  assign tmp45486 = s1 ? tmp45487 : tmp45489;
  assign tmp45485 = ~(s2 ? tmp45399 : tmp45486);
  assign tmp45478 = s3 ? tmp45479 : tmp45485;
  assign tmp45463 = s4 ? tmp45464 : tmp45478;
  assign tmp45495 = s0 ? tmp45456 : tmp43949;
  assign tmp45494 = s1 ? tmp45495 : tmp44756;
  assign tmp45498 = l2 ? tmp43906 : tmp44847;
  assign tmp45497 = l1 ? tmp45498 : tmp44531;
  assign tmp45500 = l1 ? tmp44031 : tmp44519;
  assign tmp45499 = ~(s0 ? tmp45500 : 1);
  assign tmp45496 = ~(s1 ? tmp45497 : tmp45499);
  assign tmp45493 = s2 ? tmp45494 : tmp45496;
  assign tmp45503 = l1 ? tmp43906 : tmp43907;
  assign tmp45502 = s1 ? tmp45503 : tmp45419;
  assign tmp45506 = l1 ? tmp45472 : tmp44538;
  assign tmp45507 = ~(l1 ? tmp44031 : tmp44544);
  assign tmp45505 = ~(s0 ? tmp45506 : tmp45507);
  assign tmp45504 = ~(s1 ? tmp45422 : tmp45505);
  assign tmp45501 = ~(s2 ? tmp45502 : tmp45504);
  assign tmp45492 = s3 ? tmp45493 : tmp45501;
  assign tmp45511 = s0 ? tmp45430 : tmp45467;
  assign tmp45510 = s1 ? tmp45511 : tmp44609;
  assign tmp45512 = l1 ? tmp44009 : tmp44531;
  assign tmp45509 = s2 ? tmp45510 : tmp45512;
  assign tmp45517 = l2 ? tmp43900 : tmp43906;
  assign tmp45516 = ~(l1 ? tmp45517 : tmp44538);
  assign tmp45515 = s0 ? tmp45305 : tmp45516;
  assign tmp45514 = s1 ? tmp45515 : tmp45436;
  assign tmp45513 = ~(s2 ? tmp45514 : tmp45437);
  assign tmp45508 = ~(s3 ? tmp45509 : tmp45513);
  assign tmp45491 = s4 ? tmp45492 : tmp45508;
  assign tmp45520 = s2 ? tmp45442 : tmp44782;
  assign tmp45519 = s3 ? tmp45520 : tmp45446;
  assign tmp45522 = s1 ? tmp45459 : tmp45460;
  assign tmp45521 = ~(s3 ? tmp45453 : tmp45522);
  assign tmp45518 = ~(s4 ? tmp45519 : tmp45521);
  assign tmp45490 = s5 ? tmp45491 : tmp45518;
  assign tmp45462 = s6 ? tmp45463 : tmp45490;
  assign tmp45461 = s7 ? tmp43890 : tmp45462;
  assign tmp45371 = s8 ? tmp45372 : tmp45461;
  assign tmp45370 = s9 ? tmp45371 : tmp45461;
  assign tmp45524 = s8 ? tmp45461 : tmp43890;
  assign tmp45529 = ~(s4 ? tmp45440 : tmp45521);
  assign tmp45528 = s5 ? tmp45407 : tmp45529;
  assign tmp45527 = s6 ? tmp45374 : tmp45528;
  assign tmp45526 = s7 ? tmp45527 : tmp45462;
  assign tmp45525 = s8 ? tmp45526 : tmp45462;
  assign tmp45523 = s9 ? tmp45524 : tmp45525;
  assign tmp45369 = s10 ? tmp45370 : tmp45523;
  assign tmp45533 = s7 ? tmp45373 : tmp45462;
  assign tmp45532 = s8 ? tmp45533 : tmp45462;
  assign tmp45531 = s9 ? tmp45524 : tmp45532;
  assign tmp45530 = s10 ? tmp45370 : tmp45531;
  assign tmp45368 = s11 ? tmp45369 : tmp45530;
  assign tmp45196 = s12 ? tmp45197 : tmp45368;
  assign tmp45543 = ~(l2 ? tmp43896 : tmp43902);
  assign tmp45542 = l1 ? 1 : tmp45543;
  assign tmp45546 = ~(l2 ? tmp43896 : tmp43898);
  assign tmp45545 = ~(l1 ? tmp44044 : tmp45546);
  assign tmp45544 = ~(s0 ? tmp44404 : tmp45545);
  assign tmp45541 = s1 ? tmp45542 : tmp45544;
  assign tmp45552 = ~(l3 ? 1 : tmp43897);
  assign tmp45551 = l2 ? tmp43896 : tmp45552;
  assign tmp45550 = l1 ? tmp45551 : tmp43934;
  assign tmp45549 = s0 ? tmp44409 : tmp45550;
  assign tmp45554 = ~(l1 ? tmp45551 : tmp43934);
  assign tmp45553 = ~(s0 ? tmp44148 : tmp45554);
  assign tmp45548 = s1 ? tmp45549 : tmp45553;
  assign tmp45557 = ~(l1 ? tmp44044 : tmp45543);
  assign tmp45556 = ~(s0 ? tmp45550 : tmp45557);
  assign tmp45555 = ~(s1 ? tmp44416 : tmp45556);
  assign tmp45547 = ~(s2 ? tmp45548 : tmp45555);
  assign tmp45540 = s3 ? tmp45541 : tmp45547;
  assign tmp45562 = l1 ? 1 : tmp45546;
  assign tmp45561 = s0 ? tmp45562 : tmp44423;
  assign tmp45564 = l1 ? tmp44044 : tmp45543;
  assign tmp45563 = s0 ? tmp45564 : tmp45554;
  assign tmp45560 = s1 ? tmp45561 : tmp45563;
  assign tmp45566 = s0 ? tmp45542 : 1;
  assign tmp45565 = s1 ? tmp45566 : tmp44427;
  assign tmp45559 = s2 ? tmp45560 : tmp45565;
  assign tmp45569 = l1 ? tmp43955 : tmp44005;
  assign tmp45568 = s1 ? tmp44404 : tmp45569;
  assign tmp45573 = ~(l2 ? tmp43910 : tmp43902);
  assign tmp45572 = ~(l1 ? tmp44044 : tmp45573);
  assign tmp45571 = s0 ? tmp45550 : tmp45572;
  assign tmp45575 = l1 ? tmp44044 : tmp43991;
  assign tmp45574 = ~(s0 ? tmp45575 : tmp45554);
  assign tmp45570 = s1 ? tmp45571 : tmp45574;
  assign tmp45567 = ~(s2 ? tmp45568 : tmp45570);
  assign tmp45558 = s3 ? tmp45559 : tmp45567;
  assign tmp45539 = s4 ? tmp45540 : tmp45558;
  assign tmp45582 = l1 ? tmp44044 : tmp45546;
  assign tmp45581 = s0 ? tmp45582 : tmp43949;
  assign tmp45580 = s1 ? tmp45581 : tmp44439;
  assign tmp45585 = l2 ? tmp43910 : tmp45552;
  assign tmp45584 = l1 ? tmp45585 : tmp44011;
  assign tmp45587 = l1 ? tmp44044 : tmp45573;
  assign tmp45586 = ~(s0 ? tmp45587 : 1);
  assign tmp45583 = ~(s1 ? tmp45584 : tmp45586);
  assign tmp45579 = s2 ? tmp45580 : tmp45583;
  assign tmp45590 = l1 ? tmp44213 : tmp44011;
  assign tmp45589 = s1 ? tmp44128 : tmp45590;
  assign tmp45593 = l1 ? tmp44044 : tmp43955;
  assign tmp45592 = s0 ? tmp45575 : tmp45593;
  assign tmp45595 = l1 ? tmp45551 : tmp44011;
  assign tmp45596 = ~(l1 ? tmp44044 : tmp44682);
  assign tmp45594 = ~(s0 ? tmp45595 : tmp45596);
  assign tmp45591 = ~(s1 ? tmp45592 : tmp45594);
  assign tmp45588 = ~(s2 ? tmp45589 : tmp45591);
  assign tmp45578 = s3 ? tmp45579 : tmp45588;
  assign tmp45600 = s0 ? tmp45569 : tmp45557;
  assign tmp45599 = s1 ? tmp45600 : tmp44451;
  assign tmp45601 = l1 ? tmp44410 : tmp44011;
  assign tmp45598 = s2 ? tmp45599 : tmp45601;
  assign tmp45605 = ~(l1 ? tmp44150 : tmp44011);
  assign tmp45604 = s0 ? tmp45562 : tmp45605;
  assign tmp45606 = l1 ? tmp44044 : tmp44682;
  assign tmp45603 = s1 ? tmp45604 : tmp45606;
  assign tmp45608 = l1 ? 1 : tmp43955;
  assign tmp45609 = ~(l1 ? tmp43955 : tmp44005);
  assign tmp45607 = s1 ? tmp45608 : tmp45609;
  assign tmp45602 = ~(s2 ? tmp45603 : tmp45607);
  assign tmp45597 = ~(s3 ? tmp45598 : tmp45602);
  assign tmp45577 = s4 ? tmp45578 : tmp45597;
  assign tmp45614 = s0 ? tmp45590 : tmp44159;
  assign tmp45613 = s1 ? tmp45614 : 0;
  assign tmp45612 = s2 ? tmp45613 : tmp44160;
  assign tmp45617 = l1 ? tmp44044 : tmp44045;
  assign tmp45618 = s0 ? tmp44047 : tmp44903;
  assign tmp45616 = s1 ? tmp45617 : tmp45618;
  assign tmp45621 = l2 ? 1 : tmp43910;
  assign tmp45620 = l1 ? 1 : tmp45621;
  assign tmp45619 = s1 ? tmp45087 : tmp45620;
  assign tmp45615 = ~(s2 ? tmp45616 : tmp45619);
  assign tmp45611 = s3 ? tmp45612 : tmp45615;
  assign tmp45624 = s1 ? tmp44044 : tmp45575;
  assign tmp45623 = s2 ? tmp45624 : tmp45582;
  assign tmp45627 = ~(l1 ? tmp44213 : tmp44005);
  assign tmp45626 = s1 ? tmp45575 : tmp45627;
  assign tmp45625 = s2 ? tmp45626 : tmp44047;
  assign tmp45622 = ~(s3 ? tmp45623 : tmp45625);
  assign tmp45610 = ~(s4 ? tmp45611 : tmp45622);
  assign tmp45576 = s5 ? tmp45577 : tmp45610;
  assign tmp45538 = s6 ? tmp45539 : tmp45576;
  assign tmp45537 = s7 ? tmp43890 : tmp45538;
  assign tmp45629 = s8 ? tmp45537 : tmp43890;
  assign tmp45633 = ~(s3 ? tmp45623 : tmp45626);
  assign tmp45632 = ~(s4 ? tmp45611 : tmp45633);
  assign tmp45631 = s5 ? tmp45577 : tmp45632;
  assign tmp45630 = s6 ? tmp45539 : tmp45631;
  assign tmp45628 = s9 ? tmp45629 : tmp45630;
  assign tmp45536 = s10 ? tmp45537 : tmp45628;
  assign tmp45635 = s9 ? tmp45629 : tmp45538;
  assign tmp45634 = s10 ? tmp45537 : tmp45635;
  assign tmp45535 = s11 ? tmp45536 : tmp45634;
  assign tmp45645 = l1 ? tmp45378 : tmp45546;
  assign tmp45647 = ~(l1 ? tmp44131 : tmp45546);
  assign tmp45646 = ~(s0 ? tmp44637 : tmp45647);
  assign tmp45644 = s1 ? tmp45645 : tmp45646;
  assign tmp45652 = l2 ? tmp43955 : tmp43901;
  assign tmp45651 = l1 ? tmp45652 : tmp43920;
  assign tmp45650 = s0 ? tmp44491 : tmp45651;
  assign tmp45654 = l1 ? tmp45378 : tmp44038;
  assign tmp45655 = ~(l1 ? tmp45652 : tmp43920);
  assign tmp45653 = ~(s0 ? tmp45654 : tmp45655);
  assign tmp45649 = s1 ? tmp45650 : tmp45653;
  assign tmp45657 = s0 ? tmp45654 : tmp44417;
  assign tmp45658 = ~(s0 ? tmp45651 : tmp45647);
  assign tmp45656 = ~(s1 ? tmp45657 : tmp45658);
  assign tmp45648 = ~(s2 ? tmp45649 : tmp45656);
  assign tmp45643 = s3 ? tmp45644 : tmp45648;
  assign tmp45663 = l1 ? tmp44011 : tmp45546;
  assign tmp45662 = s0 ? tmp45663 : tmp44423;
  assign tmp45665 = l1 ? tmp44131 : tmp45546;
  assign tmp45664 = s0 ? tmp45665 : tmp45655;
  assign tmp45661 = s1 ? tmp45662 : tmp45664;
  assign tmp45667 = s0 ? tmp45645 : 1;
  assign tmp45666 = s1 ? tmp45667 : tmp44427;
  assign tmp45660 = s2 ? tmp45661 : tmp45666;
  assign tmp45670 = l1 ? tmp43954 : tmp44031;
  assign tmp45669 = s1 ? tmp44404 : tmp45670;
  assign tmp45674 = ~(l2 ? tmp43910 : tmp43898);
  assign tmp45673 = ~(l1 ? tmp44131 : tmp45674);
  assign tmp45672 = s0 ? tmp45651 : tmp45673;
  assign tmp45676 = l1 ? tmp43962 : tmp45291;
  assign tmp45675 = ~(s0 ? tmp45676 : tmp45655);
  assign tmp45671 = s1 ? tmp45672 : tmp45675;
  assign tmp45668 = ~(s2 ? tmp45669 : tmp45671);
  assign tmp45659 = s3 ? tmp45660 : tmp45668;
  assign tmp45642 = s4 ? tmp45643 : tmp45659;
  assign tmp45682 = s0 ? tmp45665 : tmp43949;
  assign tmp45681 = s1 ? tmp45682 : tmp44671;
  assign tmp45684 = l1 ? tmp44492 : tmp44011;
  assign tmp45686 = l1 ? tmp44131 : tmp45674;
  assign tmp45685 = ~(s0 ? tmp45686 : 1);
  assign tmp45683 = ~(s1 ? tmp45684 : tmp45685);
  assign tmp45680 = s2 ? tmp45681 : tmp45683;
  assign tmp45689 = l1 ? tmp44135 : tmp45378;
  assign tmp45688 = s1 ? tmp44081 : tmp45689;
  assign tmp45692 = l1 ? tmp44045 : tmp43954;
  assign tmp45691 = s0 ? tmp45676 : tmp45692;
  assign tmp45694 = l1 ? tmp45652 : tmp45378;
  assign tmp45695 = ~(l1 ? tmp44131 : tmp45420);
  assign tmp45693 = ~(s0 ? tmp45694 : tmp45695);
  assign tmp45690 = ~(s1 ? tmp45691 : tmp45693);
  assign tmp45687 = ~(s2 ? tmp45688 : tmp45690);
  assign tmp45679 = s3 ? tmp45680 : tmp45687;
  assign tmp45699 = s0 ? tmp45670 : tmp45647;
  assign tmp45698 = s1 ? tmp45699 : tmp44451;
  assign tmp45697 = s2 ? tmp45698 : tmp45684;
  assign tmp45703 = l1 ? tmp44005 : tmp45546;
  assign tmp45704 = ~(l1 ? tmp44135 : tmp45378);
  assign tmp45702 = s0 ? tmp45703 : tmp45704;
  assign tmp45705 = l1 ? tmp43962 : tmp45420;
  assign tmp45701 = s1 ? tmp45702 : tmp45705;
  assign tmp45707 = ~(l1 ? tmp43954 : tmp44031);
  assign tmp45706 = s1 ? tmp44001 : tmp45707;
  assign tmp45700 = ~(s2 ? tmp45701 : tmp45706);
  assign tmp45696 = ~(s3 ? tmp45697 : tmp45700);
  assign tmp45678 = s4 ? tmp45679 : tmp45696;
  assign tmp45712 = s0 ? tmp45689 : tmp44895;
  assign tmp45713 = ~(l1 ? tmp44031 : 1);
  assign tmp45711 = s1 ? tmp45712 : tmp45713;
  assign tmp45710 = s2 ? tmp45711 : tmp44782;
  assign tmp45716 = ~(l1 ? 1 : tmp43992);
  assign tmp45715 = s1 ? tmp44044 : tmp45716;
  assign tmp45718 = l1 ? tmp44005 : tmp45621;
  assign tmp45717 = s1 ? tmp45094 : tmp45718;
  assign tmp45714 = ~(s2 ? tmp45715 : tmp45717);
  assign tmp45709 = s3 ? tmp45710 : tmp45714;
  assign tmp45722 = s0 ? tmp44062 : tmp45676;
  assign tmp45721 = s1 ? tmp44060 : tmp45722;
  assign tmp45723 = l1 ? tmp43962 : tmp45546;
  assign tmp45720 = s2 ? tmp45721 : tmp45723;
  assign tmp45726 = ~(l1 ? tmp44135 : tmp44031);
  assign tmp45725 = s1 ? tmp45676 : tmp45726;
  assign tmp45724 = s2 ? tmp45725 : tmp44062;
  assign tmp45719 = ~(s3 ? tmp45720 : tmp45724);
  assign tmp45708 = ~(s4 ? tmp45709 : tmp45719);
  assign tmp45677 = s5 ? tmp45678 : tmp45708;
  assign tmp45641 = s6 ? tmp45642 : tmp45677;
  assign tmp45640 = s7 ? tmp43890 : tmp45641;
  assign tmp45732 = l1 ? tmp44031 : tmp45546;
  assign tmp45734 = ~(l1 ? tmp43962 : tmp45546);
  assign tmp45733 = ~(s0 ? tmp44404 : tmp45734);
  assign tmp45731 = s1 ? tmp45732 : tmp45733;
  assign tmp45739 = l2 ? tmp43900 : tmp43901;
  assign tmp45738 = l1 ? tmp45739 : tmp43920;
  assign tmp45737 = s0 ? tmp44583 : tmp45738;
  assign tmp45741 = l1 ? tmp44031 : tmp44038;
  assign tmp45742 = ~(l1 ? tmp45739 : tmp43920);
  assign tmp45740 = ~(s0 ? tmp45741 : tmp45742);
  assign tmp45736 = s1 ? tmp45737 : tmp45740;
  assign tmp45744 = s0 ? tmp45741 : tmp44417;
  assign tmp45745 = ~(s0 ? tmp45738 : tmp45734);
  assign tmp45743 = ~(s1 ? tmp45744 : tmp45745);
  assign tmp45735 = ~(s2 ? tmp45736 : tmp45743);
  assign tmp45730 = s3 ? tmp45731 : tmp45735;
  assign tmp45749 = s0 ? tmp45703 : tmp44423;
  assign tmp45750 = s0 ? tmp45723 : tmp45742;
  assign tmp45748 = s1 ? tmp45749 : tmp45750;
  assign tmp45752 = s0 ? tmp45732 : 1;
  assign tmp45751 = s1 ? tmp45752 : tmp44427;
  assign tmp45747 = s2 ? tmp45748 : tmp45751;
  assign tmp45756 = ~(l1 ? tmp43962 : tmp45674);
  assign tmp45755 = s0 ? tmp45738 : tmp45756;
  assign tmp45757 = ~(s0 ? tmp45676 : tmp45742);
  assign tmp45754 = s1 ? tmp45755 : tmp45757;
  assign tmp45753 = ~(s2 ? tmp45669 : tmp45754);
  assign tmp45746 = s3 ? tmp45747 : tmp45753;
  assign tmp45729 = s4 ? tmp45730 : tmp45746;
  assign tmp45763 = s0 ? tmp45723 : tmp43949;
  assign tmp45762 = s1 ? tmp45763 : tmp44756;
  assign tmp45765 = l1 ? tmp44009 : tmp44011;
  assign tmp45767 = l1 ? tmp43962 : tmp45674;
  assign tmp45766 = ~(s0 ? tmp45767 : 1);
  assign tmp45764 = ~(s1 ? tmp45765 : tmp45766);
  assign tmp45761 = s2 ? tmp45762 : tmp45764;
  assign tmp45769 = s1 ? tmp44221 : tmp45689;
  assign tmp45772 = l1 ? tmp45739 : tmp45378;
  assign tmp45773 = ~(l1 ? tmp43962 : tmp45420);
  assign tmp45771 = ~(s0 ? tmp45772 : tmp45773);
  assign tmp45770 = ~(s1 ? tmp45691 : tmp45771);
  assign tmp45768 = ~(s2 ? tmp45769 : tmp45770);
  assign tmp45760 = s3 ? tmp45761 : tmp45768;
  assign tmp45777 = s0 ? tmp45670 : tmp45734;
  assign tmp45776 = s1 ? tmp45777 : tmp44451;
  assign tmp45775 = s2 ? tmp45776 : tmp45765;
  assign tmp45781 = ~(l1 ? tmp45517 : tmp45378);
  assign tmp45780 = s0 ? tmp45703 : tmp45781;
  assign tmp45779 = s1 ? tmp45780 : tmp45705;
  assign tmp45778 = ~(s2 ? tmp45779 : tmp45706);
  assign tmp45774 = ~(s3 ? tmp45775 : tmp45778);
  assign tmp45759 = s4 ? tmp45760 : tmp45774;
  assign tmp45758 = s5 ? tmp45759 : tmp45708;
  assign tmp45728 = s6 ? tmp45729 : tmp45758;
  assign tmp45727 = s7 ? tmp43890 : tmp45728;
  assign tmp45639 = s8 ? tmp45640 : tmp45727;
  assign tmp45638 = s9 ? tmp45639 : tmp45727;
  assign tmp45783 = s8 ? tmp45727 : tmp43890;
  assign tmp45789 = ~(s3 ? tmp45720 : tmp45725);
  assign tmp45788 = ~(s4 ? tmp45709 : tmp45789);
  assign tmp45787 = s5 ? tmp45678 : tmp45788;
  assign tmp45786 = s6 ? tmp45642 : tmp45787;
  assign tmp45791 = s5 ? tmp45759 : tmp45788;
  assign tmp45790 = s6 ? tmp45729 : tmp45791;
  assign tmp45785 = s7 ? tmp45786 : tmp45790;
  assign tmp45784 = s8 ? tmp45785 : tmp45790;
  assign tmp45782 = s9 ? tmp45783 : tmp45784;
  assign tmp45637 = s10 ? tmp45638 : tmp45782;
  assign tmp45795 = s7 ? tmp45641 : tmp45728;
  assign tmp45794 = s8 ? tmp45795 : tmp45728;
  assign tmp45793 = s9 ? tmp45783 : tmp45794;
  assign tmp45792 = s10 ? tmp45638 : tmp45793;
  assign tmp45636 = s11 ? tmp45637 : tmp45792;
  assign tmp45534 = s12 ? tmp45535 : tmp45636;
  assign tmp45195 = s13 ? tmp45196 : tmp45534;
  assign tmp44829 = s14 ? tmp44830 : tmp45195;
  assign tmp43882 = s15 ? tmp43883 : tmp44829;
  assign tmp45810 = ~(s0 ? tmp44208 : tmp44013);
  assign tmp45809 = ~(s1 ? tmp44008 : tmp45810);
  assign tmp45808 = s2 ? tmp44138 : tmp45809;
  assign tmp45807 = ~(s3 ? tmp45808 : tmp44209);
  assign tmp45806 = s4 ? tmp44195 : tmp45807;
  assign tmp45805 = s5 ? tmp45806 : tmp44154;
  assign tmp45804 = s6 ? tmp44176 : tmp45805;
  assign tmp45803 = s7 ? tmp43890 : tmp45804;
  assign tmp45802 = s8 ? tmp43889 : tmp45803;
  assign tmp45801 = s9 ? tmp45802 : tmp45803;
  assign tmp45812 = s8 ? tmp45803 : tmp43890;
  assign tmp45821 = ~(l1 ? tmp44162 : tmp44123);
  assign tmp45820 = ~(s1 ? tmp44008 : tmp45821);
  assign tmp45819 = s2 ? tmp44138 : tmp45820;
  assign tmp45818 = ~(s3 ? tmp45819 : tmp44209);
  assign tmp45817 = s4 ? tmp44195 : tmp45818;
  assign tmp45816 = s5 ? tmp45817 : tmp44154;
  assign tmp45815 = s6 ? tmp44176 : tmp45816;
  assign tmp45814 = s7 ? tmp44269 : tmp45815;
  assign tmp45813 = s8 ? tmp45814 : tmp45815;
  assign tmp45811 = s9 ? tmp45812 : tmp45813;
  assign tmp45800 = s10 ? tmp45801 : tmp45811;
  assign tmp45825 = s7 ? tmp44075 : tmp45804;
  assign tmp45824 = s8 ? tmp45825 : tmp45804;
  assign tmp45823 = s9 ? tmp45812 : tmp45824;
  assign tmp45822 = s10 ? tmp45801 : tmp45823;
  assign tmp45799 = s11 ? tmp45800 : tmp45822;
  assign tmp45838 = l1 ? tmp43905 : tmp44011;
  assign tmp45837 = ~(s0 ? tmp45838 : tmp43945);
  assign tmp45836 = s1 ? tmp44192 : tmp45837;
  assign tmp45835 = s2 ? tmp44189 : tmp45836;
  assign tmp45840 = s1 ? tmp44081 : tmp44301;
  assign tmp45839 = ~(s2 ? tmp45840 : tmp44108);
  assign tmp45834 = s3 ? tmp45835 : tmp45839;
  assign tmp45833 = s4 ? tmp44177 : tmp45834;
  assign tmp45832 = s6 ? tmp45833 : tmp44193;
  assign tmp45831 = s7 ? tmp43890 : tmp45832;
  assign tmp45830 = s8 ? tmp44373 : tmp45831;
  assign tmp45829 = s9 ? tmp45830 : tmp45831;
  assign tmp45842 = s8 ? tmp45831 : tmp43890;
  assign tmp45847 = s3 ? tmp45835 : tmp44105;
  assign tmp45846 = s4 ? tmp44177 : tmp45847;
  assign tmp45845 = s6 ? tmp45846 : tmp44193;
  assign tmp45844 = s7 ? tmp44385 : tmp45845;
  assign tmp45843 = s8 ? tmp45844 : tmp45845;
  assign tmp45841 = s9 ? tmp45842 : tmp45843;
  assign tmp45828 = s10 ? tmp45829 : tmp45841;
  assign tmp45851 = s7 ? tmp44374 : tmp45832;
  assign tmp45850 = s8 ? tmp45851 : tmp45832;
  assign tmp45849 = s9 ? tmp45842 : tmp45850;
  assign tmp45848 = s10 ? tmp45829 : tmp45849;
  assign tmp45827 = s11 ? tmp45828 : tmp45848;
  assign tmp45826 = s12 ? tmp44282 : tmp45827;
  assign tmp45798 = s13 ? tmp45799 : tmp45826;
  assign tmp45861 = l1 ? tmp43944 : tmp44038;
  assign tmp45863 = ~(l1 ? tmp43944 : tmp44038);
  assign tmp45862 = ~(s0 ? tmp44637 : tmp45863);
  assign tmp45860 = s1 ? tmp45861 : tmp45862;
  assign tmp45868 = l2 ? tmp43963 : tmp43901;
  assign tmp45867 = l1 ? tmp45868 : tmp43907;
  assign tmp45870 = l2 ? tmp43897 : 0;
  assign tmp45869 = l1 ? tmp45870 : tmp43909;
  assign tmp45866 = s0 ? tmp45867 : tmp45869;
  assign tmp45872 = ~(l1 ? tmp45870 : tmp43909);
  assign tmp45871 = ~(s0 ? tmp45861 : tmp45872);
  assign tmp45865 = s1 ? tmp45866 : tmp45871;
  assign tmp45874 = s0 ? tmp45861 : tmp44648;
  assign tmp45875 = ~(s0 ? tmp45869 : tmp45863);
  assign tmp45873 = ~(s1 ? tmp45874 : tmp45875);
  assign tmp45864 = ~(s2 ? tmp45865 : tmp45873);
  assign tmp45859 = s3 ? tmp45860 : tmp45864;
  assign tmp45879 = s0 ? tmp45861 : tmp44508;
  assign tmp45880 = s0 ? tmp45861 : tmp45872;
  assign tmp45878 = s1 ? tmp45879 : tmp45880;
  assign tmp45882 = s0 ? tmp45861 : tmp43979;
  assign tmp45881 = s1 ? tmp45882 : tmp44657;
  assign tmp45877 = s2 ? tmp45878 : tmp45881;
  assign tmp45885 = s0 ? tmp45869 : tmp44110;
  assign tmp45886 = ~(s0 ? tmp44001 : tmp45872);
  assign tmp45884 = s1 ? tmp45885 : tmp45886;
  assign tmp45883 = ~(s2 ? tmp44659 : tmp45884);
  assign tmp45876 = s3 ? tmp45877 : tmp45883;
  assign tmp45858 = s4 ? tmp45859 : tmp45876;
  assign tmp45892 = s0 ? tmp45861 : tmp43949;
  assign tmp45893 = ~(l1 ? tmp45868 : tmp43907);
  assign tmp45891 = s1 ? tmp45892 : tmp45893;
  assign tmp45896 = l2 ? tmp43963 : 0;
  assign tmp45895 = l1 ? tmp45896 : tmp44123;
  assign tmp45894 = ~(s1 ? tmp45895 : tmp44124);
  assign tmp45890 = s2 ? tmp45891 : tmp45894;
  assign tmp45900 = ~(l1 ? tmp44205 : tmp43934);
  assign tmp45899 = s0 ? tmp43983 : tmp45900;
  assign tmp45898 = s1 ? tmp45899 : tmp44316;
  assign tmp45903 = l1 ? tmp45870 : tmp44131;
  assign tmp45902 = ~(s0 ? tmp45903 : tmp44134);
  assign tmp45901 = s1 ? tmp44001 : tmp45902;
  assign tmp45897 = s2 ? tmp45898 : tmp45901;
  assign tmp45889 = s3 ? tmp45890 : tmp45897;
  assign tmp45907 = s0 ? tmp44140 : tmp45863;
  assign tmp45906 = s1 ? tmp45907 : tmp44692;
  assign tmp45908 = l1 ? tmp45868 : tmp44123;
  assign tmp45905 = s2 ? tmp45906 : tmp45908;
  assign tmp45904 = ~(s3 ? tmp45905 : tmp44209);
  assign tmp45888 = s4 ? tmp45889 : tmp45904;
  assign tmp45887 = s5 ? tmp45888 : tmp44154;
  assign tmp45857 = s6 ? tmp45858 : tmp45887;
  assign tmp45856 = s7 ? tmp43890 : tmp45857;
  assign tmp45910 = s8 ? tmp45856 : tmp43890;
  assign tmp45918 = s1 ? tmp45899 : tmp44317;
  assign tmp45917 = s2 ? tmp45918 : tmp45901;
  assign tmp45916 = s3 ? tmp45890 : tmp45917;
  assign tmp45915 = s4 ? tmp45916 : tmp45904;
  assign tmp45914 = s5 ? tmp45915 : tmp44154;
  assign tmp45913 = s6 ? tmp45858 : tmp45914;
  assign tmp45912 = s7 ? tmp44471 : tmp45913;
  assign tmp45911 = s8 ? tmp45912 : tmp45913;
  assign tmp45909 = s9 ? tmp45910 : tmp45911;
  assign tmp45855 = s10 ? tmp45856 : tmp45909;
  assign tmp45922 = s7 ? tmp44399 : tmp45857;
  assign tmp45921 = s8 ? tmp45922 : tmp45857;
  assign tmp45920 = s9 ? tmp45910 : tmp45921;
  assign tmp45919 = s10 ? tmp45856 : tmp45920;
  assign tmp45854 = s11 ? tmp45855 : tmp45919;
  assign tmp45930 = l1 ? tmp43944 : tmp43921;
  assign tmp45932 = ~(l1 ? tmp43944 : tmp43921);
  assign tmp45931 = ~(s0 ? tmp44491 : tmp45932);
  assign tmp45929 = s1 ? tmp45930 : tmp45931;
  assign tmp45936 = l1 ? tmp45870 : tmp44498;
  assign tmp45935 = s0 ? tmp45867 : tmp45936;
  assign tmp45938 = ~(l1 ? tmp45870 : tmp44498);
  assign tmp45937 = ~(s0 ? tmp45930 : tmp45938);
  assign tmp45934 = s1 ? tmp45935 : tmp45937;
  assign tmp45940 = s0 ? tmp45930 : tmp44648;
  assign tmp45941 = ~(s0 ? tmp45936 : tmp45932);
  assign tmp45939 = ~(s1 ? tmp45940 : tmp45941);
  assign tmp45933 = ~(s2 ? tmp45934 : tmp45939);
  assign tmp45928 = s3 ? tmp45929 : tmp45933;
  assign tmp45945 = s0 ? tmp45930 : tmp44508;
  assign tmp45946 = s0 ? tmp45930 : tmp45938;
  assign tmp45944 = s1 ? tmp45945 : tmp45946;
  assign tmp45948 = s0 ? tmp45930 : tmp43979;
  assign tmp45947 = s1 ? tmp45948 : tmp44512;
  assign tmp45943 = s2 ? tmp45944 : tmp45947;
  assign tmp45951 = s0 ? tmp45936 : tmp44518;
  assign tmp45952 = ~(s0 ? tmp44521 : tmp45938);
  assign tmp45950 = s1 ? tmp45951 : tmp45952;
  assign tmp45949 = ~(s2 ? tmp44514 : tmp45950);
  assign tmp45942 = s3 ? tmp45943 : tmp45949;
  assign tmp45927 = s4 ? tmp45928 : tmp45942;
  assign tmp45958 = s0 ? tmp45930 : tmp43949;
  assign tmp45957 = s1 ? tmp45958 : tmp45893;
  assign tmp45960 = l1 ? tmp45896 : tmp44531;
  assign tmp45961 = ~(s0 ? tmp44533 : tmp43979);
  assign tmp45959 = ~(s1 ? tmp45960 : tmp45961);
  assign tmp45956 = s2 ? tmp45957 : tmp45959;
  assign tmp45964 = l1 ? tmp44205 : tmp43907;
  assign tmp45963 = s1 ? tmp45964 : tmp44537;
  assign tmp45967 = l1 ? tmp45870 : tmp44538;
  assign tmp45966 = ~(s0 ? tmp45967 : tmp44543);
  assign tmp45965 = ~(s1 ? tmp44540 : tmp45966);
  assign tmp45962 = ~(s2 ? tmp45963 : tmp45965);
  assign tmp45955 = s3 ? tmp45956 : tmp45962;
  assign tmp45971 = s0 ? tmp44549 : tmp45932;
  assign tmp45970 = s1 ? tmp45971 : tmp44550;
  assign tmp45973 = ~(l1 ? tmp45868 : tmp44531);
  assign tmp45972 = ~(s1 ? tmp44010 : tmp45973);
  assign tmp45969 = s2 ? tmp45970 : tmp45972;
  assign tmp45977 = ~(l1 ? tmp44213 : tmp44538);
  assign tmp45976 = s0 ? tmp44489 : tmp45977;
  assign tmp45975 = s1 ? tmp45976 : tmp44558;
  assign tmp45974 = ~(s2 ? tmp45975 : tmp44560);
  assign tmp45968 = ~(s3 ? tmp45969 : tmp45974);
  assign tmp45954 = s4 ? tmp45955 : tmp45968;
  assign tmp45953 = s5 ? tmp45954 : tmp44562;
  assign tmp45926 = s6 ? tmp45927 : tmp45953;
  assign tmp45925 = s7 ? tmp43890 : tmp45926;
  assign tmp45979 = s8 ? tmp45925 : tmp43890;
  assign tmp45985 = s1 ? tmp45976 : tmp44559;
  assign tmp45984 = ~(s2 ? tmp45985 : tmp44560);
  assign tmp45983 = ~(s3 ? tmp45969 : tmp45984);
  assign tmp45982 = s4 ? tmp45955 : tmp45983;
  assign tmp45981 = s5 ? tmp45982 : tmp44562;
  assign tmp45980 = s6 ? tmp45927 : tmp45981;
  assign tmp45978 = s9 ? tmp45979 : tmp45980;
  assign tmp45924 = s10 ? tmp45925 : tmp45978;
  assign tmp45987 = s9 ? tmp45979 : tmp45926;
  assign tmp45986 = s10 ? tmp45925 : tmp45987;
  assign tmp45923 = s11 ? tmp45924 : tmp45986;
  assign tmp45853 = s12 ? tmp45854 : tmp45923;
  assign tmp45999 = s1 ? 1 : tmp44042;
  assign tmp45998 = ~(s2 ? tmp44165 : tmp45999);
  assign tmp45997 = s3 ? tmp44781 : tmp45998;
  assign tmp45996 = ~(s4 ? tmp45997 : tmp44794);
  assign tmp45995 = s5 ? tmp44666 : tmp45996;
  assign tmp45994 = s6 ? tmp44632 : tmp45995;
  assign tmp45993 = s7 ? tmp43890 : tmp45994;
  assign tmp46002 = s5 ? tmp44751 : tmp45996;
  assign tmp46001 = s6 ? tmp44723 : tmp46002;
  assign tmp46000 = s7 ? tmp43890 : tmp46001;
  assign tmp45992 = s8 ? tmp45993 : tmp46000;
  assign tmp46006 = s5 ? tmp44751 : tmp44700;
  assign tmp46005 = s6 ? tmp44723 : tmp46006;
  assign tmp46004 = s7 ? tmp43890 : tmp46005;
  assign tmp46003 = s8 ? tmp46000 : tmp46004;
  assign tmp45991 = s9 ? tmp45992 : tmp46003;
  assign tmp46008 = s8 ? tmp46000 : tmp43890;
  assign tmp46012 = s5 ? tmp44751 : tmp44793;
  assign tmp46011 = s6 ? tmp44723 : tmp46012;
  assign tmp46010 = s7 ? tmp45994 : tmp46011;
  assign tmp46009 = s8 ? tmp46010 : tmp46001;
  assign tmp46007 = s9 ? tmp46008 : tmp46009;
  assign tmp45990 = s10 ? tmp45991 : tmp46007;
  assign tmp46016 = s7 ? tmp45994 : tmp46005;
  assign tmp46015 = s8 ? tmp46016 : tmp46001;
  assign tmp46014 = s9 ? tmp46008 : tmp46015;
  assign tmp46013 = s10 ? tmp45991 : tmp46014;
  assign tmp45989 = s11 ? tmp45990 : tmp46013;
  assign tmp46023 = s5 ? tmp44815 : tmp45996;
  assign tmp46022 = s6 ? tmp44809 : tmp46023;
  assign tmp46021 = s7 ? tmp43890 : tmp46022;
  assign tmp46020 = s8 ? tmp46021 : tmp46000;
  assign tmp46024 = s8 ? tmp46000 : tmp44721;
  assign tmp46019 = s9 ? tmp46020 : tmp46024;
  assign tmp46027 = s7 ? tmp46022 : tmp44796;
  assign tmp46026 = s8 ? tmp46027 : tmp46001;
  assign tmp46025 = s9 ? tmp46008 : tmp46026;
  assign tmp46018 = s10 ? tmp46019 : tmp46025;
  assign tmp46031 = s7 ? tmp46022 : tmp44722;
  assign tmp46030 = s8 ? tmp46031 : tmp46001;
  assign tmp46029 = s9 ? tmp46008 : tmp46030;
  assign tmp46028 = s10 ? tmp46019 : tmp46029;
  assign tmp46017 = s11 ? tmp46018 : tmp46028;
  assign tmp45988 = s12 ? tmp45989 : tmp46017;
  assign tmp45852 = s13 ? tmp45853 : tmp45988;
  assign tmp45797 = s14 ? tmp45798 : tmp45852;
  assign tmp46046 = l1 ? 1 : tmp44044;
  assign tmp46045 = s1 ? tmp46046 : tmp44166;
  assign tmp46047 = s1 ? tmp45281 : tmp44053;
  assign tmp46044 = ~(s2 ? tmp46045 : tmp46047);
  assign tmp46043 = s3 ? tmp45272 : tmp46044;
  assign tmp46050 = s1 ? tmp45286 : tmp45234;
  assign tmp46049 = s2 ? tmp46050 : tmp44017;
  assign tmp46048 = ~(s3 ? tmp46049 : tmp45289);
  assign tmp46042 = ~(s4 ? tmp46043 : tmp46048);
  assign tmp46041 = s5 ? tmp45236 : tmp46042;
  assign tmp46040 = s6 ? tmp45203 : tmp46041;
  assign tmp46039 = s7 ? tmp43890 : tmp46040;
  assign tmp46053 = s5 ? tmp45324 : tmp46042;
  assign tmp46052 = s6 ? tmp45295 : tmp46053;
  assign tmp46051 = s7 ? tmp43890 : tmp46052;
  assign tmp46038 = s8 ? tmp46039 : tmp46051;
  assign tmp46054 = s8 ? tmp46051 : tmp45293;
  assign tmp46037 = s9 ? tmp46038 : tmp46054;
  assign tmp46056 = s8 ? tmp46051 : tmp43890;
  assign tmp46060 = s5 ? tmp45355 : tmp46042;
  assign tmp46059 = s6 ? tmp45203 : tmp46060;
  assign tmp46058 = s7 ? tmp46059 : tmp45362;
  assign tmp46057 = s8 ? tmp46058 : tmp46052;
  assign tmp46055 = s9 ? tmp46056 : tmp46057;
  assign tmp46036 = s10 ? tmp46037 : tmp46055;
  assign tmp46064 = s7 ? tmp46040 : tmp45294;
  assign tmp46063 = s8 ? tmp46064 : tmp46052;
  assign tmp46062 = s9 ? tmp46056 : tmp46063;
  assign tmp46061 = s10 ? tmp46037 : tmp46062;
  assign tmp46035 = s11 ? tmp46036 : tmp46061;
  assign tmp46071 = s5 ? tmp45491 : tmp45439;
  assign tmp46070 = s6 ? tmp45463 : tmp46071;
  assign tmp46069 = s7 ? tmp43890 : tmp46070;
  assign tmp46068 = s8 ? tmp45372 : tmp46069;
  assign tmp46067 = s9 ? tmp46068 : tmp46069;
  assign tmp46073 = s8 ? tmp46069 : tmp43890;
  assign tmp46077 = s5 ? tmp45491 : tmp45529;
  assign tmp46076 = s6 ? tmp45463 : tmp46077;
  assign tmp46075 = s7 ? tmp45527 : tmp46076;
  assign tmp46074 = s8 ? tmp46075 : tmp46076;
  assign tmp46072 = s9 ? tmp46073 : tmp46074;
  assign tmp46066 = s10 ? tmp46067 : tmp46072;
  assign tmp46081 = s7 ? tmp45373 : tmp46070;
  assign tmp46080 = s8 ? tmp46081 : tmp46070;
  assign tmp46079 = s9 ? tmp46073 : tmp46080;
  assign tmp46078 = s10 ? tmp46067 : tmp46079;
  assign tmp46065 = s11 ? tmp46066 : tmp46078;
  assign tmp46034 = s12 ? tmp46035 : tmp46065;
  assign tmp46033 = s13 ? tmp46034 : tmp45534;
  assign tmp46032 = s14 ? tmp44830 : tmp46033;
  assign tmp45796 = s15 ? tmp45797 : tmp46032;
  assign tmp43881 = s16 ? tmp43882 : tmp45796;
  assign tmp46089 = s8 ? tmp45803 : tmp44215;
  assign tmp46088 = s9 ? tmp45802 : tmp46089;
  assign tmp46092 = s7 ? tmp45815 : tmp44216;
  assign tmp46091 = s8 ? tmp44268 : tmp46092;
  assign tmp46090 = s9 ? tmp44266 : tmp46091;
  assign tmp46087 = s10 ? tmp46088 : tmp46090;
  assign tmp46096 = s7 ? tmp45804 : tmp44216;
  assign tmp46095 = s8 ? tmp44280 : tmp46096;
  assign tmp46094 = s9 ? tmp44266 : tmp46095;
  assign tmp46093 = s10 ? tmp46088 : tmp46094;
  assign tmp46086 = s11 ? tmp46087 : tmp46093;
  assign tmp46101 = s8 ? tmp45831 : tmp44215;
  assign tmp46100 = s9 ? tmp45830 : tmp46101;
  assign tmp46104 = s7 ? tmp45845 : tmp44216;
  assign tmp46103 = s8 ? tmp44384 : tmp46104;
  assign tmp46102 = s9 ? tmp44266 : tmp46103;
  assign tmp46099 = s10 ? tmp46100 : tmp46102;
  assign tmp46108 = s7 ? tmp45832 : tmp44216;
  assign tmp46107 = s8 ? tmp44391 : tmp46108;
  assign tmp46106 = s9 ? tmp44266 : tmp46107;
  assign tmp46105 = s10 ? tmp46100 : tmp46106;
  assign tmp46098 = s11 ? tmp46099 : tmp46105;
  assign tmp46097 = s12 ? tmp44282 : tmp46098;
  assign tmp46085 = s13 ? tmp46086 : tmp46097;
  assign tmp46114 = s8 ? tmp45856 : tmp44453;
  assign tmp46113 = s9 ? tmp45856 : tmp46114;
  assign tmp46117 = s7 ? tmp45913 : tmp44454;
  assign tmp46116 = s8 ? tmp44470 : tmp46117;
  assign tmp46115 = s9 ? tmp44468 : tmp46116;
  assign tmp46112 = s10 ? tmp46113 : tmp46115;
  assign tmp46121 = s7 ? tmp45857 : tmp44454;
  assign tmp46120 = s8 ? tmp44479 : tmp46121;
  assign tmp46119 = s9 ? tmp44468 : tmp46120;
  assign tmp46118 = s10 ? tmp46113 : tmp46119;
  assign tmp46111 = s11 ? tmp46112 : tmp46118;
  assign tmp46125 = s8 ? tmp45925 : tmp44577;
  assign tmp46124 = s9 ? tmp45925 : tmp46125;
  assign tmp46127 = s7 ? tmp45980 : tmp44578;
  assign tmp46126 = s9 ? tmp44614 : tmp46127;
  assign tmp46123 = s10 ? tmp46124 : tmp46126;
  assign tmp46130 = s7 ? tmp45926 : tmp44578;
  assign tmp46129 = s9 ? tmp44614 : tmp46130;
  assign tmp46128 = s10 ? tmp46124 : tmp46129;
  assign tmp46122 = s11 ? tmp46123 : tmp46128;
  assign tmp46110 = s12 ? tmp46111 : tmp46122;
  assign tmp46135 = s8 ? tmp44630 : tmp46004;
  assign tmp46136 = s8 ? tmp46004 : tmp44721;
  assign tmp46134 = s9 ? tmp46135 : tmp46136;
  assign tmp46139 = s7 ? tmp46011 : tmp44796;
  assign tmp46138 = s8 ? tmp44790 : tmp46139;
  assign tmp46137 = s9 ? tmp44788 : tmp46138;
  assign tmp46133 = s10 ? tmp46134 : tmp46137;
  assign tmp46143 = s7 ? tmp46005 : tmp44722;
  assign tmp46142 = s8 ? tmp44802 : tmp46143;
  assign tmp46141 = s9 ? tmp44788 : tmp46142;
  assign tmp46140 = s10 ? tmp46134 : tmp46141;
  assign tmp46132 = s11 ? tmp46133 : tmp46140;
  assign tmp46131 = s12 ? tmp46132 : tmp44803;
  assign tmp46109 = s13 ? tmp46110 : tmp46131;
  assign tmp46084 = s14 ? tmp46085 : tmp46109;
  assign tmp46150 = s8 ? tmp46069 : tmp45461;
  assign tmp46149 = s9 ? tmp46068 : tmp46150;
  assign tmp46153 = s7 ? tmp46076 : tmp45462;
  assign tmp46152 = s8 ? tmp45526 : tmp46153;
  assign tmp46151 = s9 ? tmp45524 : tmp46152;
  assign tmp46148 = s10 ? tmp46149 : tmp46151;
  assign tmp46157 = s7 ? tmp46070 : tmp45462;
  assign tmp46156 = s8 ? tmp45533 : tmp46157;
  assign tmp46155 = s9 ? tmp45524 : tmp46156;
  assign tmp46154 = s10 ? tmp46149 : tmp46155;
  assign tmp46147 = s11 ? tmp46148 : tmp46154;
  assign tmp46146 = s12 ? tmp45197 : tmp46147;
  assign tmp46145 = s13 ? tmp46146 : tmp45534;
  assign tmp46144 = s14 ? tmp44830 : tmp46145;
  assign tmp46083 = s15 ? tmp46084 : tmp46144;
  assign tmp46164 = s9 ? tmp46135 : tmp46004;
  assign tmp46166 = s8 ? tmp46004 : tmp43890;
  assign tmp46168 = s7 ? tmp44791 : tmp46011;
  assign tmp46167 = s8 ? tmp46168 : tmp46011;
  assign tmp46165 = s9 ? tmp46166 : tmp46167;
  assign tmp46163 = s10 ? tmp46164 : tmp46165;
  assign tmp46172 = s7 ? tmp44631 : tmp46005;
  assign tmp46171 = s8 ? tmp46172 : tmp46005;
  assign tmp46170 = s9 ? tmp46166 : tmp46171;
  assign tmp46169 = s10 ? tmp46164 : tmp46170;
  assign tmp46162 = s11 ? tmp46163 : tmp46169;
  assign tmp46161 = s12 ? tmp46162 : tmp44803;
  assign tmp46160 = s13 ? tmp45853 : tmp46161;
  assign tmp46159 = s14 ? tmp45798 : tmp46160;
  assign tmp46175 = s12 ? tmp45197 : tmp46065;
  assign tmp46174 = s13 ? tmp46175 : tmp45534;
  assign tmp46173 = s14 ? tmp44830 : tmp46174;
  assign tmp46158 = s15 ? tmp46159 : tmp46173;
  assign tmp46082 = s16 ? tmp46083 : tmp46158;
  assign tmp43880 = ~(s17 ? tmp43881 : tmp46082);
  assign s0n = tmp43880;

  initial
   begin
    s0 = 0;
    s1 = 0;
    s2 = 0;
    s3 = 0;
    s4 = 0;
    s5 = 0;
    s6 = 0;
    s7 = 0;
    s8 = 0;
    s9 = 0;
    s10 = 0;
    s11 = 0;
    s12 = 0;
    s13 = 0;
    s14 = 0;
    s15 = 0;
    s16 = 0;
    s17 = 0;
    s18 = 0;
   end

  always @(posedge clock)
   begin
    s0 = s0n;
    s1 = s1n;
    s2 = s2n;
    s3 = s3n;
    s4 = s4n;
    s5 = s5n;
    s6 = s6n;
    s7 = s7n;
    s8 = s8n;
    s9 = s9n;
    s10 = s10n;
    s11 = s11n;
    s12 = s12n;
    s13 = s13n;
    s14 = s14n;
    s15 = s15n;
    s16 = s16n;
    s17 = s17n;
    s18 = s18n;
   end
endmodule



