/**************************************
* Simulation for inputfiles   
*   inputfiles/uav/map_8_states/map.dfa +                          
*   inputfiles/uav/map_8_states/adversary.dfa
***************************************/

module main;
  // Input of DUT:
  reg clk;
  reg l3;
  reg l2;
  reg l1;
  
  // Output of the DUT:
  wire l3__1;
  wire l2__1;
  wire l1__1;

  //Instantiate the DUT:
  shield s(clk, l1, l2, l3, l1__1, l2__1, l3__1);
  
  // make clock toggle:
  always #5 clk = ~clk;
  
  // Sequence of input stimuli to test with:
  initial begin
    clk = 0;

    l3 = 0;
    l2 = 0;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1);

    $display("Go around the building: 1 -> 2 -> 5 -> 6 -> 1");    

    //time=11 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 0;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d",  
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1);

    //time=21 -------------------------------------------------
    #9
    l3 = 1;
    l2 = 1;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d (Error by Design)",  
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1);
 
    //time=31 -------------------------------------------------
    #9
    l3 = 1;
    l2 = 0;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1);

    //time=61 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 0;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1); 

    $display("Go to loction 4 (on path of adversary) and stay there:");
    $display("    1 -> 4 -> 4 -> 1 -> 4 -> 1 -> 6");  

    //time=71 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 1;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d",  
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1);

    //time=81 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 1;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d (Error by Design)", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1); 

    //time=91 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 0;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1); 

    //time=101 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 1;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1); 

    //time=111 -------------------------------------------------
    #9
    l3 = 0;
    l2 = 0;
    l1 = 0;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1); 


    //time=121 -------------------------------------------------
    #9
    l3 = 1;
    l2 = 0;
    l1 = 1;
    #1
    $display("Time = %d, loc_design=%d%d%d, loc_shield=%d%d%d", 
             $time, 
             l3, l2, l1, l3__1, l2__1, l1__1); 

    #1 $finish;         
  end
endmodule


module shield(clock, l1, l2, l3, l1__1, l2__1, l3__1, recovery__1, recovery__2);
  input clock;
  input l1;
  input l2;
  input l3;
  output l1__1;
  output l2__1;
  output l3__1;
  output recovery__1;
  output recovery__2;

  wire s0n;
  wire s1n;
  wire s2n;
  wire s3n;
  wire s4n;
  wire s5n;
  wire s6n;
  wire s7n;
  wire s8n;
  wire s9n;
  wire s10n;
  wire s11n;
  wire s12n;
  wire s13n;
  wire s14n;
  wire s15n;
  wire s16n;
  wire tmp1;
  wire tmp2;
  wire tmp3;
  wire tmp4;
  wire tmp5;
  wire tmp6;
  wire tmp7;
  wire tmp8;
  wire tmp9;
  wire tmp10;
  wire tmp11;
  wire tmp12;
  wire tmp13;
  wire tmp14;
  wire tmp15;
  wire tmp16;
  wire tmp17;
  wire tmp18;
  wire tmp19;
  wire tmp20;
  wire tmp21;
  wire tmp22;
  wire tmp23;
  wire tmp24;
  wire tmp25;
  wire tmp26;
  wire tmp27;
  wire tmp28;
  wire tmp29;
  wire tmp30;
  wire tmp31;
  wire tmp32;
  wire tmp33;
  wire tmp34;
  wire tmp35;
  wire tmp36;
  wire tmp37;
  wire tmp38;
  wire tmp39;
  wire tmp40;
  wire tmp41;
  wire tmp42;
  wire tmp43;
  wire tmp44;
  wire tmp45;
  wire tmp46;
  wire tmp47;
  wire tmp48;
  wire tmp49;
  wire tmp50;
  wire tmp51;
  wire tmp52;
  wire tmp53;
  wire tmp54;
  wire tmp55;
  wire tmp56;
  wire tmp57;
  wire tmp58;
  wire tmp59;
  wire tmp60;
  wire tmp61;
  wire tmp62;
  wire tmp63;
  wire tmp64;
  wire tmp65;
  wire tmp66;
  wire tmp67;
  wire tmp68;
  wire tmp69;
  wire tmp70;
  wire tmp71;
  wire tmp72;
  wire tmp73;
  wire tmp74;
  wire tmp75;
  wire tmp76;
  wire tmp77;
  wire tmp78;
  wire tmp79;
  wire tmp80;
  wire tmp81;
  wire tmp82;
  wire tmp83;
  wire tmp84;
  wire tmp85;
  wire tmp86;
  wire tmp87;
  wire tmp88;
  wire tmp89;
  wire tmp90;
  wire tmp91;
  wire tmp92;
  wire tmp93;
  wire tmp94;
  wire tmp95;
  wire tmp96;
  wire tmp97;
  wire tmp98;
  wire tmp99;
  wire tmp100;
  wire tmp101;
  wire tmp102;
  wire tmp103;
  wire tmp104;
  wire tmp105;
  wire tmp106;
  wire tmp107;
  wire tmp108;
  wire tmp109;
  wire tmp110;
  wire tmp111;
  wire tmp112;
  wire tmp113;
  wire tmp114;
  wire tmp115;
  wire tmp116;
  wire tmp117;
  wire tmp118;
  wire tmp119;
  wire tmp120;
  wire tmp121;
  wire tmp122;
  wire tmp123;
  wire tmp124;
  wire tmp125;
  wire tmp126;
  wire tmp127;
  wire tmp128;
  wire tmp129;
  wire tmp130;
  wire tmp131;
  wire tmp132;
  wire tmp133;
  wire tmp134;
  wire tmp135;
  wire tmp136;
  wire tmp137;
  wire tmp138;
  wire tmp139;
  wire tmp140;
  wire tmp141;
  wire tmp142;
  wire tmp143;
  wire tmp144;
  wire tmp145;
  wire tmp146;
  wire tmp147;
  wire tmp148;
  wire tmp149;
  wire tmp150;
  wire tmp151;
  wire tmp152;
  wire tmp153;
  wire tmp154;
  wire tmp155;
  wire tmp156;
  wire tmp157;
  wire tmp158;
  wire tmp159;
  wire tmp160;
  wire tmp161;
  wire tmp162;
  wire tmp163;
  wire tmp164;
  wire tmp165;
  wire tmp166;
  wire tmp167;
  wire tmp168;
  wire tmp169;
  wire tmp170;
  wire tmp171;
  wire tmp172;
  wire tmp173;
  wire tmp174;
  wire tmp175;
  wire tmp176;
  wire tmp177;
  wire tmp178;
  wire tmp179;
  wire tmp180;
  wire tmp181;
  wire tmp182;
  wire tmp183;
  wire tmp184;
  wire tmp185;
  wire tmp186;
  wire tmp187;
  wire tmp188;
  wire tmp189;
  wire tmp190;
  wire tmp191;
  wire tmp192;
  wire tmp193;
  wire tmp194;
  wire tmp195;
  wire tmp196;
  wire tmp197;
  wire tmp198;
  wire tmp199;
  wire tmp200;
  wire tmp201;
  wire tmp202;
  wire tmp203;
  wire tmp204;
  wire tmp205;
  wire tmp206;
  wire tmp207;
  wire tmp208;
  wire tmp209;
  wire tmp210;
  wire tmp211;
  wire tmp212;
  wire tmp213;
  wire tmp214;
  wire tmp215;
  wire tmp216;
  wire tmp217;
  wire tmp218;
  wire tmp219;
  wire tmp220;
  wire tmp221;
  wire tmp222;
  wire tmp223;
  wire tmp224;
  wire tmp225;
  wire tmp226;
  wire tmp227;
  wire tmp228;
  wire tmp229;
  wire tmp230;
  wire tmp231;
  wire tmp232;
  wire tmp233;
  wire tmp234;
  wire tmp235;
  wire tmp236;
  wire tmp237;
  wire tmp238;
  wire tmp239;
  wire tmp240;
  wire tmp241;
  wire tmp242;
  wire tmp243;
  wire tmp244;
  wire tmp245;
  wire tmp246;
  wire tmp247;
  wire tmp248;
  wire tmp249;
  wire tmp250;
  wire tmp251;
  wire tmp252;
  wire tmp253;
  wire tmp254;
  wire tmp255;
  wire tmp256;
  wire tmp257;
  wire tmp258;
  wire tmp259;
  wire tmp260;
  wire tmp261;
  wire tmp262;
  wire tmp263;
  wire tmp264;
  wire tmp265;
  wire tmp266;
  wire tmp267;
  wire tmp268;
  wire tmp269;
  wire tmp270;
  wire tmp271;
  wire tmp272;
  wire tmp273;
  wire tmp274;
  wire tmp275;
  wire tmp276;
  wire tmp277;
  wire tmp278;
  wire tmp279;
  wire tmp280;
  wire tmp281;
  wire tmp282;
  wire tmp283;
  wire tmp284;
  wire tmp285;
  wire tmp286;
  wire tmp287;
  wire tmp288;
  wire tmp289;
  wire tmp290;
  wire tmp291;
  wire tmp292;
  wire tmp293;
  wire tmp294;
  wire tmp295;
  wire tmp296;
  wire tmp297;
  wire tmp298;
  wire tmp299;
  wire tmp300;
  wire tmp301;
  wire tmp302;
  wire tmp303;
  wire tmp304;
  wire tmp305;
  wire tmp306;
  wire tmp307;
  wire tmp308;
  wire tmp309;
  wire tmp310;
  wire tmp311;
  wire tmp312;
  wire tmp313;
  wire tmp314;
  wire tmp315;
  wire tmp316;
  wire tmp317;
  wire tmp318;
  wire tmp319;
  wire tmp320;
  wire tmp321;
  wire tmp322;
  wire tmp323;
  wire tmp324;
  wire tmp325;
  wire tmp326;
  wire tmp327;
  wire tmp328;
  wire tmp329;
  wire tmp330;
  wire tmp331;
  wire tmp332;
  wire tmp333;
  wire tmp334;
  wire tmp335;
  wire tmp336;
  wire tmp337;
  wire tmp338;
  wire tmp339;
  wire tmp340;
  wire tmp341;
  wire tmp342;
  wire tmp343;
  wire tmp344;
  wire tmp345;
  wire tmp346;
  wire tmp347;
  wire tmp348;
  wire tmp349;
  wire tmp350;
  wire tmp351;
  wire tmp352;
  wire tmp353;
  wire tmp354;
  wire tmp355;
  wire tmp356;
  wire tmp357;
  wire tmp358;
  wire tmp359;
  wire tmp360;
  wire tmp361;
  wire tmp362;
  wire tmp363;
  wire tmp364;
  wire tmp365;
  wire tmp366;
  wire tmp367;
  wire tmp368;
  wire tmp369;
  wire tmp370;
  wire tmp371;
  wire tmp372;
  wire tmp373;
  wire tmp374;
  wire tmp375;
  wire tmp376;
  wire tmp377;
  wire tmp378;
  wire tmp379;
  wire tmp380;
  wire tmp381;
  wire tmp382;
  wire tmp383;
  wire tmp384;
  wire tmp385;
  wire tmp386;
  wire tmp387;
  wire tmp388;
  wire tmp389;
  wire tmp390;
  wire tmp391;
  wire tmp392;
  wire tmp393;
  wire tmp394;
  wire tmp395;
  wire tmp396;
  wire tmp397;
  wire tmp398;
  wire tmp399;
  wire tmp400;
  wire tmp401;
  wire tmp402;
  wire tmp403;
  wire tmp404;
  wire tmp405;
  wire tmp406;
  wire tmp407;
  wire tmp408;
  wire tmp409;
  wire tmp410;
  wire tmp411;
  wire tmp412;
  wire tmp413;
  wire tmp414;
  wire tmp415;
  wire tmp416;
  wire tmp417;
  wire tmp418;
  wire tmp419;
  wire tmp420;
  wire tmp421;
  wire tmp422;
  wire tmp423;
  wire tmp424;
  wire tmp425;
  wire tmp426;
  wire tmp427;
  wire tmp428;
  wire tmp429;
  wire tmp430;
  wire tmp431;
  wire tmp432;
  wire tmp433;
  wire tmp434;
  wire tmp435;
  wire tmp436;
  wire tmp437;
  wire tmp438;
  wire tmp439;
  wire tmp440;
  wire tmp441;
  wire tmp442;
  wire tmp443;
  wire tmp444;
  wire tmp445;
  wire tmp446;
  wire tmp447;
  wire tmp448;
  wire tmp449;
  wire tmp450;
  wire tmp451;
  wire tmp452;
  wire tmp453;
  wire tmp454;
  wire tmp455;
  wire tmp456;
  wire tmp457;
  wire tmp458;
  wire tmp459;
  wire tmp460;
  wire tmp461;
  wire tmp462;
  wire tmp463;
  wire tmp464;
  wire tmp465;
  wire tmp466;
  wire tmp467;
  wire tmp468;
  wire tmp469;
  wire tmp470;
  wire tmp471;
  wire tmp472;
  wire tmp473;
  wire tmp474;
  wire tmp475;
  wire tmp476;
  wire tmp477;
  wire tmp478;
  wire tmp479;
  wire tmp480;
  wire tmp481;
  wire tmp482;
  wire tmp483;
  wire tmp484;
  wire tmp485;
  wire tmp486;
  wire tmp487;
  wire tmp488;
  wire tmp489;
  wire tmp490;
  wire tmp491;
  wire tmp492;
  wire tmp493;
  wire tmp494;
  wire tmp495;
  wire tmp496;
  wire tmp497;
  wire tmp498;
  wire tmp499;
  wire tmp500;
  wire tmp501;
  wire tmp502;
  wire tmp503;
  wire tmp504;
  wire tmp505;
  wire tmp506;
  wire tmp507;
  wire tmp508;
  wire tmp509;
  wire tmp510;
  wire tmp511;
  wire tmp512;
  wire tmp513;
  wire tmp514;
  wire tmp515;
  wire tmp516;
  wire tmp517;
  wire tmp518;
  wire tmp519;
  wire tmp520;
  wire tmp521;
  wire tmp522;
  wire tmp523;
  wire tmp524;
  wire tmp525;
  wire tmp526;
  wire tmp527;
  wire tmp528;
  wire tmp529;
  wire tmp530;
  wire tmp531;
  wire tmp532;
  wire tmp533;
  wire tmp534;
  wire tmp535;
  wire tmp536;
  wire tmp537;
  wire tmp538;
  wire tmp539;
  wire tmp540;
  wire tmp541;
  wire tmp542;
  wire tmp543;
  wire tmp544;
  wire tmp545;
  wire tmp546;
  wire tmp547;
  wire tmp548;
  wire tmp549;
  wire tmp550;
  wire tmp551;
  wire tmp552;
  wire tmp553;
  wire tmp554;
  wire tmp555;
  wire tmp556;
  wire tmp557;
  wire tmp558;
  wire tmp559;
  wire tmp560;
  wire tmp561;
  wire tmp562;
  wire tmp563;
  wire tmp564;
  wire tmp565;
  wire tmp566;
  wire tmp567;
  wire tmp568;
  wire tmp569;
  wire tmp570;
  wire tmp571;
  wire tmp572;
  wire tmp573;
  wire tmp574;
  wire tmp575;
  wire tmp576;
  wire tmp577;
  wire tmp578;
  wire tmp579;
  wire tmp580;
  wire tmp581;
  wire tmp582;
  wire tmp583;
  wire tmp584;
  wire tmp585;
  wire tmp586;
  wire tmp587;
  wire tmp588;
  wire tmp589;
  wire tmp590;
  wire tmp591;
  wire tmp592;
  wire tmp593;
  wire tmp594;
  wire tmp595;
  wire tmp596;
  wire tmp597;
  wire tmp598;
  wire tmp599;
  wire tmp600;
  wire tmp601;
  wire tmp602;
  wire tmp603;
  wire tmp604;
  wire tmp605;
  wire tmp606;
  wire tmp607;
  wire tmp608;
  wire tmp609;
  wire tmp610;
  wire tmp611;
  wire tmp612;
  wire tmp613;
  wire tmp614;
  wire tmp615;
  wire tmp616;
  wire tmp617;
  wire tmp618;
  wire tmp619;
  wire tmp620;
  wire tmp621;
  wire tmp622;
  wire tmp623;
  wire tmp624;
  wire tmp625;
  wire tmp626;
  wire tmp627;
  wire tmp628;
  wire tmp629;
  wire tmp630;
  wire tmp631;
  wire tmp632;
  wire tmp633;
  wire tmp634;
  wire tmp635;
  wire tmp636;
  wire tmp637;
  wire tmp638;
  wire tmp639;
  wire tmp640;
  wire tmp641;
  wire tmp642;
  wire tmp643;
  wire tmp644;
  wire tmp645;
  wire tmp646;
  wire tmp647;
  wire tmp648;
  wire tmp649;
  wire tmp650;
  wire tmp651;
  wire tmp652;
  wire tmp653;
  wire tmp654;
  wire tmp655;
  wire tmp656;
  wire tmp657;
  wire tmp658;
  wire tmp659;
  wire tmp660;
  wire tmp661;
  wire tmp662;
  wire tmp663;
  wire tmp664;
  wire tmp665;
  wire tmp666;
  wire tmp667;
  wire tmp668;
  wire tmp669;
  wire tmp670;
  wire tmp671;
  wire tmp672;
  wire tmp673;
  wire tmp674;
  wire tmp675;
  wire tmp676;
  wire tmp677;
  wire tmp678;
  wire tmp679;
  wire tmp680;
  wire tmp681;
  wire tmp682;
  wire tmp683;
  wire tmp684;
  wire tmp685;
  wire tmp686;
  wire tmp687;
  wire tmp688;
  wire tmp689;
  wire tmp690;
  wire tmp691;
  wire tmp692;
  wire tmp693;
  wire tmp694;
  wire tmp695;
  wire tmp696;
  wire tmp697;
  wire tmp698;
  wire tmp699;
  wire tmp700;
  wire tmp701;
  wire tmp702;
  wire tmp703;
  wire tmp704;
  wire tmp705;
  wire tmp706;
  wire tmp707;
  wire tmp708;
  wire tmp709;
  wire tmp710;
  wire tmp711;
  wire tmp712;
  wire tmp713;
  wire tmp714;
  wire tmp715;
  wire tmp716;
  wire tmp717;
  wire tmp718;
  wire tmp719;
  wire tmp720;
  wire tmp721;
  wire tmp722;
  wire tmp723;
  wire tmp724;
  wire tmp725;
  wire tmp726;
  wire tmp727;
  wire tmp728;
  wire tmp729;
  wire tmp730;
  wire tmp731;
  wire tmp732;
  wire tmp733;
  wire tmp734;
  wire tmp735;
  wire tmp736;
  wire tmp737;
  wire tmp738;
  wire tmp739;
  wire tmp740;
  wire tmp741;
  wire tmp742;
  wire tmp743;
  wire tmp744;
  wire tmp745;
  wire tmp746;
  wire tmp747;
  wire tmp748;
  wire tmp749;
  wire tmp750;
  wire tmp751;
  wire tmp752;
  wire tmp753;
  wire tmp754;
  wire tmp755;
  wire tmp756;
  wire tmp757;
  wire tmp758;
  wire tmp759;
  wire tmp760;
  wire tmp761;
  wire tmp762;
  wire tmp763;
  wire tmp764;
  wire tmp765;
  wire tmp766;
  wire tmp767;
  wire tmp768;
  wire tmp769;
  wire tmp770;
  wire tmp771;
  wire tmp772;
  wire tmp773;
  wire tmp774;
  wire tmp775;
  wire tmp776;
  wire tmp777;
  wire tmp778;
  wire tmp779;
  wire tmp780;
  wire tmp781;
  wire tmp782;
  wire tmp783;
  wire tmp784;
  wire tmp785;
  wire tmp786;
  wire tmp787;
  wire tmp788;
  wire tmp789;
  wire tmp790;
  wire tmp791;
  wire tmp792;
  wire tmp793;
  wire tmp794;
  wire tmp795;
  wire tmp796;
  wire tmp797;
  wire tmp798;
  wire tmp799;
  wire tmp800;
  wire tmp801;
  wire tmp802;
  wire tmp803;
  wire tmp804;
  wire tmp805;
  wire tmp806;
  wire tmp807;
  wire tmp808;
  wire tmp809;
  wire tmp810;
  wire tmp811;
  wire tmp812;
  wire tmp813;
  wire tmp814;
  wire tmp815;
  wire tmp816;
  wire tmp817;
  wire tmp818;
  wire tmp819;
  wire tmp820;
  wire tmp821;
  wire tmp822;
  wire tmp823;
  wire tmp824;
  wire tmp825;
  wire tmp826;
  wire tmp827;
  wire tmp828;
  wire tmp829;
  wire tmp830;
  wire tmp831;
  wire tmp832;
  wire tmp833;
  wire tmp834;
  wire tmp835;
  wire tmp836;
  wire tmp837;
  wire tmp838;
  wire tmp839;
  wire tmp840;
  wire tmp841;
  wire tmp842;
  wire tmp843;
  wire tmp844;
  wire tmp845;
  wire tmp846;
  wire tmp847;
  wire tmp848;
  wire tmp849;
  wire tmp850;
  wire tmp851;
  wire tmp852;
  wire tmp853;
  wire tmp854;
  wire tmp855;
  wire tmp856;
  wire tmp857;
  wire tmp858;
  wire tmp859;
  wire tmp860;
  wire tmp861;
  wire tmp862;
  wire tmp863;
  wire tmp864;
  wire tmp865;
  wire tmp866;
  wire tmp867;
  wire tmp868;
  wire tmp869;
  wire tmp870;
  wire tmp871;
  wire tmp872;
  wire tmp873;
  wire tmp874;
  wire tmp875;
  wire tmp876;
  wire tmp877;
  wire tmp878;
  wire tmp879;
  wire tmp880;
  wire tmp881;
  wire tmp882;
  wire tmp883;
  wire tmp884;
  wire tmp885;
  wire tmp886;
  wire tmp887;
  wire tmp888;
  wire tmp889;
  wire tmp890;
  wire tmp891;
  wire tmp892;
  wire tmp893;
  wire tmp894;
  wire tmp895;
  wire tmp896;
  wire tmp897;
  wire tmp898;
  wire tmp899;
  wire tmp900;
  wire tmp901;
  wire tmp902;
  wire tmp903;
  wire tmp904;
  wire tmp905;
  wire tmp906;
  wire tmp907;
  wire tmp908;
  wire tmp909;
  wire tmp910;
  wire tmp911;
  wire tmp912;
  wire tmp913;
  wire tmp914;
  wire tmp915;
  wire tmp916;
  wire tmp917;
  wire tmp918;
  wire tmp919;
  wire tmp920;
  wire tmp921;
  wire tmp922;
  wire tmp923;
  wire tmp924;
  wire tmp925;
  wire tmp926;
  wire tmp927;
  wire tmp928;
  wire tmp929;
  wire tmp930;
  wire tmp931;
  wire tmp932;
  wire tmp933;
  wire tmp934;
  wire tmp935;
  wire tmp936;
  wire tmp937;
  wire tmp938;
  wire tmp939;
  wire tmp940;
  wire tmp941;
  wire tmp942;
  wire tmp943;
  wire tmp944;
  wire tmp945;
  wire tmp946;
  wire tmp947;
  wire tmp948;
  wire tmp949;
  wire tmp950;
  wire tmp951;
  wire tmp952;
  wire tmp953;
  wire tmp954;
  wire tmp955;
  wire tmp956;
  wire tmp957;
  wire tmp958;
  wire tmp959;
  wire tmp960;
  wire tmp961;
  wire tmp962;
  wire tmp963;
  wire tmp964;
  wire tmp965;
  wire tmp966;
  wire tmp967;
  wire tmp968;
  wire tmp969;
  wire tmp970;
  wire tmp971;
  wire tmp972;
  wire tmp973;
  wire tmp974;
  wire tmp975;
  wire tmp976;
  wire tmp977;
  wire tmp978;
  wire tmp979;
  wire tmp980;
  wire tmp981;
  wire tmp982;
  wire tmp983;
  wire tmp984;
  wire tmp985;
  wire tmp986;
  wire tmp987;
  wire tmp988;
  wire tmp989;
  wire tmp990;
  wire tmp991;
  wire tmp992;
  wire tmp993;
  wire tmp994;
  wire tmp995;
  wire tmp996;
  wire tmp997;
  wire tmp998;
  wire tmp999;
  wire tmp1000;
  wire tmp1001;
  wire tmp1002;
  wire tmp1003;
  wire tmp1004;
  wire tmp1005;
  wire tmp1006;
  wire tmp1007;
  wire tmp1008;
  wire tmp1009;
  wire tmp1010;
  wire tmp1011;
  wire tmp1012;
  wire tmp1013;
  wire tmp1014;
  wire tmp1015;
  wire tmp1016;
  wire tmp1017;
  wire tmp1018;
  wire tmp1019;
  wire tmp1020;
  wire tmp1021;
  wire tmp1022;
  wire tmp1023;
  wire tmp1024;
  wire tmp1025;
  wire tmp1026;
  wire tmp1027;
  wire tmp1028;
  wire tmp1029;
  wire tmp1030;
  wire tmp1031;
  wire tmp1032;
  wire tmp1033;
  wire tmp1034;
  wire tmp1035;
  wire tmp1036;
  wire tmp1037;
  wire tmp1038;
  wire tmp1039;
  wire tmp1040;
  wire tmp1041;
  wire tmp1042;
  wire tmp1043;
  wire tmp1044;
  wire tmp1045;
  wire tmp1046;
  wire tmp1047;
  wire tmp1048;
  wire tmp1049;
  wire tmp1050;
  wire tmp1051;
  wire tmp1052;
  wire tmp1053;
  wire tmp1054;
  wire tmp1055;
  wire tmp1056;
  wire tmp1057;
  wire tmp1058;
  wire tmp1059;
  wire tmp1060;
  wire tmp1061;
  wire tmp1062;
  wire tmp1063;
  wire tmp1064;
  wire tmp1065;
  wire tmp1066;
  wire tmp1067;
  wire tmp1068;
  wire tmp1069;
  wire tmp1070;
  wire tmp1071;
  wire tmp1072;
  wire tmp1073;
  wire tmp1074;
  wire tmp1075;
  wire tmp1076;
  wire tmp1077;
  wire tmp1078;
  wire tmp1079;
  wire tmp1080;
  wire tmp1081;
  wire tmp1082;
  wire tmp1083;
  wire tmp1084;
  wire tmp1085;
  wire tmp1086;
  wire tmp1087;
  wire tmp1088;
  wire tmp1089;
  wire tmp1090;
  wire tmp1091;
  wire tmp1092;
  wire tmp1093;
  wire tmp1094;
  wire tmp1095;
  wire tmp1096;
  wire tmp1097;
  wire tmp1098;
  wire tmp1099;
  wire tmp1100;
  wire tmp1101;
  wire tmp1102;
  wire tmp1103;
  wire tmp1104;
  wire tmp1105;
  wire tmp1106;
  wire tmp1107;
  wire tmp1108;
  wire tmp1109;
  wire tmp1110;
  wire tmp1111;
  wire tmp1112;
  wire tmp1113;
  wire tmp1114;
  wire tmp1115;
  wire tmp1116;
  wire tmp1117;
  wire tmp1118;
  wire tmp1119;
  wire tmp1120;
  wire tmp1121;
  wire tmp1122;
  wire tmp1123;
  wire tmp1124;
  wire tmp1125;
  wire tmp1126;
  wire tmp1127;
  wire tmp1128;
  wire tmp1129;
  wire tmp1130;
  wire tmp1131;
  wire tmp1132;
  wire tmp1133;
  wire tmp1134;
  wire tmp1135;
  wire tmp1136;
  wire tmp1137;
  wire tmp1138;
  wire tmp1139;
  wire tmp1140;
  wire tmp1141;
  wire tmp1142;
  wire tmp1143;
  wire tmp1144;
  wire tmp1145;
  wire tmp1146;
  wire tmp1147;
  wire tmp1148;
  wire tmp1149;
  wire tmp1150;
  wire tmp1151;
  wire tmp1152;
  wire tmp1153;
  wire tmp1154;
  wire tmp1155;
  wire tmp1156;
  wire tmp1157;
  wire tmp1158;
  wire tmp1159;
  wire tmp1160;
  wire tmp1161;
  wire tmp1162;
  wire tmp1163;
  wire tmp1164;
  wire tmp1165;
  wire tmp1166;
  wire tmp1167;
  wire tmp1168;
  wire tmp1169;
  wire tmp1170;
  wire tmp1171;
  wire tmp1172;
  wire tmp1173;
  wire tmp1174;
  wire tmp1175;
  wire tmp1176;
  wire tmp1177;
  wire tmp1178;
  wire tmp1179;
  wire tmp1180;
  wire tmp1181;
  wire tmp1182;
  wire tmp1183;
  wire tmp1184;
  wire tmp1185;
  wire tmp1186;
  wire tmp1187;
  wire tmp1188;
  wire tmp1189;
  wire tmp1190;
  wire tmp1191;
  wire tmp1192;
  wire tmp1193;
  wire tmp1194;
  wire tmp1195;
  wire tmp1196;
  wire tmp1197;
  wire tmp1198;
  wire tmp1199;
  wire tmp1200;
  wire tmp1201;
  wire tmp1202;
  wire tmp1203;
  wire tmp1204;
  wire tmp1205;
  wire tmp1206;
  wire tmp1207;
  wire tmp1208;
  wire tmp1209;
  wire tmp1210;
  wire tmp1211;
  wire tmp1212;
  wire tmp1213;
  wire tmp1214;
  wire tmp1215;
  wire tmp1216;
  wire tmp1217;
  wire tmp1218;
  wire tmp1219;
  wire tmp1220;
  wire tmp1221;
  wire tmp1222;
  wire tmp1223;
  wire tmp1224;
  wire tmp1225;
  wire tmp1226;
  wire tmp1227;
  wire tmp1228;
  wire tmp1229;
  wire tmp1230;
  wire tmp1231;
  wire tmp1232;
  wire tmp1233;
  wire tmp1234;
  wire tmp1235;
  wire tmp1236;
  wire tmp1237;
  wire tmp1238;
  wire tmp1239;
  wire tmp1240;
  wire tmp1241;
  wire tmp1242;
  wire tmp1243;
  wire tmp1244;
  wire tmp1245;
  wire tmp1246;
  wire tmp1247;
  wire tmp1248;
  wire tmp1249;
  wire tmp1250;
  wire tmp1251;
  wire tmp1252;
  wire tmp1253;
  wire tmp1254;
  wire tmp1255;
  wire tmp1256;
  wire tmp1257;
  wire tmp1258;
  wire tmp1259;
  wire tmp1260;
  wire tmp1261;
  wire tmp1262;
  wire tmp1263;
  wire tmp1264;
  wire tmp1265;
  wire tmp1266;
  wire tmp1267;
  wire tmp1268;
  wire tmp1269;
  wire tmp1270;
  wire tmp1271;
  wire tmp1272;
  wire tmp1273;
  wire tmp1274;
  wire tmp1275;
  wire tmp1276;
  wire tmp1277;
  wire tmp1278;
  wire tmp1279;
  wire tmp1280;
  wire tmp1281;
  wire tmp1282;
  wire tmp1283;
  wire tmp1284;
  wire tmp1285;
  wire tmp1286;
  wire tmp1287;
  wire tmp1288;
  wire tmp1289;
  wire tmp1290;
  wire tmp1291;
  wire tmp1292;
  wire tmp1293;
  wire tmp1294;
  wire tmp1295;
  wire tmp1296;
  wire tmp1297;
  wire tmp1298;
  wire tmp1299;
  wire tmp1300;
  wire tmp1301;
  wire tmp1302;
  wire tmp1303;
  wire tmp1304;
  wire tmp1305;
  wire tmp1306;
  wire tmp1307;
  wire tmp1308;
  wire tmp1309;
  wire tmp1310;
  wire tmp1311;
  wire tmp1312;
  wire tmp1313;
  wire tmp1314;
  wire tmp1315;
  wire tmp1316;
  wire tmp1317;
  wire tmp1318;
  wire tmp1319;
  wire tmp1320;
  wire tmp1321;
  wire tmp1322;
  wire tmp1323;
  wire tmp1324;
  wire tmp1325;
  wire tmp1326;
  wire tmp1327;
  wire tmp1328;
  wire tmp1329;
  wire tmp1330;
  wire tmp1331;
  wire tmp1332;
  wire tmp1333;
  wire tmp1334;
  wire tmp1335;
  wire tmp1336;
  wire tmp1337;
  wire tmp1338;
  wire tmp1339;
  wire tmp1340;
  wire tmp1341;
  wire tmp1342;
  wire tmp1343;
  wire tmp1344;
  wire tmp1345;
  wire tmp1346;
  wire tmp1347;
  wire tmp1348;
  wire tmp1349;
  wire tmp1350;
  wire tmp1351;
  wire tmp1352;
  wire tmp1353;
  wire tmp1354;
  wire tmp1355;
  wire tmp1356;
  wire tmp1357;
  wire tmp1358;
  wire tmp1359;
  wire tmp1360;
  wire tmp1361;
  wire tmp1362;
  wire tmp1363;
  wire tmp1364;
  wire tmp1365;
  wire tmp1366;
  wire tmp1367;
  wire tmp1368;
  wire tmp1369;
  wire tmp1370;
  wire tmp1371;
  wire tmp1372;
  wire tmp1373;
  wire tmp1374;
  wire tmp1375;
  wire tmp1376;
  wire tmp1377;
  wire tmp1378;
  wire tmp1379;
  wire tmp1380;
  wire tmp1381;
  wire tmp1382;
  wire tmp1383;
  wire tmp1384;
  wire tmp1385;
  wire tmp1386;
  wire tmp1387;
  wire tmp1388;
  wire tmp1389;
  wire tmp1390;
  wire tmp1391;
  wire tmp1392;
  wire tmp1393;
  wire tmp1394;
  wire tmp1395;
  wire tmp1396;
  wire tmp1397;
  wire tmp1398;
  wire tmp1399;
  wire tmp1400;
  wire tmp1401;
  wire tmp1402;
  wire tmp1403;
  wire tmp1404;
  wire tmp1405;
  wire tmp1406;
  wire tmp1407;
  wire tmp1408;
  wire tmp1409;
  wire tmp1410;
  wire tmp1411;
  wire tmp1412;
  wire tmp1413;
  wire tmp1414;
  wire tmp1415;
  wire tmp1416;
  wire tmp1417;
  wire tmp1418;
  wire tmp1419;
  wire tmp1420;
  wire tmp1421;
  wire tmp1422;
  wire tmp1423;
  wire tmp1424;
  wire tmp1425;
  wire tmp1426;
  wire tmp1427;
  wire tmp1428;
  wire tmp1429;
  wire tmp1430;
  wire tmp1431;
  wire tmp1432;
  wire tmp1433;
  wire tmp1434;
  wire tmp1435;
  wire tmp1436;
  wire tmp1437;
  wire tmp1438;
  wire tmp1439;
  wire tmp1440;
  wire tmp1441;
  wire tmp1442;
  wire tmp1443;
  wire tmp1444;
  wire tmp1445;
  wire tmp1446;
  wire tmp1447;
  wire tmp1448;
  wire tmp1449;
  wire tmp1450;
  wire tmp1451;
  wire tmp1452;
  wire tmp1453;
  wire tmp1454;
  wire tmp1455;
  wire tmp1456;
  wire tmp1457;
  wire tmp1458;
  wire tmp1459;
  wire tmp1460;
  wire tmp1461;
  wire tmp1462;
  wire tmp1463;
  wire tmp1464;
  wire tmp1465;
  wire tmp1466;
  wire tmp1467;
  wire tmp1468;
  wire tmp1469;
  wire tmp1470;
  wire tmp1471;
  wire tmp1472;
  wire tmp1473;
  wire tmp1474;
  wire tmp1475;
  wire tmp1476;
  wire tmp1477;
  wire tmp1478;
  wire tmp1479;
  wire tmp1480;
  wire tmp1481;
  wire tmp1482;
  wire tmp1483;
  wire tmp1484;
  wire tmp1485;
  wire tmp1486;
  wire tmp1487;
  wire tmp1488;
  wire tmp1489;
  wire tmp1490;
  wire tmp1491;
  wire tmp1492;
  wire tmp1493;
  wire tmp1494;
  wire tmp1495;
  wire tmp1496;
  wire tmp1497;
  wire tmp1498;
  wire tmp1499;
  wire tmp1500;
  wire tmp1501;
  wire tmp1502;
  wire tmp1503;
  wire tmp1504;
  wire tmp1505;
  wire tmp1506;
  wire tmp1507;
  wire tmp1508;
  wire tmp1509;
  wire tmp1510;
  wire tmp1511;
  wire tmp1512;
  wire tmp1513;
  wire tmp1514;
  wire tmp1515;
  wire tmp1516;
  wire tmp1517;
  wire tmp1518;
  wire tmp1519;
  wire tmp1520;
  wire tmp1521;
  wire tmp1522;
  wire tmp1523;
  wire tmp1524;
  wire tmp1525;
  wire tmp1526;
  wire tmp1527;
  wire tmp1528;
  wire tmp1529;
  wire tmp1530;
  wire tmp1531;
  wire tmp1532;
  wire tmp1533;
  wire tmp1534;
  wire tmp1535;
  wire tmp1536;
  wire tmp1537;
  wire tmp1538;
  wire tmp1539;
  wire tmp1540;
  wire tmp1541;
  wire tmp1542;
  wire tmp1543;
  wire tmp1544;
  wire tmp1545;
  wire tmp1546;
  wire tmp1547;
  wire tmp1548;
  wire tmp1549;
  wire tmp1550;
  wire tmp1551;
  wire tmp1552;
  wire tmp1553;
  wire tmp1554;
  wire tmp1555;
  wire tmp1556;
  wire tmp1557;
  wire tmp1558;
  wire tmp1559;
  wire tmp1560;
  wire tmp1561;
  wire tmp1562;
  wire tmp1563;
  wire tmp1564;
  wire tmp1565;
  wire tmp1566;
  wire tmp1567;
  wire tmp1568;
  wire tmp1569;
  wire tmp1570;
  wire tmp1571;
  wire tmp1572;
  wire tmp1573;
  wire tmp1574;
  wire tmp1575;
  wire tmp1576;
  wire tmp1577;
  wire tmp1578;
  wire tmp1579;
  wire tmp1580;
  wire tmp1581;
  wire tmp1582;
  wire tmp1583;
  wire tmp1584;
  wire tmp1585;
  wire tmp1586;
  wire tmp1587;
  wire tmp1588;
  wire tmp1589;
  wire tmp1590;
  wire tmp1591;
  wire tmp1592;
  wire tmp1593;
  wire tmp1594;
  wire tmp1595;
  wire tmp1596;
  wire tmp1597;
  wire tmp1598;
  wire tmp1599;
  wire tmp1600;
  wire tmp1601;
  wire tmp1602;
  wire tmp1603;
  wire tmp1604;
  wire tmp1605;
  wire tmp1606;
  wire tmp1607;
  wire tmp1608;
  wire tmp1609;
  wire tmp1610;
  wire tmp1611;
  wire tmp1612;
  wire tmp1613;
  wire tmp1614;
  wire tmp1615;
  wire tmp1616;
  wire tmp1617;
  wire tmp1618;
  wire tmp1619;
  wire tmp1620;
  wire tmp1621;
  wire tmp1622;
  wire tmp1623;
  wire tmp1624;
  wire tmp1625;
  wire tmp1626;
  wire tmp1627;
  wire tmp1628;
  wire tmp1629;
  wire tmp1630;
  wire tmp1631;
  wire tmp1632;
  wire tmp1633;
  wire tmp1634;
  wire tmp1635;
  wire tmp1636;
  wire tmp1637;
  wire tmp1638;
  wire tmp1639;
  wire tmp1640;
  wire tmp1641;
  wire tmp1642;
  wire tmp1643;
  wire tmp1644;
  wire tmp1645;
  wire tmp1646;
  wire tmp1647;
  wire tmp1648;
  wire tmp1649;
  wire tmp1650;
  wire tmp1651;
  wire tmp1652;
  wire tmp1653;
  wire tmp1654;
  wire tmp1655;
  wire tmp1656;
  wire tmp1657;
  wire tmp1658;
  wire tmp1659;
  wire tmp1660;
  wire tmp1661;
  wire tmp1662;
  wire tmp1663;
  wire tmp1664;
  wire tmp1665;
  wire tmp1666;
  wire tmp1667;
  wire tmp1668;
  wire tmp1669;
  wire tmp1670;
  wire tmp1671;
  wire tmp1672;
  wire tmp1673;
  wire tmp1674;
  wire tmp1675;
  wire tmp1676;
  wire tmp1677;
  wire tmp1678;
  wire tmp1679;
  wire tmp1680;
  wire tmp1681;
  wire tmp1682;
  wire tmp1683;
  wire tmp1684;
  wire tmp1685;
  wire tmp1686;
  wire tmp1687;
  wire tmp1688;
  wire tmp1689;
  wire tmp1690;
  wire tmp1691;
  wire tmp1692;
  wire tmp1693;
  wire tmp1694;
  wire tmp1695;
  wire tmp1696;
  wire tmp1697;
  wire tmp1698;
  wire tmp1699;
  wire tmp1700;
  wire tmp1701;
  wire tmp1702;
  wire tmp1703;
  wire tmp1704;
  wire tmp1705;
  wire tmp1706;
  wire tmp1707;
  wire tmp1708;
  wire tmp1709;
  wire tmp1710;
  wire tmp1711;
  wire tmp1712;
  wire tmp1713;
  wire tmp1714;
  wire tmp1715;
  wire tmp1716;
  wire tmp1717;
  wire tmp1718;
  wire tmp1719;
  wire tmp1720;
  wire tmp1721;
  wire tmp1722;
  wire tmp1723;
  wire tmp1724;
  wire tmp1725;
  wire tmp1726;
  wire tmp1727;
  wire tmp1728;
  wire tmp1729;
  wire tmp1730;
  wire tmp1731;
  wire tmp1732;
  wire tmp1733;
  wire tmp1734;
  wire tmp1735;
  wire tmp1736;
  wire tmp1737;
  wire tmp1738;
  wire tmp1739;
  wire tmp1740;
  wire tmp1741;
  wire tmp1742;
  wire tmp1743;
  wire tmp1744;
  wire tmp1745;
  wire tmp1746;
  wire tmp1747;
  wire tmp1748;
  wire tmp1749;
  wire tmp1750;
  wire tmp1751;
  wire tmp1752;
  wire tmp1753;
  wire tmp1754;
  wire tmp1755;
  wire tmp1756;
  wire tmp1757;
  wire tmp1758;
  wire tmp1759;
  wire tmp1760;
  wire tmp1761;
  wire tmp1762;
  wire tmp1763;
  wire tmp1764;
  wire tmp1765;
  wire tmp1766;
  wire tmp1767;
  wire tmp1768;
  wire tmp1769;
  wire tmp1770;
  wire tmp1771;
  wire tmp1772;
  wire tmp1773;
  wire tmp1774;
  wire tmp1775;
  wire tmp1776;
  wire tmp1777;
  wire tmp1778;
  wire tmp1779;
  wire tmp1780;
  wire tmp1781;
  wire tmp1782;
  wire tmp1783;
  wire tmp1784;
  wire tmp1785;
  wire tmp1786;
  wire tmp1787;
  wire tmp1788;
  wire tmp1789;
  wire tmp1790;
  wire tmp1791;
  wire tmp1792;
  wire tmp1793;
  wire tmp1794;
  wire tmp1795;
  wire tmp1796;
  wire tmp1797;
  wire tmp1798;
  wire tmp1799;
  wire tmp1800;
  wire tmp1801;
  wire tmp1802;
  wire tmp1803;
  wire tmp1804;
  wire tmp1805;
  wire tmp1806;
  wire tmp1807;
  wire tmp1808;
  wire tmp1809;
  wire tmp1810;
  wire tmp1811;
  wire tmp1812;
  wire tmp1813;
  wire tmp1814;
  wire tmp1815;
  wire tmp1816;
  wire tmp1817;
  wire tmp1818;
  wire tmp1819;
  wire tmp1820;
  wire tmp1821;
  wire tmp1822;
  wire tmp1823;
  wire tmp1824;
  wire tmp1825;
  wire tmp1826;
  wire tmp1827;
  wire tmp1828;
  wire tmp1829;
  wire tmp1830;
  wire tmp1831;
  wire tmp1832;
  wire tmp1833;
  wire tmp1834;
  wire tmp1835;
  wire tmp1836;
  wire tmp1837;
  wire tmp1838;
  wire tmp1839;
  wire tmp1840;
  wire tmp1841;
  wire tmp1842;
  wire tmp1843;
  wire tmp1844;
  wire tmp1845;
  wire tmp1846;
  wire tmp1847;
  wire tmp1848;
  wire tmp1849;
  wire tmp1850;
  wire tmp1851;
  wire tmp1852;
  wire tmp1853;
  wire tmp1854;
  wire tmp1855;
  wire tmp1856;
  wire tmp1857;
  wire tmp1858;
  wire tmp1859;
  wire tmp1860;
  wire tmp1861;
  wire tmp1862;
  wire tmp1863;
  wire tmp1864;
  wire tmp1865;
  wire tmp1866;
  wire tmp1867;
  wire tmp1868;
  wire tmp1869;
  wire tmp1870;
  wire tmp1871;
  wire tmp1872;
  wire tmp1873;
  wire tmp1874;
  wire tmp1875;
  wire tmp1876;
  wire tmp1877;
  wire tmp1878;
  wire tmp1879;
  wire tmp1880;
  wire tmp1881;
  wire tmp1882;
  wire tmp1883;
  wire tmp1884;
  wire tmp1885;
  wire tmp1886;
  wire tmp1887;
  wire tmp1888;
  wire tmp1889;
  wire tmp1890;
  wire tmp1891;
  wire tmp1892;
  wire tmp1893;
  wire tmp1894;
  wire tmp1895;
  wire tmp1896;
  wire tmp1897;
  wire tmp1898;
  wire tmp1899;
  wire tmp1900;
  wire tmp1901;
  wire tmp1902;
  wire tmp1903;
  wire tmp1904;
  wire tmp1905;
  wire tmp1906;
  wire tmp1907;
  wire tmp1908;
  wire tmp1909;
  wire tmp1910;
  wire tmp1911;
  wire tmp1912;
  wire tmp1913;
  wire tmp1914;
  wire tmp1915;
  wire tmp1916;
  wire tmp1917;
  wire tmp1918;
  wire tmp1919;
  wire tmp1920;
  wire tmp1921;
  wire tmp1922;
  wire tmp1923;
  wire tmp1924;
  wire tmp1925;
  wire tmp1926;
  wire tmp1927;
  wire tmp1928;
  wire tmp1929;
  wire tmp1930;
  wire tmp1931;
  wire tmp1932;
  wire tmp1933;
  wire tmp1934;
  wire tmp1935;
  wire tmp1936;
  wire tmp1937;
  wire tmp1938;
  wire tmp1939;
  wire tmp1940;
  wire tmp1941;
  wire tmp1942;
  wire tmp1943;
  wire tmp1944;
  wire tmp1945;
  wire tmp1946;
  wire tmp1947;
  wire tmp1948;
  wire tmp1949;
  wire tmp1950;
  wire tmp1951;
  wire tmp1952;
  wire tmp1953;
  wire tmp1954;
  wire tmp1955;
  wire tmp1956;
  wire tmp1957;
  wire tmp1958;
  wire tmp1959;
  wire tmp1960;
  wire tmp1961;
  wire tmp1962;
  wire tmp1963;
  wire tmp1964;
  wire tmp1965;
  wire tmp1966;
  wire tmp1967;
  wire tmp1968;
  wire tmp1969;
  wire tmp1970;
  wire tmp1971;
  wire tmp1972;
  wire tmp1973;
  wire tmp1974;
  wire tmp1975;
  wire tmp1976;
  wire tmp1977;
  wire tmp1978;
  wire tmp1979;
  wire tmp1980;
  wire tmp1981;
  wire tmp1982;
  wire tmp1983;
  wire tmp1984;
  wire tmp1985;
  wire tmp1986;
  wire tmp1987;
  wire tmp1988;
  wire tmp1989;
  wire tmp1990;
  wire tmp1991;
  wire tmp1992;
  wire tmp1993;
  wire tmp1994;
  wire tmp1995;
  wire tmp1996;
  wire tmp1997;
  wire tmp1998;
  wire tmp1999;
  wire tmp2000;
  wire tmp2001;
  wire tmp2002;
  wire tmp2003;
  wire tmp2004;
  wire tmp2005;
  wire tmp2006;
  wire tmp2007;
  wire tmp2008;
  wire tmp2009;
  wire tmp2010;
  wire tmp2011;
  wire tmp2012;
  wire tmp2013;
  wire tmp2014;
  wire tmp2015;
  wire tmp2016;
  wire tmp2017;
  wire tmp2018;
  wire tmp2019;
  wire tmp2020;
  wire tmp2021;
  wire tmp2022;
  wire tmp2023;
  wire tmp2024;
  wire tmp2025;
  wire tmp2026;
  wire tmp2027;
  wire tmp2028;
  wire tmp2029;
  wire tmp2030;
  wire tmp2031;
  wire tmp2032;
  wire tmp2033;
  wire tmp2034;
  wire tmp2035;
  wire tmp2036;
  wire tmp2037;
  wire tmp2038;
  wire tmp2039;
  wire tmp2040;
  wire tmp2041;
  wire tmp2042;
  wire tmp2043;
  wire tmp2044;
  wire tmp2045;
  wire tmp2046;
  wire tmp2047;
  wire tmp2048;
  wire tmp2049;
  wire tmp2050;
  wire tmp2051;
  wire tmp2052;
  wire tmp2053;
  wire tmp2054;
  wire tmp2055;
  wire tmp2056;
  wire tmp2057;
  wire tmp2058;
  wire tmp2059;
  wire tmp2060;
  wire tmp2061;
  wire tmp2062;
  wire tmp2063;
  wire tmp2064;
  wire tmp2065;
  wire tmp2066;
  wire tmp2067;
  wire tmp2068;
  wire tmp2069;
  wire tmp2070;
  wire tmp2071;
  wire tmp2072;
  wire tmp2073;
  wire tmp2074;
  wire tmp2075;
  wire tmp2076;
  wire tmp2077;
  wire tmp2078;
  wire tmp2079;
  wire tmp2080;
  wire tmp2081;
  wire tmp2082;
  wire tmp2083;
  wire tmp2084;
  wire tmp2085;
  wire tmp2086;
  wire tmp2087;
  wire tmp2088;
  wire tmp2089;
  wire tmp2090;
  wire tmp2091;
  wire tmp2092;
  wire tmp2093;
  wire tmp2094;
  wire tmp2095;
  wire tmp2096;
  wire tmp2097;
  wire tmp2098;
  wire tmp2099;
  wire tmp2100;
  wire tmp2101;
  wire tmp2102;
  wire tmp2103;
  wire tmp2104;
  wire tmp2105;
  wire tmp2106;
  wire tmp2107;
  wire tmp2108;
  wire tmp2109;
  wire tmp2110;
  wire tmp2111;
  wire tmp2112;
  wire tmp2113;
  wire tmp2114;
  wire tmp2115;
  wire tmp2116;
  wire tmp2117;
  wire tmp2118;
  wire tmp2119;
  wire tmp2120;
  wire tmp2121;
  wire tmp2122;
  wire tmp2123;
  wire tmp2124;
  wire tmp2125;
  wire tmp2126;
  wire tmp2127;
  wire tmp2128;
  wire tmp2129;
  wire tmp2130;
  wire tmp2131;
  wire tmp2132;
  wire tmp2133;
  wire tmp2134;
  wire tmp2135;
  wire tmp2136;
  wire tmp2137;
  wire tmp2138;
  wire tmp2139;
  wire tmp2140;
  wire tmp2141;
  wire tmp2142;
  wire tmp2143;
  wire tmp2144;
  wire tmp2145;
  wire tmp2146;
  wire tmp2147;
  wire tmp2148;
  wire tmp2149;
  wire tmp2150;
  wire tmp2151;
  wire tmp2152;
  wire tmp2153;
  wire tmp2154;
  wire tmp2155;
  wire tmp2156;
  wire tmp2157;
  wire tmp2158;
  wire tmp2159;
  wire tmp2160;
  wire tmp2161;
  wire tmp2162;
  wire tmp2163;
  wire tmp2164;
  wire tmp2165;
  wire tmp2166;
  wire tmp2167;
  wire tmp2168;
  wire tmp2169;
  wire tmp2170;
  wire tmp2171;
  wire tmp2172;
  wire tmp2173;
  wire tmp2174;
  wire tmp2175;
  wire tmp2176;
  wire tmp2177;
  wire tmp2178;
  wire tmp2179;
  wire tmp2180;
  wire tmp2181;
  wire tmp2182;
  wire tmp2183;
  wire tmp2184;
  wire tmp2185;
  wire tmp2186;
  wire tmp2187;
  wire tmp2188;
  wire tmp2189;
  wire tmp2190;
  wire tmp2191;
  wire tmp2192;
  wire tmp2193;
  wire tmp2194;
  wire tmp2195;
  wire tmp2196;
  wire tmp2197;
  wire tmp2198;
  wire tmp2199;
  wire tmp2200;
  wire tmp2201;
  wire tmp2202;
  wire tmp2203;
  wire tmp2204;
  wire tmp2205;
  wire tmp2206;
  wire tmp2207;
  wire tmp2208;
  wire tmp2209;
  wire tmp2210;
  wire tmp2211;
  wire tmp2212;
  wire tmp2213;
  wire tmp2214;
  wire tmp2215;
  wire tmp2216;
  wire tmp2217;
  wire tmp2218;
  wire tmp2219;
  wire tmp2220;
  wire tmp2221;
  wire tmp2222;
  wire tmp2223;
  wire tmp2224;
  wire tmp2225;
  wire tmp2226;
  wire tmp2227;
  wire tmp2228;
  wire tmp2229;
  wire tmp2230;
  wire tmp2231;
  wire tmp2232;
  wire tmp2233;
  wire tmp2234;
  wire tmp2235;
  wire tmp2236;
  wire tmp2237;
  wire tmp2238;
  wire tmp2239;
  wire tmp2240;
  wire tmp2241;
  wire tmp2242;
  wire tmp2243;
  wire tmp2244;
  wire tmp2245;
  wire tmp2246;
  wire tmp2247;
  wire tmp2248;
  wire tmp2249;
  wire tmp2250;
  wire tmp2251;
  wire tmp2252;
  wire tmp2253;
  wire tmp2254;
  wire tmp2255;
  wire tmp2256;
  wire tmp2257;
  wire tmp2258;
  wire tmp2259;
  wire tmp2260;
  wire tmp2261;
  wire tmp2262;
  wire tmp2263;
  wire tmp2264;
  wire tmp2265;
  wire tmp2266;
  wire tmp2267;
  wire tmp2268;
  wire tmp2269;
  wire tmp2270;
  wire tmp2271;
  wire tmp2272;
  wire tmp2273;
  wire tmp2274;
  wire tmp2275;
  wire tmp2276;
  wire tmp2277;
  wire tmp2278;
  wire tmp2279;
  wire tmp2280;
  wire tmp2281;
  wire tmp2282;
  wire tmp2283;
  wire tmp2284;
  wire tmp2285;
  wire tmp2286;
  wire tmp2287;
  wire tmp2288;
  wire tmp2289;
  wire tmp2290;
  wire tmp2291;
  wire tmp2292;
  wire tmp2293;
  wire tmp2294;
  wire tmp2295;
  wire tmp2296;
  wire tmp2297;
  wire tmp2298;
  wire tmp2299;
  wire tmp2300;
  wire tmp2301;
  wire tmp2302;
  wire tmp2303;
  wire tmp2304;
  wire tmp2305;
  wire tmp2306;
  wire tmp2307;
  wire tmp2308;
  wire tmp2309;
  wire tmp2310;
  wire tmp2311;
  wire tmp2312;
  wire tmp2313;
  wire tmp2314;
  wire tmp2315;
  wire tmp2316;
  wire tmp2317;
  wire tmp2318;
  wire tmp2319;
  wire tmp2320;
  wire tmp2321;
  wire tmp2322;
  wire tmp2323;
  wire tmp2324;
  wire tmp2325;
  wire tmp2326;
  wire tmp2327;
  wire tmp2328;
  wire tmp2329;
  wire tmp2330;
  wire tmp2331;
  wire tmp2332;
  wire tmp2333;
  wire tmp2334;
  wire tmp2335;
  wire tmp2336;
  wire tmp2337;
  wire tmp2338;
  wire tmp2339;
  wire tmp2340;
  wire tmp2341;
  wire tmp2342;
  wire tmp2343;
  wire tmp2344;
  wire tmp2345;
  wire tmp2346;
  wire tmp2347;
  wire tmp2348;
  wire tmp2349;
  wire tmp2350;
  wire tmp2351;
  wire tmp2352;
  wire tmp2353;
  wire tmp2354;
  wire tmp2355;
  wire tmp2356;
  wire tmp2357;
  wire tmp2358;
  wire tmp2359;
  wire tmp2360;
  wire tmp2361;
  wire tmp2362;
  wire tmp2363;
  wire tmp2364;
  wire tmp2365;
  wire tmp2366;
  wire tmp2367;
  wire tmp2368;
  wire tmp2369;
  wire tmp2370;
  wire tmp2371;
  wire tmp2372;
  wire tmp2373;
  wire tmp2374;
  wire tmp2375;
  wire tmp2376;
  wire tmp2377;
  wire tmp2378;
  wire tmp2379;
  wire tmp2380;
  wire tmp2381;
  wire tmp2382;
  wire tmp2383;
  wire tmp2384;
  wire tmp2385;
  wire tmp2386;
  wire tmp2387;
  wire tmp2388;
  wire tmp2389;
  wire tmp2390;
  wire tmp2391;
  wire tmp2392;
  wire tmp2393;
  wire tmp2394;
  wire tmp2395;
  wire tmp2396;
  wire tmp2397;
  wire tmp2398;
  wire tmp2399;
  wire tmp2400;
  wire tmp2401;
  wire tmp2402;
  wire tmp2403;
  wire tmp2404;
  wire tmp2405;
  wire tmp2406;
  wire tmp2407;
  wire tmp2408;
  wire tmp2409;
  wire tmp2410;
  wire tmp2411;
  wire tmp2412;
  wire tmp2413;
  wire tmp2414;
  wire tmp2415;
  wire tmp2416;
  wire tmp2417;
  wire tmp2418;
  wire tmp2419;
  wire tmp2420;
  wire tmp2421;
  wire tmp2422;
  wire tmp2423;
  wire tmp2424;
  wire tmp2425;
  wire tmp2426;
  wire tmp2427;
  wire tmp2428;
  wire tmp2429;
  wire tmp2430;
  wire tmp2431;
  wire tmp2432;
  wire tmp2433;
  wire tmp2434;
  wire tmp2435;
  wire tmp2436;
  wire tmp2437;
  wire tmp2438;
  wire tmp2439;
  wire tmp2440;
  wire tmp2441;
  wire tmp2442;
  wire tmp2443;
  wire tmp2444;
  wire tmp2445;
  wire tmp2446;
  wire tmp2447;
  wire tmp2448;
  wire tmp2449;
  wire tmp2450;
  wire tmp2451;
  wire tmp2452;
  wire tmp2453;
  wire tmp2454;
  wire tmp2455;
  wire tmp2456;
  wire tmp2457;
  wire tmp2458;
  wire tmp2459;
  wire tmp2460;
  wire tmp2461;
  wire tmp2462;
  wire tmp2463;
  wire tmp2464;
  wire tmp2465;
  wire tmp2466;
  wire tmp2467;
  wire tmp2468;
  wire tmp2469;
  wire tmp2470;
  wire tmp2471;
  wire tmp2472;
  wire tmp2473;
  wire tmp2474;
  wire tmp2475;
  wire tmp2476;
  wire tmp2477;
  wire tmp2478;
  wire tmp2479;
  wire tmp2480;
  wire tmp2481;
  wire tmp2482;
  wire tmp2483;
  wire tmp2484;
  wire tmp2485;
  wire tmp2486;
  wire tmp2487;
  wire tmp2488;
  wire tmp2489;
  wire tmp2490;
  wire tmp2491;
  wire tmp2492;
  wire tmp2493;
  wire tmp2494;
  wire tmp2495;
  wire tmp2496;
  wire tmp2497;
  wire tmp2498;
  wire tmp2499;
  wire tmp2500;
  wire tmp2501;
  wire tmp2502;
  wire tmp2503;
  wire tmp2504;
  wire tmp2505;
  wire tmp2506;
  wire tmp2507;
  wire tmp2508;
  wire tmp2509;
  wire tmp2510;
  wire tmp2511;
  wire tmp2512;
  wire tmp2513;
  wire tmp2514;
  wire tmp2515;
  wire tmp2516;
  wire tmp2517;
  wire tmp2518;
  wire tmp2519;
  wire tmp2520;
  wire tmp2521;
  wire tmp2522;
  wire tmp2523;
  wire tmp2524;
  wire tmp2525;
  wire tmp2526;
  wire tmp2527;
  wire tmp2528;
  wire tmp2529;
  wire tmp2530;
  wire tmp2531;
  wire tmp2532;
  wire tmp2533;
  wire tmp2534;
  wire tmp2535;
  wire tmp2536;
  wire tmp2537;
  wire tmp2538;
  wire tmp2539;
  wire tmp2540;
  wire tmp2541;
  wire tmp2542;
  wire tmp2543;
  wire tmp2544;
  wire tmp2545;
  wire tmp2546;
  wire tmp2547;
  wire tmp2548;
  wire tmp2549;
  wire tmp2550;
  wire tmp2551;
  wire tmp2552;
  wire tmp2553;
  wire tmp2554;
  wire tmp2555;
  wire tmp2556;
  wire tmp2557;
  wire tmp2558;
  wire tmp2559;
  wire tmp2560;
  wire tmp2561;
  wire tmp2562;
  wire tmp2563;
  wire tmp2564;
  wire tmp2565;
  wire tmp2566;
  wire tmp2567;
  wire tmp2568;
  wire tmp2569;
  wire tmp2570;
  wire tmp2571;
  wire tmp2572;
  wire tmp2573;
  wire tmp2574;
  wire tmp2575;
  wire tmp2576;
  wire tmp2577;
  wire tmp2578;
  wire tmp2579;
  wire tmp2580;
  wire tmp2581;
  wire tmp2582;
  wire tmp2583;
  wire tmp2584;
  wire tmp2585;
  wire tmp2586;
  wire tmp2587;
  wire tmp2588;
  wire tmp2589;
  wire tmp2590;
  wire tmp2591;
  wire tmp2592;
  wire tmp2593;
  wire tmp2594;
  wire tmp2595;
  wire tmp2596;
  wire tmp2597;
  wire tmp2598;
  wire tmp2599;
  wire tmp2600;
  wire tmp2601;
  wire tmp2602;
  wire tmp2603;
  wire tmp2604;
  wire tmp2605;
  wire tmp2606;
  wire tmp2607;
  wire tmp2608;
  wire tmp2609;
  wire tmp2610;
  wire tmp2611;
  wire tmp2612;
  wire tmp2613;
  wire tmp2614;
  wire tmp2615;
  wire tmp2616;
  wire tmp2617;
  wire tmp2618;
  wire tmp2619;
  wire tmp2620;
  wire tmp2621;
  wire tmp2622;
  wire tmp2623;
  wire tmp2624;
  wire tmp2625;
  wire tmp2626;
  wire tmp2627;
  wire tmp2628;
  wire tmp2629;
  wire tmp2630;
  wire tmp2631;
  wire tmp2632;
  wire tmp2633;
  wire tmp2634;
  wire tmp2635;
  wire tmp2636;
  wire tmp2637;
  wire tmp2638;
  wire tmp2639;
  wire tmp2640;
  wire tmp2641;
  wire tmp2642;
  wire tmp2643;
  wire tmp2644;
  wire tmp2645;
  wire tmp2646;
  wire tmp2647;
  wire tmp2648;
  wire tmp2649;
  wire tmp2650;
  wire tmp2651;
  wire tmp2652;
  wire tmp2653;
  wire tmp2654;
  wire tmp2655;
  wire tmp2656;
  wire tmp2657;
  wire tmp2658;
  wire tmp2659;
  wire tmp2660;
  wire tmp2661;
  wire tmp2662;
  wire tmp2663;
  wire tmp2664;
  wire tmp2665;
  wire tmp2666;
  wire tmp2667;
  wire tmp2668;
  wire tmp2669;
  wire tmp2670;
  wire tmp2671;
  wire tmp2672;
  wire tmp2673;
  wire tmp2674;
  wire tmp2675;
  wire tmp2676;
  wire tmp2677;
  wire tmp2678;
  wire tmp2679;
  wire tmp2680;
  wire tmp2681;
  wire tmp2682;
  wire tmp2683;
  wire tmp2684;
  wire tmp2685;
  wire tmp2686;
  wire tmp2687;
  wire tmp2688;
  wire tmp2689;
  wire tmp2690;
  wire tmp2691;
  wire tmp2692;
  wire tmp2693;
  wire tmp2694;
  wire tmp2695;
  wire tmp2696;
  wire tmp2697;
  wire tmp2698;
  wire tmp2699;
  wire tmp2700;
  wire tmp2701;
  wire tmp2702;
  wire tmp2703;
  wire tmp2704;
  wire tmp2705;
  wire tmp2706;
  wire tmp2707;
  wire tmp2708;
  wire tmp2709;
  wire tmp2710;
  wire tmp2711;
  wire tmp2712;
  wire tmp2713;
  wire tmp2714;
  wire tmp2715;
  wire tmp2716;
  wire tmp2717;
  wire tmp2718;
  wire tmp2719;
  wire tmp2720;
  wire tmp2721;
  wire tmp2722;
  wire tmp2723;
  wire tmp2724;
  wire tmp2725;
  wire tmp2726;
  wire tmp2727;
  wire tmp2728;
  wire tmp2729;
  wire tmp2730;
  wire tmp2731;
  wire tmp2732;
  wire tmp2733;
  wire tmp2734;
  wire tmp2735;
  wire tmp2736;
  wire tmp2737;
  wire tmp2738;
  wire tmp2739;
  wire tmp2740;
  wire tmp2741;
  wire tmp2742;
  wire tmp2743;
  wire tmp2744;
  wire tmp2745;
  wire tmp2746;
  wire tmp2747;
  wire tmp2748;
  wire tmp2749;
  wire tmp2750;
  wire tmp2751;
  wire tmp2752;
  wire tmp2753;
  wire tmp2754;
  wire tmp2755;
  wire tmp2756;
  wire tmp2757;
  wire tmp2758;
  wire tmp2759;
  wire tmp2760;
  wire tmp2761;
  wire tmp2762;
  wire tmp2763;
  wire tmp2764;
  wire tmp2765;
  wire tmp2766;
  wire tmp2767;
  wire tmp2768;
  wire tmp2769;
  wire tmp2770;
  wire tmp2771;
  wire tmp2772;
  wire tmp2773;
  wire tmp2774;
  wire tmp2775;
  wire tmp2776;
  wire tmp2777;
  wire tmp2778;
  wire tmp2779;
  wire tmp2780;
  wire tmp2781;
  wire tmp2782;
  wire tmp2783;
  wire tmp2784;
  wire tmp2785;
  wire tmp2786;
  wire tmp2787;
  wire tmp2788;
  wire tmp2789;
  wire tmp2790;
  wire tmp2791;
  wire tmp2792;
  wire tmp2793;
  wire tmp2794;
  wire tmp2795;
  wire tmp2796;
  wire tmp2797;
  wire tmp2798;
  wire tmp2799;
  wire tmp2800;
  wire tmp2801;
  wire tmp2802;
  wire tmp2803;
  wire tmp2804;
  wire tmp2805;
  wire tmp2806;
  wire tmp2807;
  wire tmp2808;
  wire tmp2809;
  wire tmp2810;
  wire tmp2811;
  wire tmp2812;
  wire tmp2813;
  wire tmp2814;
  wire tmp2815;
  wire tmp2816;
  wire tmp2817;
  wire tmp2818;
  wire tmp2819;
  wire tmp2820;
  wire tmp2821;
  wire tmp2822;
  wire tmp2823;
  wire tmp2824;
  wire tmp2825;
  wire tmp2826;
  wire tmp2827;
  wire tmp2828;
  wire tmp2829;
  wire tmp2830;
  wire tmp2831;
  wire tmp2832;
  wire tmp2833;
  wire tmp2834;
  wire tmp2835;
  wire tmp2836;
  wire tmp2837;
  wire tmp2838;
  wire tmp2839;
  wire tmp2840;
  wire tmp2841;
  wire tmp2842;
  wire tmp2843;
  wire tmp2844;
  wire tmp2845;
  wire tmp2846;
  wire tmp2847;
  wire tmp2848;
  wire tmp2849;
  wire tmp2850;
  wire tmp2851;
  wire tmp2852;
  wire tmp2853;
  wire tmp2854;
  wire tmp2855;
  wire tmp2856;
  wire tmp2857;
  wire tmp2858;
  wire tmp2859;
  wire tmp2860;
  wire tmp2861;
  wire tmp2862;
  wire tmp2863;
  wire tmp2864;
  wire tmp2865;
  wire tmp2866;
  wire tmp2867;
  wire tmp2868;
  wire tmp2869;
  wire tmp2870;
  wire tmp2871;
  wire tmp2872;
  wire tmp2873;
  wire tmp2874;
  wire tmp2875;
  wire tmp2876;
  wire tmp2877;
  wire tmp2878;
  wire tmp2879;
  wire tmp2880;
  wire tmp2881;
  wire tmp2882;
  wire tmp2883;
  wire tmp2884;
  wire tmp2885;
  wire tmp2886;
  wire tmp2887;
  wire tmp2888;
  wire tmp2889;
  wire tmp2890;
  wire tmp2891;
  wire tmp2892;
  wire tmp2893;
  wire tmp2894;
  wire tmp2895;
  wire tmp2896;
  wire tmp2897;
  wire tmp2898;
  wire tmp2899;
  wire tmp2900;
  wire tmp2901;
  wire tmp2902;
  wire tmp2903;
  wire tmp2904;
  wire tmp2905;
  wire tmp2906;
  wire tmp2907;
  wire tmp2908;
  wire tmp2909;
  wire tmp2910;
  wire tmp2911;
  wire tmp2912;
  wire tmp2913;
  wire tmp2914;
  wire tmp2915;
  wire tmp2916;
  wire tmp2917;
  wire tmp2918;
  wire tmp2919;
  wire tmp2920;
  wire tmp2921;
  wire tmp2922;
  wire tmp2923;
  wire tmp2924;
  wire tmp2925;
  wire tmp2926;
  wire tmp2927;
  wire tmp2928;
  wire tmp2929;
  wire tmp2930;
  wire tmp2931;
  wire tmp2932;
  wire tmp2933;
  wire tmp2934;
  wire tmp2935;
  wire tmp2936;
  wire tmp2937;
  wire tmp2938;
  wire tmp2939;
  wire tmp2940;
  wire tmp2941;
  wire tmp2942;
  wire tmp2943;
  wire tmp2944;
  wire tmp2945;
  wire tmp2946;
  wire tmp2947;
  wire tmp2948;
  wire tmp2949;
  wire tmp2950;
  wire tmp2951;
  wire tmp2952;
  wire tmp2953;
  wire tmp2954;
  wire tmp2955;
  wire tmp2956;
  wire tmp2957;
  wire tmp2958;
  wire tmp2959;
  wire tmp2960;
  wire tmp2961;
  wire tmp2962;
  wire tmp2963;
  wire tmp2964;
  wire tmp2965;
  wire tmp2966;
  wire tmp2967;
  wire tmp2968;
  wire tmp2969;
  wire tmp2970;
  wire tmp2971;
  wire tmp2972;
  wire tmp2973;
  wire tmp2974;
  wire tmp2975;
  wire tmp2976;
  wire tmp2977;
  wire tmp2978;
  wire tmp2979;
  wire tmp2980;
  wire tmp2981;
  wire tmp2982;
  wire tmp2983;
  wire tmp2984;
  wire tmp2985;
  wire tmp2986;
  wire tmp2987;
  wire tmp2988;
  wire tmp2989;
  wire tmp2990;
  wire tmp2991;
  wire tmp2992;
  wire tmp2993;
  wire tmp2994;
  wire tmp2995;
  wire tmp2996;
  wire tmp2997;
  wire tmp2998;
  wire tmp2999;
  wire tmp3000;
  wire tmp3001;
  wire tmp3002;
  wire tmp3003;
  wire tmp3004;
  wire tmp3005;
  wire tmp3006;
  wire tmp3007;
  wire tmp3008;
  wire tmp3009;
  wire tmp3010;
  wire tmp3011;
  wire tmp3012;
  wire tmp3013;
  wire tmp3014;
  wire tmp3015;
  wire tmp3016;
  wire tmp3017;
  wire tmp3018;
  wire tmp3019;
  wire tmp3020;
  wire tmp3021;
  wire tmp3022;
  wire tmp3023;
  wire tmp3024;
  wire tmp3025;
  wire tmp3026;
  wire tmp3027;
  wire tmp3028;
  wire tmp3029;
  wire tmp3030;
  wire tmp3031;
  wire tmp3032;
  wire tmp3033;
  wire tmp3034;
  wire tmp3035;
  wire tmp3036;
  wire tmp3037;
  wire tmp3038;
  wire tmp3039;
  wire tmp3040;
  wire tmp3041;
  wire tmp3042;
  wire tmp3043;
  wire tmp3044;
  wire tmp3045;
  wire tmp3046;
  wire tmp3047;
  wire tmp3048;
  wire tmp3049;
  wire tmp3050;
  wire tmp3051;
  wire tmp3052;
  wire tmp3053;
  wire tmp3054;
  wire tmp3055;
  wire tmp3056;
  wire tmp3057;
  wire tmp3058;
  wire tmp3059;
  wire tmp3060;
  wire tmp3061;
  wire tmp3062;
  wire tmp3063;
  wire tmp3064;
  wire tmp3065;
  wire tmp3066;
  wire tmp3067;
  wire tmp3068;
  wire tmp3069;
  wire tmp3070;
  wire tmp3071;
  wire tmp3072;
  wire tmp3073;
  wire tmp3074;
  wire tmp3075;
  wire tmp3076;
  wire tmp3077;
  wire tmp3078;
  wire tmp3079;
  wire tmp3080;
  wire tmp3081;
  wire tmp3082;
  wire tmp3083;
  wire tmp3084;
  wire tmp3085;
  wire tmp3086;
  wire tmp3087;
  wire tmp3088;
  wire tmp3089;
  wire tmp3090;
  wire tmp3091;
  wire tmp3092;
  wire tmp3093;
  wire tmp3094;
  wire tmp3095;
  wire tmp3096;
  wire tmp3097;
  wire tmp3098;
  wire tmp3099;
  wire tmp3100;
  wire tmp3101;
  wire tmp3102;
  wire tmp3103;
  wire tmp3104;
  wire tmp3105;
  wire tmp3106;
  wire tmp3107;
  wire tmp3108;
  wire tmp3109;
  wire tmp3110;
  wire tmp3111;
  wire tmp3112;
  wire tmp3113;
  wire tmp3114;
  wire tmp3115;
  wire tmp3116;
  wire tmp3117;
  wire tmp3118;
  wire tmp3119;
  wire tmp3120;
  wire tmp3121;
  wire tmp3122;
  wire tmp3123;
  wire tmp3124;
  wire tmp3125;
  wire tmp3126;
  wire tmp3127;
  wire tmp3128;
  wire tmp3129;
  wire tmp3130;
  wire tmp3131;
  wire tmp3132;
  wire tmp3133;
  wire tmp3134;
  wire tmp3135;
  wire tmp3136;
  wire tmp3137;
  wire tmp3138;
  wire tmp3139;
  wire tmp3140;
  wire tmp3141;
  wire tmp3142;
  wire tmp3143;
  wire tmp3144;
  wire tmp3145;
  wire tmp3146;
  wire tmp3147;
  wire tmp3148;
  wire tmp3149;
  wire tmp3150;
  wire tmp3151;
  wire tmp3152;
  wire tmp3153;
  wire tmp3154;
  wire tmp3155;
  wire tmp3156;
  wire tmp3157;
  wire tmp3158;
  wire tmp3159;
  wire tmp3160;
  wire tmp3161;
  wire tmp3162;
  wire tmp3163;
  wire tmp3164;
  wire tmp3165;
  wire tmp3166;
  wire tmp3167;
  wire tmp3168;
  wire tmp3169;
  wire tmp3170;
  wire tmp3171;
  wire tmp3172;
  wire tmp3173;
  wire tmp3174;
  wire tmp3175;
  wire tmp3176;
  wire tmp3177;
  wire tmp3178;
  wire tmp3179;
  wire tmp3180;
  wire tmp3181;
  wire tmp3182;
  wire tmp3183;
  wire tmp3184;
  wire tmp3185;
  wire tmp3186;
  wire tmp3187;
  wire tmp3188;
  wire tmp3189;
  wire tmp3190;
  wire tmp3191;
  wire tmp3192;
  wire tmp3193;
  wire tmp3194;
  wire tmp3195;
  wire tmp3196;
  wire tmp3197;
  wire tmp3198;
  wire tmp3199;
  wire tmp3200;
  wire tmp3201;
  wire tmp3202;
  wire tmp3203;
  wire tmp3204;
  wire tmp3205;
  wire tmp3206;
  wire tmp3207;
  wire tmp3208;
  wire tmp3209;
  wire tmp3210;
  wire tmp3211;
  wire tmp3212;
  wire tmp3213;
  wire tmp3214;
  wire tmp3215;
  wire tmp3216;
  wire tmp3217;
  wire tmp3218;
  wire tmp3219;
  wire tmp3220;
  wire tmp3221;
  wire tmp3222;
  wire tmp3223;
  wire tmp3224;
  wire tmp3225;
  wire tmp3226;
  wire tmp3227;
  wire tmp3228;
  wire tmp3229;
  wire tmp3230;
  wire tmp3231;
  wire tmp3232;
  wire tmp3233;
  wire tmp3234;
  wire tmp3235;
  wire tmp3236;
  wire tmp3237;
  wire tmp3238;
  wire tmp3239;
  wire tmp3240;
  wire tmp3241;
  wire tmp3242;
  wire tmp3243;
  wire tmp3244;
  wire tmp3245;
  wire tmp3246;
  wire tmp3247;
  wire tmp3248;
  wire tmp3249;
  wire tmp3250;
  wire tmp3251;
  wire tmp3252;
  wire tmp3253;
  wire tmp3254;
  wire tmp3255;
  wire tmp3256;
  wire tmp3257;
  wire tmp3258;
  wire tmp3259;
  wire tmp3260;
  wire tmp3261;
  wire tmp3262;
  wire tmp3263;
  wire tmp3264;
  wire tmp3265;
  wire tmp3266;
  wire tmp3267;
  wire tmp3268;
  wire tmp3269;
  wire tmp3270;
  wire tmp3271;
  wire tmp3272;
  wire tmp3273;
  wire tmp3274;
  wire tmp3275;
  wire tmp3276;
  wire tmp3277;
  wire tmp3278;
  wire tmp3279;
  wire tmp3280;
  wire tmp3281;
  wire tmp3282;
  wire tmp3283;
  wire tmp3284;
  wire tmp3285;
  wire tmp3286;
  wire tmp3287;
  wire tmp3288;
  wire tmp3289;
  wire tmp3290;
  wire tmp3291;
  wire tmp3292;
  wire tmp3293;
  wire tmp3294;
  wire tmp3295;
  wire tmp3296;
  wire tmp3297;
  wire tmp3298;
  wire tmp3299;
  wire tmp3300;
  wire tmp3301;
  wire tmp3302;
  wire tmp3303;
  wire tmp3304;
  wire tmp3305;
  wire tmp3306;
  wire tmp3307;
  wire tmp3308;
  wire tmp3309;
  wire tmp3310;
  wire tmp3311;
  wire tmp3312;
  wire tmp3313;
  wire tmp3314;
  wire tmp3315;
  wire tmp3316;
  wire tmp3317;
  wire tmp3318;
  wire tmp3319;
  wire tmp3320;
  wire tmp3321;
  wire tmp3322;
  wire tmp3323;
  wire tmp3324;
  wire tmp3325;
  wire tmp3326;
  wire tmp3327;
  wire tmp3328;
  wire tmp3329;
  wire tmp3330;
  wire tmp3331;
  wire tmp3332;
  wire tmp3333;
  wire tmp3334;
  wire tmp3335;
  wire tmp3336;
  wire tmp3337;
  wire tmp3338;
  wire tmp3339;
  wire tmp3340;
  wire tmp3341;
  wire tmp3342;
  wire tmp3343;
  wire tmp3344;
  wire tmp3345;
  wire tmp3346;
  wire tmp3347;
  wire tmp3348;
  wire tmp3349;
  wire tmp3350;
  wire tmp3351;
  wire tmp3352;
  wire tmp3353;
  wire tmp3354;
  wire tmp3355;
  wire tmp3356;
  wire tmp3357;
  wire tmp3358;
  wire tmp3359;
  wire tmp3360;
  wire tmp3361;
  wire tmp3362;
  wire tmp3363;
  wire tmp3364;
  wire tmp3365;
  wire tmp3366;
  wire tmp3367;
  wire tmp3368;
  wire tmp3369;
  wire tmp3370;
  wire tmp3371;
  wire tmp3372;
  wire tmp3373;
  wire tmp3374;
  wire tmp3375;
  wire tmp3376;
  wire tmp3377;
  wire tmp3378;
  wire tmp3379;
  wire tmp3380;
  wire tmp3381;
  wire tmp3382;
  wire tmp3383;
  wire tmp3384;
  wire tmp3385;
  wire tmp3386;
  wire tmp3387;
  wire tmp3388;
  wire tmp3389;
  wire tmp3390;
  wire tmp3391;
  wire tmp3392;
  wire tmp3393;
  wire tmp3394;
  wire tmp3395;
  wire tmp3396;
  wire tmp3397;
  wire tmp3398;
  wire tmp3399;
  wire tmp3400;
  wire tmp3401;
  wire tmp3402;
  wire tmp3403;
  wire tmp3404;
  wire tmp3405;
  wire tmp3406;
  wire tmp3407;
  wire tmp3408;
  wire tmp3409;
  wire tmp3410;
  wire tmp3411;
  wire tmp3412;
  wire tmp3413;
  wire tmp3414;
  wire tmp3415;
  wire tmp3416;
  wire tmp3417;
  wire tmp3418;
  wire tmp3419;
  wire tmp3420;
  wire tmp3421;
  wire tmp3422;
  wire tmp3423;
  wire tmp3424;
  wire tmp3425;
  wire tmp3426;
  wire tmp3427;
  wire tmp3428;
  wire tmp3429;
  wire tmp3430;
  wire tmp3431;
  wire tmp3432;
  wire tmp3433;
  wire tmp3434;
  wire tmp3435;
  wire tmp3436;
  wire tmp3437;
  wire tmp3438;
  wire tmp3439;
  wire tmp3440;
  wire tmp3441;
  wire tmp3442;
  wire tmp3443;
  wire tmp3444;
  wire tmp3445;
  wire tmp3446;
  wire tmp3447;
  wire tmp3448;
  wire tmp3449;
  wire tmp3450;
  wire tmp3451;
  wire tmp3452;
  wire tmp3453;
  wire tmp3454;
  wire tmp3455;
  wire tmp3456;
  wire tmp3457;
  wire tmp3458;
  wire tmp3459;
  wire tmp3460;
  wire tmp3461;
  wire tmp3462;
  wire tmp3463;
  wire tmp3464;
  wire tmp3465;
  wire tmp3466;
  wire tmp3467;
  wire tmp3468;
  wire tmp3469;
  wire tmp3470;
  wire tmp3471;
  wire tmp3472;
  wire tmp3473;
  wire tmp3474;
  wire tmp3475;
  wire tmp3476;
  wire tmp3477;
  wire tmp3478;
  wire tmp3479;
  wire tmp3480;
  wire tmp3481;
  wire tmp3482;
  wire tmp3483;
  wire tmp3484;
  wire tmp3485;
  wire tmp3486;
  wire tmp3487;
  wire tmp3488;
  wire tmp3489;
  wire tmp3490;
  wire tmp3491;
  wire tmp3492;
  wire tmp3493;
  wire tmp3494;
  wire tmp3495;
  wire tmp3496;
  wire tmp3497;
  wire tmp3498;
  wire tmp3499;
  wire tmp3500;
  wire tmp3501;
  wire tmp3502;
  wire tmp3503;
  wire tmp3504;
  wire tmp3505;
  wire tmp3506;
  wire tmp3507;
  wire tmp3508;
  wire tmp3509;
  wire tmp3510;
  wire tmp3511;
  wire tmp3512;
  wire tmp3513;
  wire tmp3514;
  wire tmp3515;
  wire tmp3516;
  wire tmp3517;
  wire tmp3518;
  wire tmp3519;
  wire tmp3520;
  wire tmp3521;
  wire tmp3522;
  wire tmp3523;
  wire tmp3524;
  wire tmp3525;
  wire tmp3526;
  wire tmp3527;
  wire tmp3528;
  wire tmp3529;
  wire tmp3530;
  wire tmp3531;
  wire tmp3532;
  wire tmp3533;
  wire tmp3534;
  wire tmp3535;
  wire tmp3536;
  wire tmp3537;
  wire tmp3538;
  wire tmp3539;
  wire tmp3540;
  wire tmp3541;
  wire tmp3542;
  wire tmp3543;
  wire tmp3544;
  wire tmp3545;
  wire tmp3546;
  wire tmp3547;
  wire tmp3548;
  wire tmp3549;
  wire tmp3550;
  wire tmp3551;
  wire tmp3552;
  wire tmp3553;
  wire tmp3554;
  wire tmp3555;
  wire tmp3556;
  wire tmp3557;
  wire tmp3558;
  wire tmp3559;
  wire tmp3560;
  wire tmp3561;
  wire tmp3562;
  wire tmp3563;
  wire tmp3564;
  wire tmp3565;
  wire tmp3566;
  wire tmp3567;
  wire tmp3568;
  wire tmp3569;
  wire tmp3570;
  wire tmp3571;
  wire tmp3572;
  wire tmp3573;
  wire tmp3574;
  wire tmp3575;
  wire tmp3576;
  wire tmp3577;
  wire tmp3578;
  wire tmp3579;
  wire tmp3580;
  wire tmp3581;
  wire tmp3582;
  wire tmp3583;
  wire tmp3584;
  wire tmp3585;
  wire tmp3586;
  wire tmp3587;
  wire tmp3588;
  wire tmp3589;
  wire tmp3590;
  wire tmp3591;
  wire tmp3592;
  wire tmp3593;
  wire tmp3594;
  wire tmp3595;
  wire tmp3596;
  wire tmp3597;
  wire tmp3598;
  wire tmp3599;
  wire tmp3600;
  wire tmp3601;
  wire tmp3602;
  wire tmp3603;
  wire tmp3604;
  wire tmp3605;
  wire tmp3606;
  wire tmp3607;
  wire tmp3608;
  wire tmp3609;
  wire tmp3610;
  wire tmp3611;
  wire tmp3612;
  wire tmp3613;
  wire tmp3614;
  wire tmp3615;
  wire tmp3616;
  wire tmp3617;
  wire tmp3618;
  wire tmp3619;
  wire tmp3620;
  wire tmp3621;
  wire tmp3622;
  wire tmp3623;
  wire tmp3624;
  wire tmp3625;
  wire tmp3626;
  wire tmp3627;
  wire tmp3628;
  wire tmp3629;
  wire tmp3630;
  wire tmp3631;
  wire tmp3632;
  wire tmp3633;
  wire tmp3634;
  wire tmp3635;
  wire tmp3636;
  wire tmp3637;
  wire tmp3638;
  wire tmp3639;
  wire tmp3640;
  wire tmp3641;
  wire tmp3642;
  wire tmp3643;
  wire tmp3644;
  wire tmp3645;
  wire tmp3646;
  wire tmp3647;
  wire tmp3648;
  wire tmp3649;
  wire tmp3650;
  wire tmp3651;
  wire tmp3652;
  wire tmp3653;
  wire tmp3654;
  wire tmp3655;
  wire tmp3656;
  wire tmp3657;
  wire tmp3658;
  wire tmp3659;
  wire tmp3660;
  wire tmp3661;
  wire tmp3662;
  wire tmp3663;
  wire tmp3664;
  wire tmp3665;
  wire tmp3666;
  wire tmp3667;
  wire tmp3668;
  wire tmp3669;
  wire tmp3670;
  wire tmp3671;
  wire tmp3672;
  wire tmp3673;
  wire tmp3674;
  wire tmp3675;
  wire tmp3676;
  wire tmp3677;
  wire tmp3678;
  wire tmp3679;
  wire tmp3680;
  wire tmp3681;
  wire tmp3682;
  wire tmp3683;
  wire tmp3684;
  wire tmp3685;
  wire tmp3686;
  wire tmp3687;
  wire tmp3688;
  wire tmp3689;
  wire tmp3690;
  wire tmp3691;
  wire tmp3692;
  wire tmp3693;
  wire tmp3694;
  wire tmp3695;
  wire tmp3696;
  wire tmp3697;
  wire tmp3698;
  wire tmp3699;
  wire tmp3700;
  wire tmp3701;
  wire tmp3702;
  wire tmp3703;
  wire tmp3704;
  wire tmp3705;
  wire tmp3706;
  wire tmp3707;
  wire tmp3708;
  wire tmp3709;
  wire tmp3710;
  wire tmp3711;
  wire tmp3712;
  wire tmp3713;
  wire tmp3714;
  wire tmp3715;
  wire tmp3716;
  wire tmp3717;
  wire tmp3718;
  wire tmp3719;
  wire tmp3720;
  wire tmp3721;
  wire tmp3722;
  wire tmp3723;
  wire tmp3724;
  wire tmp3725;
  wire tmp3726;
  wire tmp3727;
  wire tmp3728;
  wire tmp3729;
  wire tmp3730;
  wire tmp3731;
  wire tmp3732;
  wire tmp3733;
  wire tmp3734;
  wire tmp3735;
  wire tmp3736;
  wire tmp3737;
  wire tmp3738;
  wire tmp3739;
  wire tmp3740;
  wire tmp3741;
  wire tmp3742;
  wire tmp3743;
  wire tmp3744;
  wire tmp3745;
  wire tmp3746;
  wire tmp3747;
  wire tmp3748;
  wire tmp3749;
  wire tmp3750;
  wire tmp3751;
  wire tmp3752;
  wire tmp3753;
  wire tmp3754;
  wire tmp3755;
  wire tmp3756;
  wire tmp3757;
  wire tmp3758;
  wire tmp3759;
  wire tmp3760;
  wire tmp3761;
  wire tmp3762;
  wire tmp3763;
  wire tmp3764;
  wire tmp3765;
  wire tmp3766;
  wire tmp3767;
  wire tmp3768;
  wire tmp3769;
  wire tmp3770;
  wire tmp3771;
  wire tmp3772;
  wire tmp3773;
  wire tmp3774;
  wire tmp3775;
  wire tmp3776;
  wire tmp3777;
  wire tmp3778;
  wire tmp3779;
  wire tmp3780;
  wire tmp3781;
  wire tmp3782;
  wire tmp3783;
  wire tmp3784;
  wire tmp3785;
  wire tmp3786;
  wire tmp3787;
  wire tmp3788;
  wire tmp3789;
  wire tmp3790;
  wire tmp3791;
  wire tmp3792;
  wire tmp3793;
  wire tmp3794;
  wire tmp3795;
  wire tmp3796;
  wire tmp3797;
  wire tmp3798;
  wire tmp3799;
  wire tmp3800;
  wire tmp3801;
  wire tmp3802;
  wire tmp3803;
  wire tmp3804;
  wire tmp3805;
  wire tmp3806;
  wire tmp3807;
  wire tmp3808;
  wire tmp3809;
  wire tmp3810;
  wire tmp3811;
  wire tmp3812;
  wire tmp3813;
  wire tmp3814;
  wire tmp3815;
  wire tmp3816;
  wire tmp3817;
  wire tmp3818;
  wire tmp3819;
  wire tmp3820;
  wire tmp3821;
  wire tmp3822;
  wire tmp3823;
  wire tmp3824;
  wire tmp3825;
  wire tmp3826;
  wire tmp3827;
  wire tmp3828;
  wire tmp3829;
  wire tmp3830;
  wire tmp3831;
  wire tmp3832;
  wire tmp3833;
  wire tmp3834;
  wire tmp3835;
  wire tmp3836;
  wire tmp3837;
  wire tmp3838;
  wire tmp3839;
  wire tmp3840;
  wire tmp3841;
  wire tmp3842;
  wire tmp3843;
  wire tmp3844;
  wire tmp3845;
  wire tmp3846;
  wire tmp3847;
  wire tmp3848;
  wire tmp3849;
  wire tmp3850;
  wire tmp3851;
  wire tmp3852;
  wire tmp3853;
  wire tmp3854;
  wire tmp3855;
  wire tmp3856;
  wire tmp3857;
  wire tmp3858;
  wire tmp3859;
  wire tmp3860;
  wire tmp3861;
  wire tmp3862;
  wire tmp3863;
  wire tmp3864;
  wire tmp3865;
  wire tmp3866;
  wire tmp3867;
  wire tmp3868;
  wire tmp3869;
  wire tmp3870;
  wire tmp3871;
  wire tmp3872;
  wire tmp3873;
  wire tmp3874;
  wire tmp3875;
  wire tmp3876;
  wire tmp3877;
  wire tmp3878;
  wire tmp3879;
  wire tmp3880;
  wire tmp3881;
  wire tmp3882;
  wire tmp3883;
  wire tmp3884;
  wire tmp3885;
  wire tmp3886;
  wire tmp3887;
  wire tmp3888;
  wire tmp3889;
  wire tmp3890;
  wire tmp3891;
  wire tmp3892;
  wire tmp3893;
  wire tmp3894;
  wire tmp3895;
  wire tmp3896;
  wire tmp3897;
  wire tmp3898;
  wire tmp3899;
  wire tmp3900;
  wire tmp3901;
  wire tmp3902;
  wire tmp3903;
  wire tmp3904;
  wire tmp3905;
  wire tmp3906;
  wire tmp3907;
  wire tmp3908;
  wire tmp3909;
  wire tmp3910;
  wire tmp3911;
  wire tmp3912;
  wire tmp3913;
  wire tmp3914;
  wire tmp3915;
  wire tmp3916;
  wire tmp3917;
  wire tmp3918;
  wire tmp3919;
  wire tmp3920;
  wire tmp3921;
  wire tmp3922;
  wire tmp3923;
  wire tmp3924;
  wire tmp3925;
  wire tmp3926;
  wire tmp3927;
  wire tmp3928;
  wire tmp3929;
  wire tmp3930;
  wire tmp3931;
  wire tmp3932;
  wire tmp3933;
  wire tmp3934;
  wire tmp3935;
  wire tmp3936;
  wire tmp3937;
  wire tmp3938;
  wire tmp3939;
  wire tmp3940;
  wire tmp3941;
  wire tmp3942;
  wire tmp3943;
  wire tmp3944;
  wire tmp3945;
  wire tmp3946;
  wire tmp3947;
  wire tmp3948;
  wire tmp3949;
  wire tmp3950;
  wire tmp3951;
  wire tmp3952;
  wire tmp3953;
  wire tmp3954;
  wire tmp3955;
  wire tmp3956;
  wire tmp3957;
  wire tmp3958;
  wire tmp3959;
  wire tmp3960;
  wire tmp3961;
  wire tmp3962;
  wire tmp3963;
  wire tmp3964;
  wire tmp3965;
  wire tmp3966;
  wire tmp3967;
  wire tmp3968;
  wire tmp3969;
  wire tmp3970;
  wire tmp3971;
  wire tmp3972;
  wire tmp3973;
  wire tmp3974;
  wire tmp3975;
  wire tmp3976;
  wire tmp3977;
  wire tmp3978;
  wire tmp3979;
  wire tmp3980;
  wire tmp3981;
  wire tmp3982;
  wire tmp3983;
  wire tmp3984;
  wire tmp3985;
  wire tmp3986;
  wire tmp3987;
  wire tmp3988;
  wire tmp3989;
  wire tmp3990;
  wire tmp3991;
  wire tmp3992;
  wire tmp3993;
  wire tmp3994;
  wire tmp3995;
  wire tmp3996;
  wire tmp3997;
  wire tmp3998;
  wire tmp3999;
  wire tmp4000;
  wire tmp4001;
  wire tmp4002;
  wire tmp4003;
  wire tmp4004;
  wire tmp4005;
  wire tmp4006;
  wire tmp4007;
  wire tmp4008;
  wire tmp4009;
  wire tmp4010;
  wire tmp4011;
  wire tmp4012;
  wire tmp4013;
  wire tmp4014;
  wire tmp4015;
  wire tmp4016;
  wire tmp4017;
  wire tmp4018;
  wire tmp4019;
  wire tmp4020;
  wire tmp4021;
  wire tmp4022;
  wire tmp4023;
  wire tmp4024;
  wire tmp4025;
  wire tmp4026;
  wire tmp4027;
  wire tmp4028;
  wire tmp4029;
  wire tmp4030;
  wire tmp4031;
  wire tmp4032;
  wire tmp4033;
  wire tmp4034;
  wire tmp4035;
  wire tmp4036;
  wire tmp4037;
  wire tmp4038;
  wire tmp4039;
  wire tmp4040;
  wire tmp4041;
  wire tmp4042;
  wire tmp4043;
  wire tmp4044;
  wire tmp4045;
  wire tmp4046;
  wire tmp4047;
  wire tmp4048;
  wire tmp4049;
  wire tmp4050;
  wire tmp4051;
  wire tmp4052;
  wire tmp4053;
  wire tmp4054;
  wire tmp4055;
  wire tmp4056;
  wire tmp4057;
  wire tmp4058;
  wire tmp4059;
  wire tmp4060;
  wire tmp4061;
  wire tmp4062;
  wire tmp4063;
  wire tmp4064;
  wire tmp4065;
  wire tmp4066;
  wire tmp4067;
  wire tmp4068;
  wire tmp4069;
  wire tmp4070;
  wire tmp4071;
  wire tmp4072;
  wire tmp4073;
  wire tmp4074;
  wire tmp4075;
  wire tmp4076;
  wire tmp4077;
  wire tmp4078;
  wire tmp4079;
  wire tmp4080;
  wire tmp4081;
  wire tmp4082;
  wire tmp4083;
  wire tmp4084;
  wire tmp4085;
  wire tmp4086;
  wire tmp4087;
  wire tmp4088;
  wire tmp4089;
  wire tmp4090;
  wire tmp4091;
  wire tmp4092;
  wire tmp4093;
  wire tmp4094;
  wire tmp4095;
  wire tmp4096;
  wire tmp4097;
  wire tmp4098;
  wire tmp4099;
  wire tmp4100;
  wire tmp4101;
  wire tmp4102;
  wire tmp4103;
  wire tmp4104;
  wire tmp4105;
  wire tmp4106;
  wire tmp4107;
  wire tmp4108;
  wire tmp4109;
  wire tmp4110;
  wire tmp4111;
  wire tmp4112;
  wire tmp4113;
  wire tmp4114;
  wire tmp4115;
  wire tmp4116;
  wire tmp4117;
  wire tmp4118;
  wire tmp4119;
  wire tmp4120;
  wire tmp4121;
  wire tmp4122;
  wire tmp4123;
  wire tmp4124;
  wire tmp4125;
  wire tmp4126;
  wire tmp4127;
  wire tmp4128;
  wire tmp4129;
  wire tmp4130;
  wire tmp4131;
  wire tmp4132;
  wire tmp4133;
  wire tmp4134;
  wire tmp4135;
  wire tmp4136;
  wire tmp4137;
  wire tmp4138;
  wire tmp4139;
  wire tmp4140;
  wire tmp4141;
  wire tmp4142;
  wire tmp4143;
  wire tmp4144;
  wire tmp4145;
  wire tmp4146;
  wire tmp4147;
  wire tmp4148;
  wire tmp4149;
  wire tmp4150;
  wire tmp4151;
  wire tmp4152;
  wire tmp4153;
  wire tmp4154;
  wire tmp4155;
  wire tmp4156;
  wire tmp4157;
  wire tmp4158;
  wire tmp4159;
  wire tmp4160;
  wire tmp4161;
  wire tmp4162;
  wire tmp4163;
  wire tmp4164;
  wire tmp4165;
  wire tmp4166;
  wire tmp4167;
  wire tmp4168;
  wire tmp4169;
  wire tmp4170;
  wire tmp4171;
  wire tmp4172;
  wire tmp4173;
  wire tmp4174;
  wire tmp4175;
  wire tmp4176;
  wire tmp4177;
  wire tmp4178;
  wire tmp4179;
  wire tmp4180;
  wire tmp4181;
  wire tmp4182;
  wire tmp4183;
  wire tmp4184;
  wire tmp4185;
  wire tmp4186;
  wire tmp4187;
  wire tmp4188;
  wire tmp4189;
  wire tmp4190;
  wire tmp4191;
  wire tmp4192;
  wire tmp4193;
  wire tmp4194;
  wire tmp4195;
  wire tmp4196;
  wire tmp4197;
  wire tmp4198;
  wire tmp4199;
  wire tmp4200;
  wire tmp4201;
  wire tmp4202;
  wire tmp4203;
  wire tmp4204;
  wire tmp4205;
  wire tmp4206;
  wire tmp4207;
  wire tmp4208;
  wire tmp4209;
  wire tmp4210;
  wire tmp4211;
  wire tmp4212;
  wire tmp4213;
  wire tmp4214;
  wire tmp4215;
  wire tmp4216;
  wire tmp4217;
  wire tmp4218;
  wire tmp4219;
  wire tmp4220;
  wire tmp4221;
  wire tmp4222;
  wire tmp4223;
  wire tmp4224;
  wire tmp4225;
  wire tmp4226;
  wire tmp4227;
  wire tmp4228;
  wire tmp4229;
  wire tmp4230;
  wire tmp4231;
  wire tmp4232;
  wire tmp4233;
  wire tmp4234;
  wire tmp4235;
  wire tmp4236;
  wire tmp4237;
  wire tmp4238;
  wire tmp4239;
  wire tmp4240;
  wire tmp4241;
  wire tmp4242;
  wire tmp4243;
  wire tmp4244;
  wire tmp4245;
  wire tmp4246;
  wire tmp4247;
  wire tmp4248;
  wire tmp4249;
  wire tmp4250;
  wire tmp4251;
  wire tmp4252;
  wire tmp4253;
  wire tmp4254;
  wire tmp4255;
  wire tmp4256;
  wire tmp4257;
  wire tmp4258;
  wire tmp4259;
  wire tmp4260;
  wire tmp4261;
  wire tmp4262;
  wire tmp4263;
  wire tmp4264;
  wire tmp4265;
  wire tmp4266;
  wire tmp4267;
  wire tmp4268;
  wire tmp4269;
  wire tmp4270;
  wire tmp4271;
  wire tmp4272;
  wire tmp4273;
  wire tmp4274;
  wire tmp4275;
  wire tmp4276;
  wire tmp4277;
  wire tmp4278;
  wire tmp4279;
  wire tmp4280;
  wire tmp4281;
  wire tmp4282;
  wire tmp4283;
  wire tmp4284;
  wire tmp4285;
  wire tmp4286;
  wire tmp4287;
  wire tmp4288;
  wire tmp4289;
  wire tmp4290;
  wire tmp4291;
  wire tmp4292;
  wire tmp4293;
  wire tmp4294;
  wire tmp4295;
  wire tmp4296;
  wire tmp4297;
  wire tmp4298;
  wire tmp4299;
  wire tmp4300;
  wire tmp4301;
  wire tmp4302;
  wire tmp4303;
  wire tmp4304;
  wire tmp4305;
  wire tmp4306;
  wire tmp4307;
  wire tmp4308;
  wire tmp4309;
  wire tmp4310;
  wire tmp4311;
  wire tmp4312;
  wire tmp4313;
  wire tmp4314;
  wire tmp4315;
  wire tmp4316;
  wire tmp4317;
  wire tmp4318;
  wire tmp4319;
  wire tmp4320;
  wire tmp4321;
  wire tmp4322;
  wire tmp4323;
  wire tmp4324;
  wire tmp4325;
  wire tmp4326;
  wire tmp4327;
  wire tmp4328;
  wire tmp4329;
  wire tmp4330;
  wire tmp4331;
  wire tmp4332;
  wire tmp4333;
  wire tmp4334;
  wire tmp4335;
  wire tmp4336;
  wire tmp4337;
  wire tmp4338;
  wire tmp4339;
  wire tmp4340;
  wire tmp4341;
  wire tmp4342;
  wire tmp4343;
  wire tmp4344;
  wire tmp4345;
  wire tmp4346;
  wire tmp4347;
  wire tmp4348;
  wire tmp4349;
  wire tmp4350;
  wire tmp4351;
  wire tmp4352;
  wire tmp4353;
  wire tmp4354;
  wire tmp4355;
  wire tmp4356;
  wire tmp4357;
  wire tmp4358;
  wire tmp4359;
  wire tmp4360;
  wire tmp4361;
  wire tmp4362;
  wire tmp4363;
  wire tmp4364;
  wire tmp4365;
  wire tmp4366;
  wire tmp4367;
  wire tmp4368;
  wire tmp4369;
  wire tmp4370;
  wire tmp4371;
  wire tmp4372;
  wire tmp4373;
  wire tmp4374;
  wire tmp4375;
  wire tmp4376;
  wire tmp4377;
  wire tmp4378;
  wire tmp4379;
  wire tmp4380;
  wire tmp4381;
  wire tmp4382;
  wire tmp4383;
  wire tmp4384;
  wire tmp4385;
  wire tmp4386;
  wire tmp4387;
  wire tmp4388;
  wire tmp4389;
  wire tmp4390;
  wire tmp4391;
  wire tmp4392;
  wire tmp4393;
  wire tmp4394;
  wire tmp4395;
  wire tmp4396;
  wire tmp4397;
  wire tmp4398;
  wire tmp4399;
  wire tmp4400;
  wire tmp4401;
  wire tmp4402;
  wire tmp4403;
  wire tmp4404;
  wire tmp4405;
  wire tmp4406;
  wire tmp4407;
  wire tmp4408;
  wire tmp4409;
  wire tmp4410;
  wire tmp4411;
  wire tmp4412;
  wire tmp4413;
  wire tmp4414;
  wire tmp4415;
  wire tmp4416;
  wire tmp4417;
  wire tmp4418;
  wire tmp4419;
  wire tmp4420;
  wire tmp4421;
  wire tmp4422;
  wire tmp4423;
  wire tmp4424;
  wire tmp4425;
  wire tmp4426;
  wire tmp4427;
  wire tmp4428;
  wire tmp4429;
  wire tmp4430;
  wire tmp4431;
  wire tmp4432;
  wire tmp4433;
  wire tmp4434;
  wire tmp4435;
  wire tmp4436;
  wire tmp4437;
  wire tmp4438;
  wire tmp4439;
  wire tmp4440;
  wire tmp4441;
  wire tmp4442;
  wire tmp4443;
  wire tmp4444;
  wire tmp4445;
  wire tmp4446;
  wire tmp4447;
  wire tmp4448;
  wire tmp4449;
  wire tmp4450;
  wire tmp4451;
  wire tmp4452;
  wire tmp4453;
  wire tmp4454;
  wire tmp4455;
  wire tmp4456;
  wire tmp4457;
  wire tmp4458;
  wire tmp4459;
  wire tmp4460;
  wire tmp4461;
  wire tmp4462;
  wire tmp4463;
  wire tmp4464;
  wire tmp4465;
  wire tmp4466;
  wire tmp4467;
  wire tmp4468;
  wire tmp4469;
  wire tmp4470;
  wire tmp4471;
  wire tmp4472;
  wire tmp4473;
  wire tmp4474;
  wire tmp4475;
  wire tmp4476;
  wire tmp4477;
  wire tmp4478;
  wire tmp4479;
  wire tmp4480;
  wire tmp4481;
  wire tmp4482;
  wire tmp4483;
  wire tmp4484;
  wire tmp4485;
  wire tmp4486;
  wire tmp4487;
  wire tmp4488;
  wire tmp4489;
  wire tmp4490;
  wire tmp4491;
  wire tmp4492;
  wire tmp4493;
  wire tmp4494;
  wire tmp4495;
  wire tmp4496;
  wire tmp4497;
  wire tmp4498;
  wire tmp4499;
  wire tmp4500;
  wire tmp4501;
  wire tmp4502;
  wire tmp4503;
  wire tmp4504;
  wire tmp4505;
  wire tmp4506;
  wire tmp4507;
  wire tmp4508;
  wire tmp4509;
  wire tmp4510;
  wire tmp4511;
  wire tmp4512;
  wire tmp4513;
  wire tmp4514;
  wire tmp4515;
  wire tmp4516;
  wire tmp4517;
  wire tmp4518;
  wire tmp4519;
  wire tmp4520;
  wire tmp4521;
  wire tmp4522;
  wire tmp4523;
  wire tmp4524;
  wire tmp4525;
  wire tmp4526;
  wire tmp4527;
  wire tmp4528;
  wire tmp4529;
  wire tmp4530;
  wire tmp4531;
  wire tmp4532;
  wire tmp4533;
  wire tmp4534;
  wire tmp4535;
  wire tmp4536;
  wire tmp4537;
  wire tmp4538;
  wire tmp4539;
  wire tmp4540;
  wire tmp4541;
  wire tmp4542;
  wire tmp4543;
  wire tmp4544;
  wire tmp4545;
  wire tmp4546;
  wire tmp4547;
  wire tmp4548;
  wire tmp4549;
  wire tmp4550;
  wire tmp4551;
  wire tmp4552;
  wire tmp4553;
  wire tmp4554;
  wire tmp4555;
  wire tmp4556;
  wire tmp4557;
  wire tmp4558;
  wire tmp4559;
  wire tmp4560;
  wire tmp4561;
  wire tmp4562;
  wire tmp4563;
  wire tmp4564;
  wire tmp4565;
  wire tmp4566;
  wire tmp4567;
  wire tmp4568;
  wire tmp4569;
  wire tmp4570;
  wire tmp4571;
  wire tmp4572;
  wire tmp4573;
  wire tmp4574;
  wire tmp4575;
  wire tmp4576;
  wire tmp4577;
  wire tmp4578;
  wire tmp4579;
  wire tmp4580;
  wire tmp4581;
  wire tmp4582;
  wire tmp4583;
  wire tmp4584;
  wire tmp4585;
  wire tmp4586;
  wire tmp4587;
  wire tmp4588;
  wire tmp4589;
  wire tmp4590;
  wire tmp4591;
  wire tmp4592;
  wire tmp4593;
  wire tmp4594;
  wire tmp4595;
  wire tmp4596;
  wire tmp4597;
  wire tmp4598;
  wire tmp4599;
  wire tmp4600;
  wire tmp4601;
  wire tmp4602;
  wire tmp4603;
  wire tmp4604;
  wire tmp4605;
  wire tmp4606;
  wire tmp4607;
  wire tmp4608;
  wire tmp4609;
  wire tmp4610;
  wire tmp4611;
  wire tmp4612;
  wire tmp4613;
  wire tmp4614;
  wire tmp4615;
  wire tmp4616;
  wire tmp4617;
  wire tmp4618;
  wire tmp4619;
  wire tmp4620;
  wire tmp4621;
  wire tmp4622;
  wire tmp4623;
  wire tmp4624;
  wire tmp4625;
  wire tmp4626;
  wire tmp4627;
  wire tmp4628;
  wire tmp4629;
  wire tmp4630;
  wire tmp4631;
  wire tmp4632;
  wire tmp4633;
  wire tmp4634;
  wire tmp4635;
  wire tmp4636;
  wire tmp4637;
  wire tmp4638;
  wire tmp4639;
  wire tmp4640;
  wire tmp4641;
  wire tmp4642;
  wire tmp4643;
  wire tmp4644;
  wire tmp4645;
  wire tmp4646;
  wire tmp4647;
  wire tmp4648;
  wire tmp4649;
  wire tmp4650;
  wire tmp4651;
  wire tmp4652;
  wire tmp4653;
  wire tmp4654;
  wire tmp4655;
  wire tmp4656;
  wire tmp4657;
  wire tmp4658;
  wire tmp4659;
  wire tmp4660;
  wire tmp4661;
  wire tmp4662;
  wire tmp4663;
  wire tmp4664;
  wire tmp4665;
  wire tmp4666;
  wire tmp4667;
  wire tmp4668;
  wire tmp4669;
  wire tmp4670;
  wire tmp4671;
  wire tmp4672;
  wire tmp4673;
  wire tmp4674;
  wire tmp4675;
  wire tmp4676;
  wire tmp4677;
  wire tmp4678;
  wire tmp4679;
  wire tmp4680;
  wire tmp4681;
  wire tmp4682;
  wire tmp4683;
  wire tmp4684;
  wire tmp4685;
  wire tmp4686;
  wire tmp4687;
  wire tmp4688;
  wire tmp4689;
  wire tmp4690;
  wire tmp4691;
  wire tmp4692;
  wire tmp4693;
  wire tmp4694;
  wire tmp4695;
  wire tmp4696;
  wire tmp4697;
  wire tmp4698;
  wire tmp4699;
  wire tmp4700;
  wire tmp4701;
  wire tmp4702;
  wire tmp4703;
  wire tmp4704;
  wire tmp4705;
  wire tmp4706;
  wire tmp4707;
  wire tmp4708;
  wire tmp4709;
  wire tmp4710;
  wire tmp4711;
  wire tmp4712;
  wire tmp4713;
  wire tmp4714;
  wire tmp4715;
  wire tmp4716;
  wire tmp4717;
  wire tmp4718;
  wire tmp4719;
  wire tmp4720;
  wire tmp4721;
  wire tmp4722;
  wire tmp4723;
  wire tmp4724;
  wire tmp4725;
  wire tmp4726;
  wire tmp4727;
  wire tmp4728;
  wire tmp4729;
  wire tmp4730;
  wire tmp4731;
  wire tmp4732;
  wire tmp4733;
  wire tmp4734;
  wire tmp4735;
  wire tmp4736;
  wire tmp4737;
  wire tmp4738;
  wire tmp4739;
  wire tmp4740;
  wire tmp4741;
  wire tmp4742;
  wire tmp4743;
  wire tmp4744;
  wire tmp4745;
  wire tmp4746;
  wire tmp4747;
  wire tmp4748;
  wire tmp4749;
  wire tmp4750;
  wire tmp4751;
  wire tmp4752;
  wire tmp4753;
  wire tmp4754;
  wire tmp4755;
  wire tmp4756;
  wire tmp4757;
  wire tmp4758;
  wire tmp4759;
  wire tmp4760;
  wire tmp4761;
  wire tmp4762;
  wire tmp4763;
  wire tmp4764;
  wire tmp4765;
  wire tmp4766;
  wire tmp4767;
  wire tmp4768;
  wire tmp4769;
  wire tmp4770;
  wire tmp4771;
  wire tmp4772;
  wire tmp4773;
  wire tmp4774;
  wire tmp4775;
  wire tmp4776;
  wire tmp4777;
  wire tmp4778;
  wire tmp4779;
  wire tmp4780;
  wire tmp4781;
  wire tmp4782;
  wire tmp4783;
  wire tmp4784;
  wire tmp4785;
  wire tmp4786;
  wire tmp4787;
  wire tmp4788;
  wire tmp4789;
  wire tmp4790;
  wire tmp4791;
  wire tmp4792;
  wire tmp4793;
  wire tmp4794;
  wire tmp4795;
  wire tmp4796;
  wire tmp4797;
  wire tmp4798;
  wire tmp4799;
  wire tmp4800;
  wire tmp4801;
  wire tmp4802;
  wire tmp4803;
  wire tmp4804;
  wire tmp4805;
  wire tmp4806;
  wire tmp4807;
  wire tmp4808;
  wire tmp4809;
  wire tmp4810;
  wire tmp4811;
  wire tmp4812;
  wire tmp4813;
  wire tmp4814;
  wire tmp4815;
  wire tmp4816;
  wire tmp4817;
  wire tmp4818;
  wire tmp4819;
  wire tmp4820;
  wire tmp4821;
  wire tmp4822;
  wire tmp4823;
  wire tmp4824;
  wire tmp4825;
  wire tmp4826;
  wire tmp4827;
  wire tmp4828;
  wire tmp4829;
  wire tmp4830;
  wire tmp4831;
  wire tmp4832;
  wire tmp4833;
  wire tmp4834;
  wire tmp4835;
  wire tmp4836;
  wire tmp4837;
  wire tmp4838;
  wire tmp4839;
  wire tmp4840;
  wire tmp4841;
  wire tmp4842;
  wire tmp4843;
  wire tmp4844;
  wire tmp4845;
  wire tmp4846;
  wire tmp4847;
  wire tmp4848;
  wire tmp4849;
  wire tmp4850;
  wire tmp4851;
  wire tmp4852;
  wire tmp4853;
  wire tmp4854;
  wire tmp4855;
  wire tmp4856;
  wire tmp4857;
  wire tmp4858;
  wire tmp4859;
  wire tmp4860;
  wire tmp4861;
  wire tmp4862;
  wire tmp4863;
  wire tmp4864;
  wire tmp4865;
  wire tmp4866;
  wire tmp4867;
  wire tmp4868;
  wire tmp4869;
  wire tmp4870;
  wire tmp4871;
  wire tmp4872;
  wire tmp4873;
  wire tmp4874;
  wire tmp4875;
  wire tmp4876;
  wire tmp4877;
  wire tmp4878;
  wire tmp4879;
  wire tmp4880;
  wire tmp4881;
  wire tmp4882;
  wire tmp4883;
  wire tmp4884;
  wire tmp4885;
  wire tmp4886;
  wire tmp4887;
  wire tmp4888;
  wire tmp4889;
  wire tmp4890;
  wire tmp4891;
  wire tmp4892;
  wire tmp4893;
  wire tmp4894;
  wire tmp4895;
  wire tmp4896;
  wire tmp4897;
  wire tmp4898;
  wire tmp4899;
  wire tmp4900;
  wire tmp4901;
  wire tmp4902;
  wire tmp4903;
  wire tmp4904;
  wire tmp4905;
  wire tmp4906;
  wire tmp4907;
  wire tmp4908;
  wire tmp4909;
  wire tmp4910;
  wire tmp4911;
  wire tmp4912;
  wire tmp4913;
  wire tmp4914;
  wire tmp4915;
  wire tmp4916;
  wire tmp4917;
  wire tmp4918;
  wire tmp4919;
  wire tmp4920;
  wire tmp4921;
  wire tmp4922;
  wire tmp4923;
  wire tmp4924;
  wire tmp4925;
  wire tmp4926;
  wire tmp4927;
  wire tmp4928;
  wire tmp4929;
  wire tmp4930;
  wire tmp4931;
  wire tmp4932;
  wire tmp4933;
  wire tmp4934;
  wire tmp4935;
  wire tmp4936;
  wire tmp4937;
  wire tmp4938;
  wire tmp4939;
  wire tmp4940;
  wire tmp4941;
  wire tmp4942;
  wire tmp4943;
  wire tmp4944;
  wire tmp4945;
  wire tmp4946;
  wire tmp4947;
  wire tmp4948;
  wire tmp4949;
  wire tmp4950;
  wire tmp4951;
  wire tmp4952;
  wire tmp4953;
  wire tmp4954;
  wire tmp4955;
  wire tmp4956;
  wire tmp4957;
  wire tmp4958;
  wire tmp4959;
  wire tmp4960;
  wire tmp4961;
  wire tmp4962;
  wire tmp4963;
  wire tmp4964;
  wire tmp4965;
  wire tmp4966;
  wire tmp4967;
  wire tmp4968;
  wire tmp4969;
  wire tmp4970;
  wire tmp4971;
  wire tmp4972;
  wire tmp4973;
  wire tmp4974;
  wire tmp4975;
  wire tmp4976;
  wire tmp4977;
  wire tmp4978;
  wire tmp4979;
  wire tmp4980;
  wire tmp4981;
  wire tmp4982;
  wire tmp4983;
  wire tmp4984;
  wire tmp4985;
  wire tmp4986;
  wire tmp4987;
  wire tmp4988;
  wire tmp4989;
  wire tmp4990;
  wire tmp4991;
  wire tmp4992;
  wire tmp4993;
  wire tmp4994;
  wire tmp4995;
  wire tmp4996;
  wire tmp4997;
  wire tmp4998;
  wire tmp4999;
  wire tmp5000;
  wire tmp5001;
  wire tmp5002;
  wire tmp5003;
  wire tmp5004;
  wire tmp5005;
  wire tmp5006;
  wire tmp5007;
  wire tmp5008;
  wire tmp5009;
  wire tmp5010;
  wire tmp5011;
  wire tmp5012;
  wire tmp5013;
  wire tmp5014;
  wire tmp5015;
  wire tmp5016;
  wire tmp5017;
  wire tmp5018;
  wire tmp5019;
  wire tmp5020;
  wire tmp5021;
  wire tmp5022;
  wire tmp5023;
  wire tmp5024;
  wire tmp5025;
  wire tmp5026;
  wire tmp5027;
  wire tmp5028;
  wire tmp5029;
  wire tmp5030;
  wire tmp5031;
  wire tmp5032;
  wire tmp5033;
  wire tmp5034;
  wire tmp5035;
  wire tmp5036;
  wire tmp5037;
  wire tmp5038;
  wire tmp5039;
  wire tmp5040;
  wire tmp5041;
  wire tmp5042;
  wire tmp5043;
  wire tmp5044;
  wire tmp5045;
  wire tmp5046;
  wire tmp5047;
  wire tmp5048;
  wire tmp5049;
  wire tmp5050;
  wire tmp5051;
  wire tmp5052;
  wire tmp5053;
  wire tmp5054;
  wire tmp5055;
  wire tmp5056;
  wire tmp5057;
  wire tmp5058;
  wire tmp5059;
  wire tmp5060;
  wire tmp5061;
  wire tmp5062;
  wire tmp5063;
  wire tmp5064;
  wire tmp5065;
  wire tmp5066;
  wire tmp5067;
  wire tmp5068;
  wire tmp5069;
  wire tmp5070;
  wire tmp5071;
  wire tmp5072;
  wire tmp5073;
  wire tmp5074;
  wire tmp5075;
  wire tmp5076;
  wire tmp5077;
  wire tmp5078;
  wire tmp5079;
  wire tmp5080;
  wire tmp5081;
  wire tmp5082;
  wire tmp5083;
  wire tmp5084;
  wire tmp5085;
  wire tmp5086;
  wire tmp5087;
  wire tmp5088;
  wire tmp5089;
  wire tmp5090;
  wire tmp5091;
  wire tmp5092;
  wire tmp5093;
  wire tmp5094;
  wire tmp5095;
  wire tmp5096;
  wire tmp5097;
  wire tmp5098;
  wire tmp5099;
  wire tmp5100;
  wire tmp5101;
  wire tmp5102;
  wire tmp5103;
  wire tmp5104;
  wire tmp5105;
  wire tmp5106;
  wire tmp5107;
  wire tmp5108;
  wire tmp5109;
  wire tmp5110;
  wire tmp5111;
  wire tmp5112;
  wire tmp5113;
  wire tmp5114;
  wire tmp5115;
  wire tmp5116;
  wire tmp5117;
  wire tmp5118;
  wire tmp5119;
  wire tmp5120;
  wire tmp5121;
  wire tmp5122;
  wire tmp5123;
  wire tmp5124;
  wire tmp5125;
  wire tmp5126;
  wire tmp5127;
  wire tmp5128;
  wire tmp5129;
  wire tmp5130;
  wire tmp5131;
  wire tmp5132;
  wire tmp5133;
  wire tmp5134;
  wire tmp5135;
  wire tmp5136;
  wire tmp5137;
  wire tmp5138;
  wire tmp5139;
  wire tmp5140;
  wire tmp5141;
  wire tmp5142;
  wire tmp5143;
  wire tmp5144;
  wire tmp5145;
  wire tmp5146;
  wire tmp5147;
  wire tmp5148;
  wire tmp5149;
  wire tmp5150;
  wire tmp5151;
  wire tmp5152;
  wire tmp5153;
  wire tmp5154;
  wire tmp5155;
  wire tmp5156;
  wire tmp5157;
  wire tmp5158;
  wire tmp5159;
  wire tmp5160;
  wire tmp5161;
  wire tmp5162;
  wire tmp5163;
  wire tmp5164;
  wire tmp5165;
  wire tmp5166;
  wire tmp5167;
  wire tmp5168;
  wire tmp5169;
  wire tmp5170;
  wire tmp5171;
  wire tmp5172;
  wire tmp5173;
  wire tmp5174;
  wire tmp5175;
  wire tmp5176;
  wire tmp5177;
  wire tmp5178;
  wire tmp5179;
  wire tmp5180;
  wire tmp5181;
  wire tmp5182;
  wire tmp5183;
  wire tmp5184;
  wire tmp5185;
  wire tmp5186;
  wire tmp5187;
  wire tmp5188;
  wire tmp5189;
  wire tmp5190;
  wire tmp5191;
  wire tmp5192;
  wire tmp5193;
  wire tmp5194;
  wire tmp5195;
  wire tmp5196;
  wire tmp5197;
  wire tmp5198;
  wire tmp5199;
  wire tmp5200;
  wire tmp5201;
  wire tmp5202;
  wire tmp5203;
  wire tmp5204;
  wire tmp5205;
  wire tmp5206;
  wire tmp5207;
  wire tmp5208;
  wire tmp5209;
  wire tmp5210;
  wire tmp5211;
  wire tmp5212;
  wire tmp5213;
  wire tmp5214;
  wire tmp5215;
  wire tmp5216;
  wire tmp5217;
  wire tmp5218;
  wire tmp5219;
  wire tmp5220;
  wire tmp5221;
  wire tmp5222;
  wire tmp5223;
  wire tmp5224;
  wire tmp5225;
  wire tmp5226;
  wire tmp5227;
  wire tmp5228;
  wire tmp5229;
  wire tmp5230;
  wire tmp5231;
  wire tmp5232;
  wire tmp5233;
  wire tmp5234;
  wire tmp5235;
  wire tmp5236;
  wire tmp5237;
  wire tmp5238;
  wire tmp5239;
  wire tmp5240;
  wire tmp5241;
  wire tmp5242;
  wire tmp5243;
  wire tmp5244;
  wire tmp5245;
  wire tmp5246;
  wire tmp5247;
  wire tmp5248;
  wire tmp5249;
  wire tmp5250;
  wire tmp5251;
  wire tmp5252;
  wire tmp5253;
  wire tmp5254;
  wire tmp5255;
  wire tmp5256;
  wire tmp5257;
  wire tmp5258;
  wire tmp5259;
  wire tmp5260;
  wire tmp5261;
  wire tmp5262;
  wire tmp5263;
  wire tmp5264;
  wire tmp5265;
  wire tmp5266;
  wire tmp5267;
  wire tmp5268;
  wire tmp5269;
  wire tmp5270;
  wire tmp5271;
  wire tmp5272;
  wire tmp5273;
  wire tmp5274;
  wire tmp5275;
  wire tmp5276;
  wire tmp5277;
  wire tmp5278;
  wire tmp5279;
  wire tmp5280;
  wire tmp5281;
  wire tmp5282;
  wire tmp5283;
  wire tmp5284;
  wire tmp5285;
  wire tmp5286;
  wire tmp5287;
  wire tmp5288;
  wire tmp5289;
  wire tmp5290;
  wire tmp5291;
  wire tmp5292;
  wire tmp5293;
  wire tmp5294;
  wire tmp5295;
  wire tmp5296;
  wire tmp5297;
  wire tmp5298;
  wire tmp5299;
  wire tmp5300;
  wire tmp5301;
  wire tmp5302;
  wire tmp5303;
  wire tmp5304;
  wire tmp5305;
  wire tmp5306;
  wire tmp5307;
  wire tmp5308;
  wire tmp5309;
  wire tmp5310;
  wire tmp5311;
  wire tmp5312;
  wire tmp5313;
  wire tmp5314;
  wire tmp5315;
  wire tmp5316;
  wire tmp5317;
  wire tmp5318;
  wire tmp5319;
  wire tmp5320;
  wire tmp5321;
  wire tmp5322;
  wire tmp5323;
  wire tmp5324;
  wire tmp5325;
  wire tmp5326;
  wire tmp5327;
  wire tmp5328;
  wire tmp5329;
  wire tmp5330;
  wire tmp5331;
  wire tmp5332;
  wire tmp5333;
  wire tmp5334;
  wire tmp5335;
  wire tmp5336;
  wire tmp5337;
  wire tmp5338;
  wire tmp5339;
  wire tmp5340;
  wire tmp5341;
  wire tmp5342;
  wire tmp5343;
  wire tmp5344;
  wire tmp5345;
  wire tmp5346;
  wire tmp5347;
  wire tmp5348;
  wire tmp5349;
  wire tmp5350;
  wire tmp5351;
  wire tmp5352;
  wire tmp5353;
  wire tmp5354;
  wire tmp5355;
  wire tmp5356;
  wire tmp5357;
  wire tmp5358;
  wire tmp5359;
  wire tmp5360;
  wire tmp5361;
  wire tmp5362;
  wire tmp5363;
  wire tmp5364;
  wire tmp5365;
  wire tmp5366;
  wire tmp5367;
  wire tmp5368;
  wire tmp5369;
  wire tmp5370;
  wire tmp5371;
  wire tmp5372;
  wire tmp5373;
  wire tmp5374;
  wire tmp5375;
  wire tmp5376;
  wire tmp5377;
  wire tmp5378;
  wire tmp5379;
  wire tmp5380;
  wire tmp5381;
  wire tmp5382;
  wire tmp5383;
  wire tmp5384;
  wire tmp5385;
  wire tmp5386;
  wire tmp5387;
  wire tmp5388;
  wire tmp5389;
  wire tmp5390;
  wire tmp5391;
  wire tmp5392;
  wire tmp5393;
  wire tmp5394;
  wire tmp5395;
  wire tmp5396;
  wire tmp5397;
  wire tmp5398;
  wire tmp5399;
  wire tmp5400;
  wire tmp5401;
  wire tmp5402;
  wire tmp5403;
  wire tmp5404;
  wire tmp5405;
  wire tmp5406;
  wire tmp5407;
  wire tmp5408;
  wire tmp5409;
  wire tmp5410;
  wire tmp5411;
  wire tmp5412;
  wire tmp5413;
  wire tmp5414;
  wire tmp5415;
  wire tmp5416;
  wire tmp5417;
  wire tmp5418;
  wire tmp5419;
  wire tmp5420;
  wire tmp5421;
  wire tmp5422;
  wire tmp5423;
  wire tmp5424;
  wire tmp5425;
  wire tmp5426;
  wire tmp5427;
  wire tmp5428;
  wire tmp5429;
  wire tmp5430;
  wire tmp5431;
  wire tmp5432;
  wire tmp5433;
  wire tmp5434;
  wire tmp5435;
  wire tmp5436;
  wire tmp5437;
  wire tmp5438;
  wire tmp5439;
  wire tmp5440;
  wire tmp5441;
  wire tmp5442;
  wire tmp5443;
  wire tmp5444;
  wire tmp5445;
  wire tmp5446;
  wire tmp5447;
  wire tmp5448;
  wire tmp5449;
  wire tmp5450;
  wire tmp5451;
  wire tmp5452;
  wire tmp5453;
  wire tmp5454;
  wire tmp5455;
  wire tmp5456;
  wire tmp5457;
  wire tmp5458;
  wire tmp5459;
  wire tmp5460;
  wire tmp5461;
  wire tmp5462;
  wire tmp5463;
  wire tmp5464;
  wire tmp5465;
  wire tmp5466;
  wire tmp5467;
  wire tmp5468;
  wire tmp5469;
  wire tmp5470;
  wire tmp5471;
  wire tmp5472;
  wire tmp5473;
  wire tmp5474;
  wire tmp5475;
  wire tmp5476;
  wire tmp5477;
  wire tmp5478;
  wire tmp5479;
  wire tmp5480;
  wire tmp5481;
  wire tmp5482;
  wire tmp5483;
  wire tmp5484;
  wire tmp5485;
  wire tmp5486;
  wire tmp5487;
  wire tmp5488;
  wire tmp5489;
  wire tmp5490;
  wire tmp5491;
  wire tmp5492;
  wire tmp5493;
  wire tmp5494;
  wire tmp5495;
  wire tmp5496;
  wire tmp5497;
  wire tmp5498;
  wire tmp5499;
  wire tmp5500;
  wire tmp5501;
  wire tmp5502;
  wire tmp5503;
  wire tmp5504;
  wire tmp5505;
  wire tmp5506;
  wire tmp5507;
  wire tmp5508;
  wire tmp5509;
  wire tmp5510;
  wire tmp5511;
  wire tmp5512;
  wire tmp5513;
  wire tmp5514;
  wire tmp5515;
  wire tmp5516;
  wire tmp5517;
  wire tmp5518;
  wire tmp5519;
  wire tmp5520;
  wire tmp5521;
  wire tmp5522;
  wire tmp5523;
  wire tmp5524;
  wire tmp5525;
  wire tmp5526;
  wire tmp5527;
  wire tmp5528;
  wire tmp5529;
  wire tmp5530;
  wire tmp5531;
  wire tmp5532;
  wire tmp5533;
  wire tmp5534;
  wire tmp5535;
  wire tmp5536;
  wire tmp5537;
  wire tmp5538;
  wire tmp5539;
  wire tmp5540;
  wire tmp5541;
  wire tmp5542;
  wire tmp5543;
  wire tmp5544;
  wire tmp5545;
  wire tmp5546;
  wire tmp5547;
  wire tmp5548;
  wire tmp5549;
  wire tmp5550;
  wire tmp5551;
  wire tmp5552;
  wire tmp5553;
  wire tmp5554;
  wire tmp5555;
  wire tmp5556;
  wire tmp5557;
  wire tmp5558;
  wire tmp5559;
  wire tmp5560;
  wire tmp5561;
  wire tmp5562;
  wire tmp5563;
  wire tmp5564;
  wire tmp5565;
  wire tmp5566;
  wire tmp5567;
  wire tmp5568;
  wire tmp5569;
  wire tmp5570;
  wire tmp5571;
  wire tmp5572;
  wire tmp5573;
  wire tmp5574;
  wire tmp5575;
  wire tmp5576;
  wire tmp5577;
  wire tmp5578;
  wire tmp5579;
  wire tmp5580;
  wire tmp5581;
  wire tmp5582;
  wire tmp5583;
  wire tmp5584;
  wire tmp5585;
  wire tmp5586;
  wire tmp5587;
  wire tmp5588;
  wire tmp5589;
  wire tmp5590;
  wire tmp5591;
  wire tmp5592;
  wire tmp5593;
  wire tmp5594;
  wire tmp5595;
  wire tmp5596;
  wire tmp5597;
  wire tmp5598;
  wire tmp5599;
  wire tmp5600;
  wire tmp5601;
  wire tmp5602;
  wire tmp5603;
  wire tmp5604;
  wire tmp5605;
  wire tmp5606;
  wire tmp5607;
  wire tmp5608;
  wire tmp5609;
  wire tmp5610;
  wire tmp5611;
  wire tmp5612;
  wire tmp5613;
  wire tmp5614;
  wire tmp5615;
  wire tmp5616;
  wire tmp5617;
  wire tmp5618;
  wire tmp5619;
  wire tmp5620;
  wire tmp5621;
  wire tmp5622;
  wire tmp5623;
  wire tmp5624;
  wire tmp5625;
  wire tmp5626;
  wire tmp5627;
  wire tmp5628;
  wire tmp5629;
  wire tmp5630;
  wire tmp5631;
  wire tmp5632;
  wire tmp5633;
  wire tmp5634;
  wire tmp5635;
  wire tmp5636;
  wire tmp5637;
  wire tmp5638;
  wire tmp5639;
  wire tmp5640;
  wire tmp5641;
  wire tmp5642;
  wire tmp5643;
  wire tmp5644;
  wire tmp5645;
  wire tmp5646;
  wire tmp5647;
  wire tmp5648;
  wire tmp5649;
  wire tmp5650;
  wire tmp5651;
  wire tmp5652;
  wire tmp5653;
  wire tmp5654;
  wire tmp5655;
  wire tmp5656;
  wire tmp5657;
  wire tmp5658;
  wire tmp5659;
  wire tmp5660;
  wire tmp5661;
  wire tmp5662;
  wire tmp5663;
  wire tmp5664;
  wire tmp5665;
  wire tmp5666;
  wire tmp5667;
  wire tmp5668;
  wire tmp5669;
  wire tmp5670;
  wire tmp5671;
  wire tmp5672;
  wire tmp5673;
  wire tmp5674;
  wire tmp5675;
  wire tmp5676;
  wire tmp5677;
  wire tmp5678;
  wire tmp5679;
  wire tmp5680;
  wire tmp5681;
  wire tmp5682;
  wire tmp5683;
  wire tmp5684;
  wire tmp5685;
  wire tmp5686;
  wire tmp5687;
  wire tmp5688;
  wire tmp5689;
  wire tmp5690;
  wire tmp5691;
  wire tmp5692;
  wire tmp5693;
  wire tmp5694;
  wire tmp5695;
  wire tmp5696;
  wire tmp5697;
  wire tmp5698;
  wire tmp5699;
  wire tmp5700;
  wire tmp5701;
  wire tmp5702;
  wire tmp5703;
  wire tmp5704;
  wire tmp5705;
  wire tmp5706;
  wire tmp5707;
  wire tmp5708;
  wire tmp5709;
  wire tmp5710;
  wire tmp5711;
  wire tmp5712;
  wire tmp5713;
  wire tmp5714;
  wire tmp5715;
  wire tmp5716;
  wire tmp5717;
  wire tmp5718;
  wire tmp5719;
  wire tmp5720;
  wire tmp5721;
  wire tmp5722;
  wire tmp5723;
  wire tmp5724;
  wire tmp5725;
  wire tmp5726;
  wire tmp5727;
  wire tmp5728;
  wire tmp5729;
  wire tmp5730;
  wire tmp5731;
  wire tmp5732;
  wire tmp5733;
  wire tmp5734;
  wire tmp5735;
  wire tmp5736;
  wire tmp5737;
  wire tmp5738;
  wire tmp5739;
  wire tmp5740;
  wire tmp5741;
  wire tmp5742;
  wire tmp5743;
  wire tmp5744;
  wire tmp5745;
  wire tmp5746;
  wire tmp5747;
  wire tmp5748;
  wire tmp5749;
  wire tmp5750;
  wire tmp5751;
  wire tmp5752;
  wire tmp5753;
  wire tmp5754;
  wire tmp5755;
  wire tmp5756;
  wire tmp5757;
  wire tmp5758;
  wire tmp5759;
  wire tmp5760;
  wire tmp5761;
  wire tmp5762;
  wire tmp5763;
  wire tmp5764;
  wire tmp5765;
  wire tmp5766;
  wire tmp5767;
  wire tmp5768;
  wire tmp5769;
  wire tmp5770;
  wire tmp5771;
  wire tmp5772;
  wire tmp5773;
  wire tmp5774;
  wire tmp5775;
  wire tmp5776;
  wire tmp5777;
  wire tmp5778;
  wire tmp5779;
  wire tmp5780;
  wire tmp5781;
  wire tmp5782;
  wire tmp5783;
  wire tmp5784;
  wire tmp5785;
  wire tmp5786;
  wire tmp5787;
  wire tmp5788;
  wire tmp5789;
  wire tmp5790;
  wire tmp5791;
  wire tmp5792;
  wire tmp5793;
  wire tmp5794;
  wire tmp5795;
  wire tmp5796;
  wire tmp5797;
  wire tmp5798;
  wire tmp5799;
  wire tmp5800;
  wire tmp5801;
  wire tmp5802;
  wire tmp5803;
  wire tmp5804;
  wire tmp5805;
  wire tmp5806;
  wire tmp5807;
  wire tmp5808;
  wire tmp5809;
  wire tmp5810;
  wire tmp5811;
  wire tmp5812;
  wire tmp5813;
  wire tmp5814;
  wire tmp5815;
  wire tmp5816;
  wire tmp5817;
  wire tmp5818;
  wire tmp5819;
  wire tmp5820;
  wire tmp5821;
  wire tmp5822;
  wire tmp5823;
  wire tmp5824;
  wire tmp5825;
  wire tmp5826;
  wire tmp5827;
  wire tmp5828;
  wire tmp5829;
  wire tmp5830;
  wire tmp5831;
  wire tmp5832;
  wire tmp5833;
  wire tmp5834;
  wire tmp5835;
  wire tmp5836;
  wire tmp5837;
  wire tmp5838;
  wire tmp5839;
  wire tmp5840;
  wire tmp5841;
  wire tmp5842;
  wire tmp5843;
  wire tmp5844;
  wire tmp5845;
  wire tmp5846;
  wire tmp5847;
  wire tmp5848;
  wire tmp5849;
  wire tmp5850;
  wire tmp5851;
  wire tmp5852;
  wire tmp5853;
  wire tmp5854;
  wire tmp5855;
  wire tmp5856;
  wire tmp5857;
  wire tmp5858;
  wire tmp5859;
  wire tmp5860;
  wire tmp5861;
  wire tmp5862;
  wire tmp5863;
  wire tmp5864;
  wire tmp5865;
  wire tmp5866;
  wire tmp5867;
  wire tmp5868;
  wire tmp5869;
  wire tmp5870;
  wire tmp5871;
  wire tmp5872;
  wire tmp5873;
  wire tmp5874;
  wire tmp5875;
  wire tmp5876;
  wire tmp5877;
  wire tmp5878;
  wire tmp5879;
  wire tmp5880;
  wire tmp5881;
  wire tmp5882;
  wire tmp5883;
  wire tmp5884;
  wire tmp5885;
  wire tmp5886;
  wire tmp5887;
  wire tmp5888;
  wire tmp5889;
  wire tmp5890;
  wire tmp5891;
  wire tmp5892;
  wire tmp5893;
  wire tmp5894;
  wire tmp5895;
  wire tmp5896;
  wire tmp5897;
  wire tmp5898;
  wire tmp5899;
  wire tmp5900;
  wire tmp5901;
  wire tmp5902;
  wire tmp5903;
  wire tmp5904;
  wire tmp5905;
  wire tmp5906;
  wire tmp5907;
  wire tmp5908;
  wire tmp5909;
  wire tmp5910;
  wire tmp5911;
  wire tmp5912;
  wire tmp5913;
  wire tmp5914;
  wire tmp5915;
  wire tmp5916;
  wire tmp5917;
  wire tmp5918;
  wire tmp5919;
  wire tmp5920;
  wire tmp5921;
  wire tmp5922;
  wire tmp5923;
  wire tmp5924;
  wire tmp5925;
  wire tmp5926;
  wire tmp5927;
  wire tmp5928;
  wire tmp5929;
  wire tmp5930;
  wire tmp5931;
  wire tmp5932;
  wire tmp5933;
  wire tmp5934;
  wire tmp5935;
  wire tmp5936;
  wire tmp5937;
  wire tmp5938;
  wire tmp5939;
  wire tmp5940;
  wire tmp5941;
  wire tmp5942;
  wire tmp5943;
  wire tmp5944;
  wire tmp5945;
  wire tmp5946;
  wire tmp5947;
  wire tmp5948;
  wire tmp5949;
  wire tmp5950;
  wire tmp5951;
  wire tmp5952;
  wire tmp5953;
  wire tmp5954;
  wire tmp5955;
  wire tmp5956;
  wire tmp5957;
  wire tmp5958;
  wire tmp5959;
  wire tmp5960;
  wire tmp5961;
  wire tmp5962;
  wire tmp5963;
  wire tmp5964;
  wire tmp5965;
  wire tmp5966;
  wire tmp5967;
  wire tmp5968;
  wire tmp5969;
  wire tmp5970;
  wire tmp5971;
  wire tmp5972;
  wire tmp5973;
  wire tmp5974;
  wire tmp5975;
  wire tmp5976;
  wire tmp5977;
  wire tmp5978;
  wire tmp5979;
  wire tmp5980;
  wire tmp5981;
  wire tmp5982;
  wire tmp5983;
  wire tmp5984;
  wire tmp5985;
  wire tmp5986;
  wire tmp5987;
  wire tmp5988;
  wire tmp5989;
  wire tmp5990;
  wire tmp5991;
  wire tmp5992;
  wire tmp5993;
  wire tmp5994;
  wire tmp5995;
  wire tmp5996;
  wire tmp5997;
  wire tmp5998;
  wire tmp5999;
  wire tmp6000;
  wire tmp6001;
  wire tmp6002;
  wire tmp6003;
  wire tmp6004;
  wire tmp6005;
  wire tmp6006;
  wire tmp6007;
  wire tmp6008;
  wire tmp6009;
  wire tmp6010;
  wire tmp6011;
  wire tmp6012;
  wire tmp6013;
  wire tmp6014;
  wire tmp6015;
  wire tmp6016;
  wire tmp6017;
  wire tmp6018;
  wire tmp6019;
  wire tmp6020;
  wire tmp6021;
  wire tmp6022;
  wire tmp6023;
  wire tmp6024;
  wire tmp6025;
  wire tmp6026;
  wire tmp6027;
  wire tmp6028;
  wire tmp6029;
  wire tmp6030;
  wire tmp6031;
  wire tmp6032;
  wire tmp6033;
  wire tmp6034;
  wire tmp6035;
  wire tmp6036;
  wire tmp6037;
  wire tmp6038;
  wire tmp6039;
  wire tmp6040;
  wire tmp6041;
  wire tmp6042;
  wire tmp6043;
  wire tmp6044;
  wire tmp6045;
  wire tmp6046;
  wire tmp6047;
  wire tmp6048;
  wire tmp6049;
  wire tmp6050;
  wire tmp6051;
  wire tmp6052;
  wire tmp6053;
  wire tmp6054;
  wire tmp6055;
  wire tmp6056;
  wire tmp6057;
  wire tmp6058;
  wire tmp6059;
  wire tmp6060;
  wire tmp6061;
  wire tmp6062;
  wire tmp6063;
  wire tmp6064;
  wire tmp6065;
  wire tmp6066;
  wire tmp6067;
  wire tmp6068;
  wire tmp6069;
  wire tmp6070;
  wire tmp6071;
  wire tmp6072;
  wire tmp6073;
  wire tmp6074;
  wire tmp6075;
  wire tmp6076;
  wire tmp6077;
  wire tmp6078;
  wire tmp6079;
  wire tmp6080;
  wire tmp6081;
  wire tmp6082;
  wire tmp6083;
  wire tmp6084;
  wire tmp6085;
  wire tmp6086;
  wire tmp6087;
  wire tmp6088;
  wire tmp6089;
  wire tmp6090;
  wire tmp6091;
  wire tmp6092;
  wire tmp6093;
  wire tmp6094;
  wire tmp6095;
  wire tmp6096;
  wire tmp6097;
  wire tmp6098;
  wire tmp6099;
  wire tmp6100;
  wire tmp6101;
  wire tmp6102;
  wire tmp6103;
  wire tmp6104;
  wire tmp6105;
  wire tmp6106;
  wire tmp6107;
  wire tmp6108;
  wire tmp6109;
  wire tmp6110;
  wire tmp6111;
  wire tmp6112;
  wire tmp6113;
  wire tmp6114;
  wire tmp6115;
  wire tmp6116;
  wire tmp6117;
  wire tmp6118;
  wire tmp6119;
  wire tmp6120;
  wire tmp6121;
  wire tmp6122;
  wire tmp6123;
  wire tmp6124;
  wire tmp6125;
  wire tmp6126;
  wire tmp6127;
  wire tmp6128;
  wire tmp6129;
  wire tmp6130;
  wire tmp6131;
  wire tmp6132;
  wire tmp6133;
  wire tmp6134;
  wire tmp6135;
  wire tmp6136;
  wire tmp6137;
  wire tmp6138;
  wire tmp6139;
  wire tmp6140;
  wire tmp6141;
  wire tmp6142;
  wire tmp6143;
  wire tmp6144;
  wire tmp6145;
  wire tmp6146;
  wire tmp6147;
  wire tmp6148;
  wire tmp6149;
  wire tmp6150;
  wire tmp6151;
  wire tmp6152;
  wire tmp6153;
  wire tmp6154;
  wire tmp6155;
  wire tmp6156;
  wire tmp6157;
  wire tmp6158;
  wire tmp6159;
  wire tmp6160;
  wire tmp6161;
  wire tmp6162;
  wire tmp6163;
  wire tmp6164;
  wire tmp6165;
  wire tmp6166;
  wire tmp6167;
  wire tmp6168;
  wire tmp6169;
  wire tmp6170;
  wire tmp6171;
  wire tmp6172;
  wire tmp6173;
  wire tmp6174;
  wire tmp6175;
  wire tmp6176;
  wire tmp6177;
  wire tmp6178;
  wire tmp6179;
  wire tmp6180;
  wire tmp6181;
  wire tmp6182;
  wire tmp6183;
  wire tmp6184;
  wire tmp6185;
  wire tmp6186;
  wire tmp6187;
  wire tmp6188;
  wire tmp6189;
  wire tmp6190;
  wire tmp6191;
  wire tmp6192;
  wire tmp6193;
  wire tmp6194;
  wire tmp6195;
  wire tmp6196;
  wire tmp6197;
  wire tmp6198;
  wire tmp6199;
  wire tmp6200;
  wire tmp6201;
  wire tmp6202;
  wire tmp6203;
  wire tmp6204;
  wire tmp6205;
  wire tmp6206;
  wire tmp6207;
  wire tmp6208;
  wire tmp6209;
  wire tmp6210;
  wire tmp6211;
  wire tmp6212;
  wire tmp6213;
  wire tmp6214;
  wire tmp6215;
  wire tmp6216;
  wire tmp6217;
  wire tmp6218;
  wire tmp6219;
  wire tmp6220;
  wire tmp6221;
  wire tmp6222;
  wire tmp6223;
  wire tmp6224;
  wire tmp6225;
  wire tmp6226;
  wire tmp6227;
  wire tmp6228;
  wire tmp6229;
  wire tmp6230;
  wire tmp6231;
  wire tmp6232;
  wire tmp6233;
  wire tmp6234;
  wire tmp6235;
  wire tmp6236;
  wire tmp6237;
  wire tmp6238;
  wire tmp6239;
  wire tmp6240;
  wire tmp6241;
  wire tmp6242;
  wire tmp6243;
  wire tmp6244;
  wire tmp6245;
  wire tmp6246;
  wire tmp6247;
  wire tmp6248;
  wire tmp6249;
  wire tmp6250;
  wire tmp6251;
  wire tmp6252;
  wire tmp6253;
  wire tmp6254;
  wire tmp6255;
  wire tmp6256;
  wire tmp6257;
  wire tmp6258;
  wire tmp6259;
  wire tmp6260;
  wire tmp6261;
  wire tmp6262;
  wire tmp6263;
  wire tmp6264;
  wire tmp6265;
  wire tmp6266;
  wire tmp6267;
  wire tmp6268;
  wire tmp6269;
  wire tmp6270;
  wire tmp6271;
  wire tmp6272;
  wire tmp6273;
  wire tmp6274;
  wire tmp6275;
  wire tmp6276;
  wire tmp6277;
  wire tmp6278;
  wire tmp6279;
  wire tmp6280;
  wire tmp6281;
  wire tmp6282;
  wire tmp6283;
  wire tmp6284;
  wire tmp6285;
  wire tmp6286;
  wire tmp6287;
  wire tmp6288;
  wire tmp6289;
  wire tmp6290;
  wire tmp6291;
  wire tmp6292;
  wire tmp6293;
  wire tmp6294;
  wire tmp6295;
  wire tmp6296;
  wire tmp6297;
  wire tmp6298;
  wire tmp6299;
  wire tmp6300;
  wire tmp6301;
  wire tmp6302;
  wire tmp6303;
  wire tmp6304;
  wire tmp6305;
  wire tmp6306;
  wire tmp6307;
  wire tmp6308;
  wire tmp6309;
  wire tmp6310;
  wire tmp6311;
  wire tmp6312;
  wire tmp6313;
  wire tmp6314;
  wire tmp6315;
  wire tmp6316;
  wire tmp6317;
  wire tmp6318;
  wire tmp6319;
  wire tmp6320;
  wire tmp6321;
  wire tmp6322;
  wire tmp6323;
  wire tmp6324;
  wire tmp6325;
  wire tmp6326;
  wire tmp6327;
  wire tmp6328;
  wire tmp6329;
  wire tmp6330;
  wire tmp6331;
  wire tmp6332;
  wire tmp6333;
  wire tmp6334;
  wire tmp6335;
  wire tmp6336;
  wire tmp6337;
  wire tmp6338;
  wire tmp6339;
  wire tmp6340;
  wire tmp6341;
  wire tmp6342;
  wire tmp6343;
  wire tmp6344;
  wire tmp6345;
  wire tmp6346;
  wire tmp6347;
  wire tmp6348;
  wire tmp6349;
  wire tmp6350;
  wire tmp6351;
  wire tmp6352;
  wire tmp6353;
  wire tmp6354;
  wire tmp6355;
  wire tmp6356;
  wire tmp6357;
  wire tmp6358;
  wire tmp6359;
  wire tmp6360;
  wire tmp6361;
  wire tmp6362;
  wire tmp6363;
  wire tmp6364;
  wire tmp6365;
  wire tmp6366;
  wire tmp6367;
  wire tmp6368;
  wire tmp6369;
  wire tmp6370;
  wire tmp6371;
  wire tmp6372;
  wire tmp6373;
  wire tmp6374;
  wire tmp6375;
  wire tmp6376;
  wire tmp6377;
  wire tmp6378;
  wire tmp6379;
  wire tmp6380;
  wire tmp6381;
  wire tmp6382;
  wire tmp6383;
  wire tmp6384;
  wire tmp6385;
  wire tmp6386;
  wire tmp6387;
  wire tmp6388;
  wire tmp6389;
  wire tmp6390;
  wire tmp6391;
  wire tmp6392;
  wire tmp6393;
  wire tmp6394;
  wire tmp6395;
  wire tmp6396;
  wire tmp6397;
  wire tmp6398;
  wire tmp6399;
  wire tmp6400;
  wire tmp6401;
  wire tmp6402;
  wire tmp6403;
  wire tmp6404;
  wire tmp6405;
  wire tmp6406;
  wire tmp6407;
  wire tmp6408;
  wire tmp6409;
  wire tmp6410;
  wire tmp6411;
  wire tmp6412;
  wire tmp6413;
  wire tmp6414;
  wire tmp6415;
  wire tmp6416;
  wire tmp6417;
  wire tmp6418;
  wire tmp6419;
  wire tmp6420;
  wire tmp6421;
  wire tmp6422;
  wire tmp6423;
  wire tmp6424;
  wire tmp6425;
  wire tmp6426;
  wire tmp6427;
  wire tmp6428;
  wire tmp6429;
  wire tmp6430;
  wire tmp6431;
  wire tmp6432;
  wire tmp6433;
  wire tmp6434;
  wire tmp6435;
  wire tmp6436;
  wire tmp6437;
  wire tmp6438;
  wire tmp6439;
  wire tmp6440;
  wire tmp6441;
  wire tmp6442;
  wire tmp6443;
  wire tmp6444;
  wire tmp6445;
  wire tmp6446;
  wire tmp6447;
  wire tmp6448;
  wire tmp6449;
  wire tmp6450;
  wire tmp6451;
  wire tmp6452;
  wire tmp6453;
  wire tmp6454;
  wire tmp6455;
  wire tmp6456;
  wire tmp6457;
  wire tmp6458;
  wire tmp6459;
  wire tmp6460;
  wire tmp6461;
  wire tmp6462;
  wire tmp6463;
  wire tmp6464;
  wire tmp6465;
  wire tmp6466;
  wire tmp6467;
  wire tmp6468;
  wire tmp6469;
  wire tmp6470;
  wire tmp6471;
  wire tmp6472;
  wire tmp6473;
  wire tmp6474;
  wire tmp6475;
  wire tmp6476;
  wire tmp6477;
  wire tmp6478;
  wire tmp6479;
  wire tmp6480;
  wire tmp6481;
  wire tmp6482;
  wire tmp6483;
  wire tmp6484;
  wire tmp6485;
  wire tmp6486;
  wire tmp6487;
  wire tmp6488;
  wire tmp6489;
  wire tmp6490;
  wire tmp6491;
  wire tmp6492;
  wire tmp6493;
  wire tmp6494;
  wire tmp6495;
  wire tmp6496;
  wire tmp6497;
  wire tmp6498;
  wire tmp6499;
  wire tmp6500;
  wire tmp6501;
  wire tmp6502;
  wire tmp6503;
  wire tmp6504;
  wire tmp6505;
  wire tmp6506;
  wire tmp6507;
  wire tmp6508;
  wire tmp6509;
  wire tmp6510;
  wire tmp6511;
  wire tmp6512;
  wire tmp6513;
  wire tmp6514;
  wire tmp6515;
  wire tmp6516;
  wire tmp6517;
  wire tmp6518;
  wire tmp6519;
  wire tmp6520;
  wire tmp6521;
  wire tmp6522;
  wire tmp6523;
  wire tmp6524;
  wire tmp6525;
  wire tmp6526;
  wire tmp6527;
  wire tmp6528;
  wire tmp6529;
  wire tmp6530;
  wire tmp6531;
  wire tmp6532;
  wire tmp6533;
  wire tmp6534;
  wire tmp6535;
  wire tmp6536;
  wire tmp6537;
  wire tmp6538;
  wire tmp6539;
  wire tmp6540;
  wire tmp6541;
  wire tmp6542;
  wire tmp6543;
  wire tmp6544;
  wire tmp6545;
  wire tmp6546;
  wire tmp6547;
  wire tmp6548;
  wire tmp6549;
  wire tmp6550;
  wire tmp6551;
  wire tmp6552;
  wire tmp6553;
  wire tmp6554;
  wire tmp6555;
  wire tmp6556;
  wire tmp6557;
  wire tmp6558;
  wire tmp6559;
  wire tmp6560;
  wire tmp6561;
  wire tmp6562;
  wire tmp6563;
  wire tmp6564;
  wire tmp6565;
  wire tmp6566;
  wire tmp6567;
  wire tmp6568;
  wire tmp6569;
  wire tmp6570;
  wire tmp6571;
  wire tmp6572;
  wire tmp6573;
  wire tmp6574;
  wire tmp6575;
  wire tmp6576;
  wire tmp6577;
  wire tmp6578;
  wire tmp6579;
  wire tmp6580;
  wire tmp6581;
  wire tmp6582;
  wire tmp6583;
  wire tmp6584;
  wire tmp6585;
  wire tmp6586;
  wire tmp6587;
  wire tmp6588;
  wire tmp6589;
  wire tmp6590;
  wire tmp6591;
  wire tmp6592;
  wire tmp6593;
  wire tmp6594;
  wire tmp6595;
  wire tmp6596;
  wire tmp6597;
  wire tmp6598;
  wire tmp6599;
  wire tmp6600;
  wire tmp6601;
  wire tmp6602;
  wire tmp6603;
  wire tmp6604;
  wire tmp6605;
  wire tmp6606;
  wire tmp6607;
  wire tmp6608;
  wire tmp6609;
  wire tmp6610;
  wire tmp6611;
  wire tmp6612;
  wire tmp6613;
  wire tmp6614;
  wire tmp6615;
  wire tmp6616;
  wire tmp6617;
  wire tmp6618;
  wire tmp6619;
  wire tmp6620;
  wire tmp6621;
  wire tmp6622;
  wire tmp6623;
  wire tmp6624;
  wire tmp6625;
  wire tmp6626;
  wire tmp6627;
  wire tmp6628;
  wire tmp6629;
  wire tmp6630;
  wire tmp6631;
  wire tmp6632;
  wire tmp6633;
  wire tmp6634;
  wire tmp6635;
  wire tmp6636;
  wire tmp6637;
  wire tmp6638;
  wire tmp6639;
  wire tmp6640;
  wire tmp6641;
  wire tmp6642;
  wire tmp6643;
  wire tmp6644;
  wire tmp6645;
  wire tmp6646;
  wire tmp6647;
  wire tmp6648;
  wire tmp6649;
  wire tmp6650;
  wire tmp6651;
  wire tmp6652;
  wire tmp6653;
  wire tmp6654;
  wire tmp6655;
  wire tmp6656;
  wire tmp6657;
  wire tmp6658;
  wire tmp6659;
  wire tmp6660;
  wire tmp6661;
  wire tmp6662;
  wire tmp6663;
  wire tmp6664;
  wire tmp6665;
  wire tmp6666;
  wire tmp6667;
  wire tmp6668;
  wire tmp6669;
  wire tmp6670;
  wire tmp6671;
  wire tmp6672;
  wire tmp6673;
  wire tmp6674;
  wire tmp6675;
  wire tmp6676;
  wire tmp6677;
  wire tmp6678;
  wire tmp6679;
  wire tmp6680;
  wire tmp6681;
  wire tmp6682;
  wire tmp6683;
  wire tmp6684;
  wire tmp6685;
  wire tmp6686;
  wire tmp6687;
  wire tmp6688;
  wire tmp6689;
  wire tmp6690;
  wire tmp6691;
  wire tmp6692;
  wire tmp6693;
  wire tmp6694;
  wire tmp6695;
  wire tmp6696;
  wire tmp6697;
  wire tmp6698;
  wire tmp6699;
  wire tmp6700;
  wire tmp6701;
  wire tmp6702;
  wire tmp6703;
  wire tmp6704;
  wire tmp6705;
  wire tmp6706;
  wire tmp6707;
  wire tmp6708;
  wire tmp6709;
  wire tmp6710;
  wire tmp6711;
  wire tmp6712;
  wire tmp6713;
  wire tmp6714;
  wire tmp6715;
  wire tmp6716;
  wire tmp6717;
  wire tmp6718;
  wire tmp6719;
  wire tmp6720;
  wire tmp6721;
  wire tmp6722;
  wire tmp6723;
  wire tmp6724;
  wire tmp6725;
  wire tmp6726;
  wire tmp6727;
  wire tmp6728;
  wire tmp6729;
  wire tmp6730;
  wire tmp6731;
  wire tmp6732;
  wire tmp6733;
  wire tmp6734;
  wire tmp6735;
  wire tmp6736;
  wire tmp6737;
  wire tmp6738;
  wire tmp6739;
  wire tmp6740;
  wire tmp6741;
  wire tmp6742;
  wire tmp6743;
  wire tmp6744;
  wire tmp6745;
  wire tmp6746;
  wire tmp6747;
  wire tmp6748;
  wire tmp6749;
  wire tmp6750;
  wire tmp6751;
  wire tmp6752;
  wire tmp6753;
  wire tmp6754;
  wire tmp6755;
  wire tmp6756;
  wire tmp6757;
  wire tmp6758;
  wire tmp6759;
  wire tmp6760;
  wire tmp6761;
  wire tmp6762;
  wire tmp6763;
  wire tmp6764;
  wire tmp6765;
  wire tmp6766;
  wire tmp6767;
  wire tmp6768;
  wire tmp6769;
  wire tmp6770;
  wire tmp6771;
  wire tmp6772;
  wire tmp6773;
  wire tmp6774;
  wire tmp6775;
  wire tmp6776;
  wire tmp6777;
  wire tmp6778;
  wire tmp6779;
  wire tmp6780;
  wire tmp6781;
  wire tmp6782;
  wire tmp6783;
  wire tmp6784;
  wire tmp6785;
  wire tmp6786;
  wire tmp6787;
  wire tmp6788;
  wire tmp6789;
  wire tmp6790;
  wire tmp6791;
  wire tmp6792;
  wire tmp6793;
  wire tmp6794;
  wire tmp6795;
  wire tmp6796;
  wire tmp6797;
  wire tmp6798;
  wire tmp6799;
  wire tmp6800;
  wire tmp6801;
  wire tmp6802;
  wire tmp6803;
  wire tmp6804;
  wire tmp6805;
  wire tmp6806;
  wire tmp6807;
  wire tmp6808;
  wire tmp6809;
  wire tmp6810;
  wire tmp6811;
  wire tmp6812;
  wire tmp6813;
  wire tmp6814;
  wire tmp6815;
  wire tmp6816;
  wire tmp6817;
  wire tmp6818;
  wire tmp6819;
  wire tmp6820;
  wire tmp6821;
  wire tmp6822;
  wire tmp6823;
  wire tmp6824;
  wire tmp6825;
  wire tmp6826;
  wire tmp6827;
  wire tmp6828;
  wire tmp6829;
  wire tmp6830;
  wire tmp6831;
  wire tmp6832;
  wire tmp6833;
  wire tmp6834;
  wire tmp6835;
  wire tmp6836;
  wire tmp6837;
  wire tmp6838;
  wire tmp6839;
  wire tmp6840;
  wire tmp6841;
  wire tmp6842;
  wire tmp6843;
  wire tmp6844;
  wire tmp6845;
  wire tmp6846;
  wire tmp6847;
  wire tmp6848;
  wire tmp6849;
  wire tmp6850;
  wire tmp6851;
  wire tmp6852;
  wire tmp6853;
  wire tmp6854;
  wire tmp6855;
  wire tmp6856;
  wire tmp6857;
  wire tmp6858;
  wire tmp6859;
  wire tmp6860;
  wire tmp6861;
  wire tmp6862;
  wire tmp6863;
  wire tmp6864;
  wire tmp6865;
  wire tmp6866;
  wire tmp6867;
  wire tmp6868;
  wire tmp6869;
  wire tmp6870;
  wire tmp6871;
  wire tmp6872;
  wire tmp6873;
  wire tmp6874;
  wire tmp6875;
  wire tmp6876;
  wire tmp6877;
  wire tmp6878;
  wire tmp6879;
  wire tmp6880;
  wire tmp6881;
  wire tmp6882;
  wire tmp6883;
  wire tmp6884;
  wire tmp6885;
  wire tmp6886;
  wire tmp6887;
  wire tmp6888;
  wire tmp6889;
  wire tmp6890;
  wire tmp6891;
  wire tmp6892;
  wire tmp6893;
  wire tmp6894;
  wire tmp6895;
  wire tmp6896;
  wire tmp6897;
  wire tmp6898;
  wire tmp6899;
  wire tmp6900;
  wire tmp6901;
  wire tmp6902;
  wire tmp6903;
  wire tmp6904;
  wire tmp6905;
  wire tmp6906;
  wire tmp6907;
  wire tmp6908;
  wire tmp6909;
  wire tmp6910;
  wire tmp6911;
  wire tmp6912;
  wire tmp6913;
  wire tmp6914;
  wire tmp6915;
  wire tmp6916;
  wire tmp6917;
  wire tmp6918;
  wire tmp6919;
  wire tmp6920;
  wire tmp6921;
  wire tmp6922;
  wire tmp6923;
  wire tmp6924;
  wire tmp6925;
  wire tmp6926;
  wire tmp6927;
  wire tmp6928;
  wire tmp6929;
  wire tmp6930;
  wire tmp6931;
  wire tmp6932;
  wire tmp6933;
  wire tmp6934;
  wire tmp6935;
  wire tmp6936;
  wire tmp6937;
  wire tmp6938;
  wire tmp6939;
  wire tmp6940;
  wire tmp6941;
  wire tmp6942;
  wire tmp6943;
  wire tmp6944;
  wire tmp6945;
  wire tmp6946;
  wire tmp6947;
  wire tmp6948;
  wire tmp6949;
  wire tmp6950;
  wire tmp6951;
  wire tmp6952;
  wire tmp6953;
  wire tmp6954;
  wire tmp6955;
  wire tmp6956;
  wire tmp6957;
  wire tmp6958;
  wire tmp6959;
  wire tmp6960;
  wire tmp6961;
  wire tmp6962;
  wire tmp6963;
  wire tmp6964;
  wire tmp6965;
  wire tmp6966;
  wire tmp6967;
  wire tmp6968;
  wire tmp6969;
  wire tmp6970;
  wire tmp6971;
  wire tmp6972;
  wire tmp6973;
  wire tmp6974;
  wire tmp6975;
  wire tmp6976;
  wire tmp6977;
  wire tmp6978;
  wire tmp6979;
  wire tmp6980;
  wire tmp6981;
  wire tmp6982;
  wire tmp6983;
  wire tmp6984;
  wire tmp6985;
  wire tmp6986;
  wire tmp6987;
  wire tmp6988;
  wire tmp6989;
  wire tmp6990;
  wire tmp6991;
  wire tmp6992;
  wire tmp6993;
  wire tmp6994;
  wire tmp6995;
  wire tmp6996;
  wire tmp6997;
  wire tmp6998;
  wire tmp6999;
  wire tmp7000;
  wire tmp7001;
  wire tmp7002;
  wire tmp7003;
  wire tmp7004;
  wire tmp7005;
  wire tmp7006;
  wire tmp7007;
  wire tmp7008;
  wire tmp7009;
  wire tmp7010;
  wire tmp7011;
  wire tmp7012;
  wire tmp7013;
  wire tmp7014;
  wire tmp7015;
  wire tmp7016;
  wire tmp7017;
  wire tmp7018;
  wire tmp7019;
  wire tmp7020;
  wire tmp7021;
  wire tmp7022;
  wire tmp7023;
  wire tmp7024;
  wire tmp7025;
  wire tmp7026;
  wire tmp7027;
  wire tmp7028;
  wire tmp7029;
  wire tmp7030;
  wire tmp7031;
  wire tmp7032;
  wire tmp7033;
  wire tmp7034;
  wire tmp7035;
  wire tmp7036;
  wire tmp7037;
  wire tmp7038;
  wire tmp7039;
  wire tmp7040;
  wire tmp7041;
  wire tmp7042;
  wire tmp7043;
  wire tmp7044;
  wire tmp7045;
  wire tmp7046;
  wire tmp7047;
  wire tmp7048;
  wire tmp7049;
  wire tmp7050;
  wire tmp7051;
  wire tmp7052;
  wire tmp7053;
  wire tmp7054;
  wire tmp7055;
  wire tmp7056;
  wire tmp7057;
  wire tmp7058;
  wire tmp7059;
  wire tmp7060;
  wire tmp7061;
  wire tmp7062;
  wire tmp7063;
  wire tmp7064;
  wire tmp7065;
  wire tmp7066;
  wire tmp7067;
  wire tmp7068;
  wire tmp7069;
  wire tmp7070;
  wire tmp7071;
  wire tmp7072;
  wire tmp7073;
  wire tmp7074;
  wire tmp7075;
  wire tmp7076;
  wire tmp7077;
  wire tmp7078;
  wire tmp7079;
  wire tmp7080;
  wire tmp7081;
  wire tmp7082;
  wire tmp7083;
  wire tmp7084;
  wire tmp7085;
  wire tmp7086;
  wire tmp7087;
  wire tmp7088;
  wire tmp7089;
  wire tmp7090;
  wire tmp7091;
  wire tmp7092;
  wire tmp7093;
  wire tmp7094;
  wire tmp7095;
  wire tmp7096;
  wire tmp7097;
  wire tmp7098;
  wire tmp7099;
  wire tmp7100;
  wire tmp7101;
  wire tmp7102;
  wire tmp7103;
  wire tmp7104;
  wire tmp7105;
  wire tmp7106;
  wire tmp7107;
  wire tmp7108;
  wire tmp7109;
  wire tmp7110;
  wire tmp7111;
  wire tmp7112;
  wire tmp7113;
  wire tmp7114;
  wire tmp7115;
  wire tmp7116;
  wire tmp7117;
  wire tmp7118;
  wire tmp7119;
  wire tmp7120;
  wire tmp7121;
  wire tmp7122;
  wire tmp7123;
  wire tmp7124;
  wire tmp7125;
  wire tmp7126;
  wire tmp7127;
  wire tmp7128;
  wire tmp7129;
  wire tmp7130;
  wire tmp7131;
  wire tmp7132;
  wire tmp7133;
  wire tmp7134;
  wire tmp7135;
  wire tmp7136;
  wire tmp7137;
  wire tmp7138;
  wire tmp7139;
  wire tmp7140;
  wire tmp7141;
  wire tmp7142;
  wire tmp7143;
  wire tmp7144;
  wire tmp7145;
  wire tmp7146;
  wire tmp7147;
  wire tmp7148;
  wire tmp7149;
  wire tmp7150;
  wire tmp7151;
  wire tmp7152;
  wire tmp7153;
  wire tmp7154;
  wire tmp7155;
  wire tmp7156;
  wire tmp7157;
  wire tmp7158;
  wire tmp7159;
  wire tmp7160;
  wire tmp7161;
  wire tmp7162;
  wire tmp7163;
  wire tmp7164;
  wire tmp7165;
  wire tmp7166;
  wire tmp7167;
  wire tmp7168;
  wire tmp7169;
  wire tmp7170;
  wire tmp7171;
  wire tmp7172;
  wire tmp7173;
  wire tmp7174;
  wire tmp7175;
  wire tmp7176;
  wire tmp7177;
  wire tmp7178;
  wire tmp7179;
  wire tmp7180;
  wire tmp7181;
  wire tmp7182;
  wire tmp7183;
  wire tmp7184;
  wire tmp7185;
  wire tmp7186;
  wire tmp7187;
  wire tmp7188;
  wire tmp7189;
  wire tmp7190;
  wire tmp7191;
  wire tmp7192;
  wire tmp7193;
  wire tmp7194;
  wire tmp7195;
  wire tmp7196;
  wire tmp7197;
  wire tmp7198;
  wire tmp7199;
  wire tmp7200;
  wire tmp7201;
  wire tmp7202;
  wire tmp7203;
  wire tmp7204;
  wire tmp7205;
  wire tmp7206;
  wire tmp7207;
  wire tmp7208;
  wire tmp7209;
  wire tmp7210;
  wire tmp7211;
  wire tmp7212;
  wire tmp7213;
  wire tmp7214;
  wire tmp7215;
  wire tmp7216;
  wire tmp7217;
  wire tmp7218;
  wire tmp7219;
  wire tmp7220;
  wire tmp7221;
  wire tmp7222;
  wire tmp7223;
  wire tmp7224;
  wire tmp7225;
  wire tmp7226;
  wire tmp7227;
  wire tmp7228;
  wire tmp7229;
  wire tmp7230;
  wire tmp7231;
  wire tmp7232;
  wire tmp7233;
  wire tmp7234;
  wire tmp7235;
  wire tmp7236;
  wire tmp7237;
  wire tmp7238;
  wire tmp7239;
  wire tmp7240;
  wire tmp7241;
  wire tmp7242;
  wire tmp7243;
  wire tmp7244;
  wire tmp7245;
  wire tmp7246;
  wire tmp7247;
  wire tmp7248;
  wire tmp7249;
  wire tmp7250;
  wire tmp7251;
  wire tmp7252;
  wire tmp7253;
  wire tmp7254;
  wire tmp7255;
  wire tmp7256;
  wire tmp7257;
  wire tmp7258;
  wire tmp7259;
  wire tmp7260;
  wire tmp7261;
  wire tmp7262;
  wire tmp7263;
  wire tmp7264;
  wire tmp7265;
  wire tmp7266;
  wire tmp7267;
  wire tmp7268;
  wire tmp7269;
  wire tmp7270;
  wire tmp7271;
  wire tmp7272;
  wire tmp7273;
  wire tmp7274;
  wire tmp7275;
  wire tmp7276;
  wire tmp7277;
  wire tmp7278;
  wire tmp7279;
  wire tmp7280;
  wire tmp7281;
  wire tmp7282;
  wire tmp7283;
  wire tmp7284;
  wire tmp7285;
  wire tmp7286;
  wire tmp7287;
  wire tmp7288;
  wire tmp7289;
  wire tmp7290;
  wire tmp7291;
  wire tmp7292;
  wire tmp7293;
  wire tmp7294;
  wire tmp7295;
  wire tmp7296;
  wire tmp7297;
  wire tmp7298;
  wire tmp7299;
  wire tmp7300;
  wire tmp7301;
  wire tmp7302;
  wire tmp7303;
  wire tmp7304;
  wire tmp7305;
  wire tmp7306;
  wire tmp7307;
  wire tmp7308;
  wire tmp7309;
  wire tmp7310;
  wire tmp7311;
  wire tmp7312;
  wire tmp7313;
  wire tmp7314;
  wire tmp7315;
  wire tmp7316;
  wire tmp7317;
  wire tmp7318;
  wire tmp7319;
  wire tmp7320;
  wire tmp7321;
  wire tmp7322;
  wire tmp7323;
  wire tmp7324;
  wire tmp7325;
  wire tmp7326;
  wire tmp7327;
  wire tmp7328;
  wire tmp7329;
  wire tmp7330;
  wire tmp7331;
  wire tmp7332;
  wire tmp7333;
  wire tmp7334;
  wire tmp7335;
  wire tmp7336;
  wire tmp7337;
  wire tmp7338;
  wire tmp7339;
  wire tmp7340;
  wire tmp7341;
  wire tmp7342;
  wire tmp7343;
  wire tmp7344;
  wire tmp7345;
  wire tmp7346;
  wire tmp7347;
  wire tmp7348;
  wire tmp7349;
  wire tmp7350;
  wire tmp7351;
  wire tmp7352;
  wire tmp7353;
  wire tmp7354;
  wire tmp7355;
  wire tmp7356;
  wire tmp7357;
  wire tmp7358;
  wire tmp7359;
  wire tmp7360;
  wire tmp7361;
  wire tmp7362;
  wire tmp7363;
  wire tmp7364;
  wire tmp7365;
  wire tmp7366;
  wire tmp7367;
  wire tmp7368;
  wire tmp7369;
  wire tmp7370;
  wire tmp7371;
  wire tmp7372;
  wire tmp7373;
  wire tmp7374;
  wire tmp7375;
  wire tmp7376;
  wire tmp7377;
  wire tmp7378;
  wire tmp7379;
  wire tmp7380;
  wire tmp7381;
  wire tmp7382;
  wire tmp7383;
  wire tmp7384;
  wire tmp7385;
  wire tmp7386;
  wire tmp7387;
  wire tmp7388;
  wire tmp7389;
  wire tmp7390;
  wire tmp7391;
  wire tmp7392;
  wire tmp7393;
  wire tmp7394;
  wire tmp7395;
  wire tmp7396;
  wire tmp7397;
  wire tmp7398;
  wire tmp7399;
  wire tmp7400;
  wire tmp7401;
  wire tmp7402;
  wire tmp7403;
  wire tmp7404;
  wire tmp7405;
  wire tmp7406;
  wire tmp7407;
  wire tmp7408;
  wire tmp7409;
  wire tmp7410;
  wire tmp7411;
  wire tmp7412;
  wire tmp7413;
  wire tmp7414;
  wire tmp7415;
  wire tmp7416;
  wire tmp7417;
  wire tmp7418;
  wire tmp7419;
  wire tmp7420;
  wire tmp7421;
  wire tmp7422;
  wire tmp7423;
  wire tmp7424;
  wire tmp7425;
  wire tmp7426;
  wire tmp7427;
  wire tmp7428;
  wire tmp7429;
  wire tmp7430;
  wire tmp7431;
  wire tmp7432;
  wire tmp7433;
  wire tmp7434;
  wire tmp7435;
  wire tmp7436;
  wire tmp7437;
  wire tmp7438;
  wire tmp7439;
  wire tmp7440;
  wire tmp7441;
  wire tmp7442;
  wire tmp7443;
  wire tmp7444;
  wire tmp7445;
  wire tmp7446;
  wire tmp7447;
  wire tmp7448;
  wire tmp7449;
  wire tmp7450;
  wire tmp7451;
  wire tmp7452;
  wire tmp7453;
  wire tmp7454;
  wire tmp7455;
  wire tmp7456;
  wire tmp7457;
  wire tmp7458;
  wire tmp7459;
  wire tmp7460;
  wire tmp7461;
  wire tmp7462;
  wire tmp7463;
  wire tmp7464;
  wire tmp7465;
  wire tmp7466;
  wire tmp7467;
  wire tmp7468;
  wire tmp7469;
  wire tmp7470;
  wire tmp7471;
  wire tmp7472;
  wire tmp7473;
  wire tmp7474;
  wire tmp7475;
  wire tmp7476;
  wire tmp7477;
  wire tmp7478;
  wire tmp7479;
  wire tmp7480;
  wire tmp7481;
  wire tmp7482;
  wire tmp7483;
  wire tmp7484;
  wire tmp7485;
  wire tmp7486;
  wire tmp7487;
  wire tmp7488;
  wire tmp7489;
  wire tmp7490;
  wire tmp7491;
  wire tmp7492;
  wire tmp7493;
  wire tmp7494;
  wire tmp7495;
  wire tmp7496;
  wire tmp7497;
  wire tmp7498;
  wire tmp7499;
  wire tmp7500;
  wire tmp7501;
  wire tmp7502;
  wire tmp7503;
  wire tmp7504;
  wire tmp7505;
  wire tmp7506;
  wire tmp7507;
  wire tmp7508;
  wire tmp7509;
  wire tmp7510;
  wire tmp7511;
  wire tmp7512;
  wire tmp7513;
  wire tmp7514;
  wire tmp7515;
  wire tmp7516;
  wire tmp7517;
  wire tmp7518;
  wire tmp7519;
  wire tmp7520;
  wire tmp7521;
  wire tmp7522;
  wire tmp7523;
  wire tmp7524;
  wire tmp7525;
  wire tmp7526;
  wire tmp7527;
  wire tmp7528;
  wire tmp7529;
  wire tmp7530;
  wire tmp7531;
  wire tmp7532;
  wire tmp7533;
  wire tmp7534;
  wire tmp7535;
  wire tmp7536;
  wire tmp7537;
  wire tmp7538;
  wire tmp7539;
  wire tmp7540;
  wire tmp7541;
  wire tmp7542;
  wire tmp7543;
  wire tmp7544;
  wire tmp7545;
  wire tmp7546;
  wire tmp7547;
  wire tmp7548;
  wire tmp7549;
  wire tmp7550;
  wire tmp7551;
  wire tmp7552;
  wire tmp7553;
  wire tmp7554;
  wire tmp7555;
  wire tmp7556;
  wire tmp7557;
  wire tmp7558;
  wire tmp7559;
  wire tmp7560;
  wire tmp7561;
  wire tmp7562;
  wire tmp7563;
  wire tmp7564;
  wire tmp7565;
  wire tmp7566;
  wire tmp7567;
  wire tmp7568;
  wire tmp7569;
  wire tmp7570;
  wire tmp7571;
  wire tmp7572;
  wire tmp7573;
  wire tmp7574;
  wire tmp7575;
  wire tmp7576;
  wire tmp7577;
  wire tmp7578;
  wire tmp7579;
  wire tmp7580;
  wire tmp7581;
  wire tmp7582;
  wire tmp7583;
  wire tmp7584;
  wire tmp7585;
  wire tmp7586;
  wire tmp7587;
  wire tmp7588;
  wire tmp7589;
  wire tmp7590;
  wire tmp7591;
  wire tmp7592;
  wire tmp7593;
  wire tmp7594;
  wire tmp7595;
  wire tmp7596;
  wire tmp7597;
  wire tmp7598;
  wire tmp7599;
  wire tmp7600;
  wire tmp7601;
  wire tmp7602;
  wire tmp7603;
  wire tmp7604;
  wire tmp7605;
  wire tmp7606;
  wire tmp7607;
  wire tmp7608;
  wire tmp7609;
  wire tmp7610;
  wire tmp7611;
  wire tmp7612;
  wire tmp7613;
  wire tmp7614;
  wire tmp7615;
  wire tmp7616;
  wire tmp7617;
  wire tmp7618;
  wire tmp7619;
  wire tmp7620;
  wire tmp7621;
  wire tmp7622;
  wire tmp7623;
  wire tmp7624;
  wire tmp7625;
  wire tmp7626;
  wire tmp7627;
  wire tmp7628;
  wire tmp7629;
  wire tmp7630;
  wire tmp7631;
  wire tmp7632;
  wire tmp7633;
  wire tmp7634;
  wire tmp7635;
  wire tmp7636;
  wire tmp7637;
  wire tmp7638;
  wire tmp7639;
  wire tmp7640;
  wire tmp7641;
  wire tmp7642;
  wire tmp7643;
  wire tmp7644;
  wire tmp7645;
  wire tmp7646;
  wire tmp7647;
  wire tmp7648;
  wire tmp7649;
  wire tmp7650;
  wire tmp7651;
  wire tmp7652;
  wire tmp7653;
  wire tmp7654;
  wire tmp7655;
  wire tmp7656;
  wire tmp7657;
  wire tmp7658;
  wire tmp7659;
  wire tmp7660;
  wire tmp7661;
  wire tmp7662;
  wire tmp7663;
  wire tmp7664;
  wire tmp7665;
  wire tmp7666;
  wire tmp7667;
  wire tmp7668;
  wire tmp7669;
  wire tmp7670;
  wire tmp7671;
  wire tmp7672;
  wire tmp7673;
  wire tmp7674;
  wire tmp7675;
  wire tmp7676;
  wire tmp7677;
  wire tmp7678;
  wire tmp7679;
  wire tmp7680;
  wire tmp7681;
  wire tmp7682;
  wire tmp7683;
  wire tmp7684;
  wire tmp7685;
  wire tmp7686;
  wire tmp7687;
  wire tmp7688;
  wire tmp7689;
  wire tmp7690;
  wire tmp7691;
  wire tmp7692;
  wire tmp7693;
  wire tmp7694;
  wire tmp7695;
  wire tmp7696;
  wire tmp7697;
  wire tmp7698;
  wire tmp7699;
  wire tmp7700;
  wire tmp7701;
  wire tmp7702;
  wire tmp7703;
  wire tmp7704;
  wire tmp7705;
  wire tmp7706;
  wire tmp7707;
  wire tmp7708;
  wire tmp7709;
  wire tmp7710;
  wire tmp7711;
  wire tmp7712;
  wire tmp7713;
  wire tmp7714;
  wire tmp7715;
  wire tmp7716;
  wire tmp7717;
  wire tmp7718;
  wire tmp7719;
  wire tmp7720;
  wire tmp7721;
  wire tmp7722;
  wire tmp7723;
  wire tmp7724;
  wire tmp7725;
  wire tmp7726;
  wire tmp7727;
  wire tmp7728;
  wire tmp7729;
  wire tmp7730;
  wire tmp7731;
  wire tmp7732;
  wire tmp7733;
  wire tmp7734;
  wire tmp7735;
  wire tmp7736;
  wire tmp7737;
  wire tmp7738;
  wire tmp7739;
  wire tmp7740;
  wire tmp7741;
  wire tmp7742;
  wire tmp7743;
  wire tmp7744;
  wire tmp7745;
  wire tmp7746;
  wire tmp7747;
  wire tmp7748;
  wire tmp7749;
  wire tmp7750;
  wire tmp7751;
  wire tmp7752;
  wire tmp7753;
  wire tmp7754;
  wire tmp7755;
  wire tmp7756;
  wire tmp7757;
  wire tmp7758;
  wire tmp7759;
  wire tmp7760;
  wire tmp7761;
  wire tmp7762;
  wire tmp7763;
  wire tmp7764;
  wire tmp7765;
  wire tmp7766;
  wire tmp7767;
  wire tmp7768;
  wire tmp7769;
  wire tmp7770;
  wire tmp7771;
  wire tmp7772;
  wire tmp7773;
  wire tmp7774;
  wire tmp7775;
  wire tmp7776;
  wire tmp7777;
  wire tmp7778;
  wire tmp7779;
  wire tmp7780;
  wire tmp7781;
  wire tmp7782;
  wire tmp7783;
  wire tmp7784;
  wire tmp7785;
  wire tmp7786;
  wire tmp7787;
  wire tmp7788;
  wire tmp7789;
  wire tmp7790;
  wire tmp7791;
  wire tmp7792;
  wire tmp7793;
  wire tmp7794;
  wire tmp7795;
  wire tmp7796;
  wire tmp7797;
  wire tmp7798;
  wire tmp7799;
  wire tmp7800;
  wire tmp7801;
  wire tmp7802;
  wire tmp7803;
  wire tmp7804;
  wire tmp7805;
  wire tmp7806;
  wire tmp7807;
  wire tmp7808;
  wire tmp7809;
  wire tmp7810;
  wire tmp7811;
  wire tmp7812;
  wire tmp7813;
  wire tmp7814;
  wire tmp7815;
  wire tmp7816;
  wire tmp7817;
  wire tmp7818;
  wire tmp7819;
  wire tmp7820;
  wire tmp7821;
  wire tmp7822;
  wire tmp7823;
  wire tmp7824;
  wire tmp7825;
  wire tmp7826;
  wire tmp7827;
  wire tmp7828;
  wire tmp7829;
  wire tmp7830;
  wire tmp7831;
  wire tmp7832;
  wire tmp7833;
  wire tmp7834;
  wire tmp7835;
  wire tmp7836;
  wire tmp7837;
  wire tmp7838;
  wire tmp7839;
  wire tmp7840;
  wire tmp7841;
  wire tmp7842;
  wire tmp7843;
  wire tmp7844;
  wire tmp7845;
  wire tmp7846;
  wire tmp7847;
  wire tmp7848;
  wire tmp7849;
  wire tmp7850;
  wire tmp7851;
  wire tmp7852;
  wire tmp7853;
  wire tmp7854;
  wire tmp7855;
  wire tmp7856;
  wire tmp7857;
  wire tmp7858;
  wire tmp7859;
  wire tmp7860;
  wire tmp7861;
  wire tmp7862;
  wire tmp7863;
  wire tmp7864;
  wire tmp7865;
  wire tmp7866;
  wire tmp7867;
  wire tmp7868;
  wire tmp7869;
  wire tmp7870;
  wire tmp7871;
  wire tmp7872;
  wire tmp7873;
  wire tmp7874;
  wire tmp7875;
  wire tmp7876;
  wire tmp7877;
  wire tmp7878;
  wire tmp7879;
  wire tmp7880;
  wire tmp7881;
  wire tmp7882;
  wire tmp7883;
  wire tmp7884;
  wire tmp7885;
  wire tmp7886;
  wire tmp7887;
  wire tmp7888;
  wire tmp7889;
  wire tmp7890;
  wire tmp7891;
  wire tmp7892;
  wire tmp7893;
  wire tmp7894;
  wire tmp7895;
  wire tmp7896;
  wire tmp7897;
  wire tmp7898;
  wire tmp7899;
  wire tmp7900;
  wire tmp7901;
  wire tmp7902;
  wire tmp7903;
  wire tmp7904;
  wire tmp7905;
  wire tmp7906;
  wire tmp7907;
  wire tmp7908;
  wire tmp7909;
  wire tmp7910;
  wire tmp7911;
  wire tmp7912;
  wire tmp7913;
  wire tmp7914;
  wire tmp7915;
  wire tmp7916;
  wire tmp7917;
  wire tmp7918;
  wire tmp7919;
  wire tmp7920;
  wire tmp7921;
  wire tmp7922;
  wire tmp7923;
  wire tmp7924;
  wire tmp7925;
  wire tmp7926;
  wire tmp7927;
  wire tmp7928;
  wire tmp7929;
  wire tmp7930;
  wire tmp7931;
  wire tmp7932;
  wire tmp7933;
  wire tmp7934;
  wire tmp7935;
  wire tmp7936;
  wire tmp7937;
  wire tmp7938;
  wire tmp7939;
  wire tmp7940;
  wire tmp7941;
  wire tmp7942;
  wire tmp7943;
  wire tmp7944;
  wire tmp7945;
  wire tmp7946;
  wire tmp7947;
  wire tmp7948;
  wire tmp7949;
  wire tmp7950;
  wire tmp7951;
  wire tmp7952;
  wire tmp7953;
  wire tmp7954;
  wire tmp7955;
  wire tmp7956;
  wire tmp7957;
  wire tmp7958;
  wire tmp7959;
  wire tmp7960;
  wire tmp7961;
  wire tmp7962;
  wire tmp7963;
  wire tmp7964;
  wire tmp7965;
  wire tmp7966;
  wire tmp7967;
  wire tmp7968;
  wire tmp7969;
  wire tmp7970;
  wire tmp7971;
  wire tmp7972;
  wire tmp7973;
  wire tmp7974;
  wire tmp7975;
  wire tmp7976;
  wire tmp7977;
  wire tmp7978;
  wire tmp7979;
  wire tmp7980;
  wire tmp7981;
  wire tmp7982;
  wire tmp7983;
  wire tmp7984;
  wire tmp7985;
  wire tmp7986;
  wire tmp7987;
  wire tmp7988;
  wire tmp7989;
  wire tmp7990;
  wire tmp7991;
  wire tmp7992;
  wire tmp7993;
  wire tmp7994;
  wire tmp7995;
  wire tmp7996;
  wire tmp7997;
  wire tmp7998;
  wire tmp7999;
  wire tmp8000;
  wire tmp8001;
  wire tmp8002;
  wire tmp8003;
  wire tmp8004;
  wire tmp8005;
  wire tmp8006;
  wire tmp8007;
  wire tmp8008;
  wire tmp8009;
  wire tmp8010;
  wire tmp8011;
  wire tmp8012;
  wire tmp8013;
  wire tmp8014;
  wire tmp8015;
  wire tmp8016;
  wire tmp8017;
  wire tmp8018;
  wire tmp8019;
  wire tmp8020;
  wire tmp8021;
  wire tmp8022;
  wire tmp8023;
  wire tmp8024;
  wire tmp8025;
  wire tmp8026;
  wire tmp8027;
  wire tmp8028;
  wire tmp8029;
  wire tmp8030;
  wire tmp8031;
  wire tmp8032;
  wire tmp8033;
  wire tmp8034;
  wire tmp8035;
  wire tmp8036;
  wire tmp8037;
  wire tmp8038;
  wire tmp8039;
  wire tmp8040;
  wire tmp8041;
  wire tmp8042;
  wire tmp8043;
  wire tmp8044;
  wire tmp8045;
  wire tmp8046;
  wire tmp8047;
  wire tmp8048;
  wire tmp8049;
  wire tmp8050;
  wire tmp8051;
  wire tmp8052;
  wire tmp8053;
  wire tmp8054;
  wire tmp8055;
  wire tmp8056;
  wire tmp8057;
  wire tmp8058;
  wire tmp8059;
  wire tmp8060;
  wire tmp8061;
  wire tmp8062;
  wire tmp8063;
  wire tmp8064;
  wire tmp8065;
  wire tmp8066;
  wire tmp8067;
  wire tmp8068;
  wire tmp8069;
  wire tmp8070;
  wire tmp8071;
  wire tmp8072;
  wire tmp8073;
  wire tmp8074;
  wire tmp8075;
  wire tmp8076;
  wire tmp8077;
  wire tmp8078;
  wire tmp8079;
  wire tmp8080;
  wire tmp8081;
  wire tmp8082;
  wire tmp8083;
  wire tmp8084;
  wire tmp8085;
  wire tmp8086;
  wire tmp8087;
  wire tmp8088;
  wire tmp8089;
  wire tmp8090;
  wire tmp8091;
  wire tmp8092;
  wire tmp8093;
  wire tmp8094;
  wire tmp8095;
  wire tmp8096;
  wire tmp8097;
  wire tmp8098;
  wire tmp8099;
  wire tmp8100;
  wire tmp8101;
  wire tmp8102;
  wire tmp8103;
  wire tmp8104;
  wire tmp8105;
  wire tmp8106;
  wire tmp8107;
  wire tmp8108;
  wire tmp8109;
  wire tmp8110;
  wire tmp8111;
  wire tmp8112;
  wire tmp8113;
  wire tmp8114;
  wire tmp8115;
  wire tmp8116;
  wire tmp8117;
  wire tmp8118;
  wire tmp8119;
  wire tmp8120;
  wire tmp8121;
  wire tmp8122;
  wire tmp8123;
  wire tmp8124;
  wire tmp8125;
  wire tmp8126;
  wire tmp8127;
  wire tmp8128;
  wire tmp8129;
  wire tmp8130;
  wire tmp8131;
  wire tmp8132;
  wire tmp8133;
  wire tmp8134;
  wire tmp8135;
  wire tmp8136;
  wire tmp8137;
  wire tmp8138;
  wire tmp8139;
  wire tmp8140;
  wire tmp8141;
  wire tmp8142;
  wire tmp8143;
  wire tmp8144;
  wire tmp8145;
  wire tmp8146;
  wire tmp8147;
  wire tmp8148;
  wire tmp8149;
  wire tmp8150;
  wire tmp8151;
  wire tmp8152;
  wire tmp8153;
  wire tmp8154;
  wire tmp8155;
  wire tmp8156;
  wire tmp8157;
  wire tmp8158;
  wire tmp8159;
  wire tmp8160;
  wire tmp8161;
  wire tmp8162;
  wire tmp8163;
  wire tmp8164;
  wire tmp8165;
  wire tmp8166;
  wire tmp8167;
  wire tmp8168;
  wire tmp8169;
  wire tmp8170;
  wire tmp8171;
  wire tmp8172;
  wire tmp8173;
  wire tmp8174;
  wire tmp8175;
  wire tmp8176;
  wire tmp8177;
  wire tmp8178;
  wire tmp8179;
  wire tmp8180;
  wire tmp8181;
  wire tmp8182;
  wire tmp8183;
  wire tmp8184;
  wire tmp8185;
  wire tmp8186;
  wire tmp8187;
  wire tmp8188;
  wire tmp8189;
  wire tmp8190;
  wire tmp8191;
  wire tmp8192;
  wire tmp8193;
  wire tmp8194;
  wire tmp8195;
  wire tmp8196;
  wire tmp8197;
  wire tmp8198;
  wire tmp8199;
  wire tmp8200;
  wire tmp8201;
  wire tmp8202;
  wire tmp8203;
  wire tmp8204;
  wire tmp8205;
  wire tmp8206;
  wire tmp8207;
  wire tmp8208;
  wire tmp8209;
  wire tmp8210;
  wire tmp8211;
  wire tmp8212;
  wire tmp8213;
  wire tmp8214;
  wire tmp8215;
  wire tmp8216;
  wire tmp8217;
  wire tmp8218;
  wire tmp8219;
  wire tmp8220;
  wire tmp8221;
  wire tmp8222;
  wire tmp8223;
  wire tmp8224;
  wire tmp8225;
  wire tmp8226;
  wire tmp8227;
  wire tmp8228;
  wire tmp8229;
  wire tmp8230;
  wire tmp8231;
  wire tmp8232;
  wire tmp8233;
  wire tmp8234;
  wire tmp8235;
  wire tmp8236;
  wire tmp8237;
  wire tmp8238;
  wire tmp8239;
  wire tmp8240;
  wire tmp8241;
  wire tmp8242;
  wire tmp8243;
  wire tmp8244;
  wire tmp8245;
  wire tmp8246;
  wire tmp8247;
  wire tmp8248;
  wire tmp8249;
  wire tmp8250;
  wire tmp8251;
  wire tmp8252;
  wire tmp8253;
  wire tmp8254;
  wire tmp8255;
  wire tmp8256;
  wire tmp8257;
  wire tmp8258;
  wire tmp8259;
  wire tmp8260;
  wire tmp8261;
  wire tmp8262;
  wire tmp8263;
  wire tmp8264;
  wire tmp8265;
  wire tmp8266;
  wire tmp8267;
  wire tmp8268;
  wire tmp8269;
  wire tmp8270;
  wire tmp8271;
  wire tmp8272;
  wire tmp8273;
  wire tmp8274;
  wire tmp8275;
  wire tmp8276;
  wire tmp8277;
  wire tmp8278;
  wire tmp8279;
  wire tmp8280;
  wire tmp8281;
  wire tmp8282;
  wire tmp8283;
  wire tmp8284;
  wire tmp8285;
  wire tmp8286;
  wire tmp8287;
  wire tmp8288;
  wire tmp8289;
  wire tmp8290;
  wire tmp8291;
  wire tmp8292;
  wire tmp8293;
  wire tmp8294;
  wire tmp8295;
  wire tmp8296;
  wire tmp8297;
  wire tmp8298;
  wire tmp8299;
  wire tmp8300;
  wire tmp8301;
  wire tmp8302;
  wire tmp8303;
  wire tmp8304;
  wire tmp8305;
  wire tmp8306;
  wire tmp8307;
  wire tmp8308;
  wire tmp8309;
  wire tmp8310;
  wire tmp8311;
  wire tmp8312;
  wire tmp8313;
  wire tmp8314;
  wire tmp8315;
  wire tmp8316;
  wire tmp8317;
  wire tmp8318;
  wire tmp8319;
  wire tmp8320;
  wire tmp8321;
  wire tmp8322;
  wire tmp8323;
  wire tmp8324;
  wire tmp8325;
  wire tmp8326;
  wire tmp8327;
  wire tmp8328;
  wire tmp8329;
  wire tmp8330;
  wire tmp8331;
  wire tmp8332;
  wire tmp8333;
  wire tmp8334;
  wire tmp8335;
  wire tmp8336;
  wire tmp8337;
  wire tmp8338;
  wire tmp8339;
  wire tmp8340;
  wire tmp8341;
  wire tmp8342;
  wire tmp8343;
  wire tmp8344;
  wire tmp8345;
  wire tmp8346;
  wire tmp8347;
  wire tmp8348;
  wire tmp8349;
  wire tmp8350;
  wire tmp8351;
  wire tmp8352;
  wire tmp8353;
  wire tmp8354;
  wire tmp8355;
  wire tmp8356;
  wire tmp8357;
  wire tmp8358;
  wire tmp8359;
  wire tmp8360;
  wire tmp8361;
  wire tmp8362;
  wire tmp8363;
  wire tmp8364;
  wire tmp8365;
  wire tmp8366;
  wire tmp8367;
  wire tmp8368;
  wire tmp8369;
  wire tmp8370;
  wire tmp8371;
  wire tmp8372;
  wire tmp8373;
  wire tmp8374;
  wire tmp8375;
  wire tmp8376;
  wire tmp8377;
  wire tmp8378;
  wire tmp8379;
  wire tmp8380;
  wire tmp8381;
  wire tmp8382;
  wire tmp8383;
  wire tmp8384;
  wire tmp8385;
  wire tmp8386;
  wire tmp8387;
  wire tmp8388;
  wire tmp8389;
  wire tmp8390;
  wire tmp8391;
  wire tmp8392;
  wire tmp8393;
  wire tmp8394;
  wire tmp8395;
  wire tmp8396;
  wire tmp8397;
  wire tmp8398;
  wire tmp8399;
  wire tmp8400;
  wire tmp8401;
  wire tmp8402;
  wire tmp8403;
  wire tmp8404;
  wire tmp8405;
  wire tmp8406;
  wire tmp8407;
  wire tmp8408;
  wire tmp8409;
  wire tmp8410;
  wire tmp8411;
  wire tmp8412;
  wire tmp8413;
  wire tmp8414;
  wire tmp8415;
  wire tmp8416;
  wire tmp8417;
  wire tmp8418;
  wire tmp8419;
  wire tmp8420;
  wire tmp8421;
  wire tmp8422;
  wire tmp8423;
  wire tmp8424;
  wire tmp8425;
  wire tmp8426;
  wire tmp8427;
  wire tmp8428;
  wire tmp8429;
  wire tmp8430;
  wire tmp8431;
  wire tmp8432;
  wire tmp8433;
  wire tmp8434;
  wire tmp8435;
  wire tmp8436;
  wire tmp8437;
  wire tmp8438;
  wire tmp8439;
  wire tmp8440;
  wire tmp8441;
  wire tmp8442;
  wire tmp8443;
  wire tmp8444;
  wire tmp8445;
  wire tmp8446;
  wire tmp8447;
  wire tmp8448;
  wire tmp8449;
  wire tmp8450;
  wire tmp8451;
  wire tmp8452;
  wire tmp8453;
  wire tmp8454;
  wire tmp8455;
  wire tmp8456;
  wire tmp8457;
  wire tmp8458;
  wire tmp8459;
  wire tmp8460;
  wire tmp8461;
  wire tmp8462;
  wire tmp8463;
  wire tmp8464;
  wire tmp8465;
  wire tmp8466;
  wire tmp8467;
  wire tmp8468;
  wire tmp8469;
  wire tmp8470;
  wire tmp8471;
  wire tmp8472;
  wire tmp8473;
  wire tmp8474;
  wire tmp8475;
  wire tmp8476;
  wire tmp8477;
  wire tmp8478;
  wire tmp8479;
  wire tmp8480;
  wire tmp8481;
  wire tmp8482;
  wire tmp8483;
  wire tmp8484;
  wire tmp8485;
  wire tmp8486;
  wire tmp8487;
  wire tmp8488;
  wire tmp8489;
  wire tmp8490;
  wire tmp8491;
  wire tmp8492;
  wire tmp8493;
  wire tmp8494;
  wire tmp8495;
  wire tmp8496;
  wire tmp8497;
  wire tmp8498;
  wire tmp8499;
  wire tmp8500;
  wire tmp8501;
  wire tmp8502;
  wire tmp8503;
  wire tmp8504;
  wire tmp8505;
  wire tmp8506;
  wire tmp8507;
  wire tmp8508;
  wire tmp8509;
  wire tmp8510;
  wire tmp8511;
  wire tmp8512;
  wire tmp8513;
  wire tmp8514;
  wire tmp8515;
  wire tmp8516;
  wire tmp8517;
  wire tmp8518;
  wire tmp8519;
  wire tmp8520;
  wire tmp8521;
  wire tmp8522;
  wire tmp8523;
  wire tmp8524;
  wire tmp8525;
  wire tmp8526;
  wire tmp8527;
  wire tmp8528;
  wire tmp8529;
  wire tmp8530;
  wire tmp8531;
  wire tmp8532;
  wire tmp8533;
  wire tmp8534;
  wire tmp8535;
  wire tmp8536;
  wire tmp8537;
  wire tmp8538;
  wire tmp8539;
  wire tmp8540;
  wire tmp8541;
  wire tmp8542;
  wire tmp8543;
  wire tmp8544;
  wire tmp8545;
  wire tmp8546;
  wire tmp8547;
  wire tmp8548;
  wire tmp8549;
  wire tmp8550;
  wire tmp8551;
  wire tmp8552;
  wire tmp8553;
  wire tmp8554;
  wire tmp8555;
  wire tmp8556;
  wire tmp8557;
  wire tmp8558;
  wire tmp8559;
  wire tmp8560;
  wire tmp8561;
  wire tmp8562;
  wire tmp8563;
  wire tmp8564;
  wire tmp8565;
  wire tmp8566;
  wire tmp8567;
  wire tmp8568;
  wire tmp8569;
  wire tmp8570;
  wire tmp8571;
  wire tmp8572;
  wire tmp8573;
  wire tmp8574;
  wire tmp8575;
  wire tmp8576;
  wire tmp8577;
  wire tmp8578;
  wire tmp8579;
  wire tmp8580;
  wire tmp8581;
  wire tmp8582;
  wire tmp8583;
  wire tmp8584;
  wire tmp8585;
  wire tmp8586;
  wire tmp8587;
  wire tmp8588;
  wire tmp8589;
  wire tmp8590;
  wire tmp8591;
  wire tmp8592;
  wire tmp8593;
  wire tmp8594;
  wire tmp8595;
  wire tmp8596;
  wire tmp8597;
  wire tmp8598;
  wire tmp8599;
  wire tmp8600;
  wire tmp8601;
  wire tmp8602;
  wire tmp8603;
  wire tmp8604;
  wire tmp8605;
  wire tmp8606;
  wire tmp8607;
  wire tmp8608;
  wire tmp8609;
  wire tmp8610;
  wire tmp8611;
  wire tmp8612;
  wire tmp8613;
  wire tmp8614;
  wire tmp8615;
  wire tmp8616;
  wire tmp8617;
  wire tmp8618;
  wire tmp8619;
  wire tmp8620;
  wire tmp8621;
  wire tmp8622;
  wire tmp8623;
  wire tmp8624;
  wire tmp8625;
  wire tmp8626;
  wire tmp8627;
  wire tmp8628;
  wire tmp8629;
  wire tmp8630;
  wire tmp8631;
  wire tmp8632;
  wire tmp8633;
  wire tmp8634;
  wire tmp8635;
  wire tmp8636;
  wire tmp8637;
  wire tmp8638;
  wire tmp8639;
  wire tmp8640;
  wire tmp8641;
  wire tmp8642;
  wire tmp8643;
  wire tmp8644;
  wire tmp8645;
  wire tmp8646;
  wire tmp8647;
  wire tmp8648;
  wire tmp8649;
  wire tmp8650;
  wire tmp8651;
  wire tmp8652;
  wire tmp8653;
  wire tmp8654;
  wire tmp8655;
  wire tmp8656;
  wire tmp8657;
  wire tmp8658;
  wire tmp8659;
  wire tmp8660;
  wire tmp8661;
  wire tmp8662;
  wire tmp8663;
  wire tmp8664;
  wire tmp8665;
  wire tmp8666;
  wire tmp8667;
  wire tmp8668;
  wire tmp8669;
  wire tmp8670;
  wire tmp8671;
  wire tmp8672;
  wire tmp8673;
  wire tmp8674;
  wire tmp8675;
  wire tmp8676;
  wire tmp8677;
  wire tmp8678;
  wire tmp8679;
  wire tmp8680;
  wire tmp8681;
  wire tmp8682;
  wire tmp8683;
  wire tmp8684;
  wire tmp8685;
  wire tmp8686;
  wire tmp8687;
  wire tmp8688;
  wire tmp8689;
  wire tmp8690;
  wire tmp8691;
  wire tmp8692;
  wire tmp8693;
  wire tmp8694;
  wire tmp8695;
  wire tmp8696;
  wire tmp8697;
  wire tmp8698;
  wire tmp8699;
  wire tmp8700;
  wire tmp8701;
  wire tmp8702;
  wire tmp8703;
  wire tmp8704;
  wire tmp8705;
  wire tmp8706;
  wire tmp8707;
  wire tmp8708;
  wire tmp8709;
  wire tmp8710;
  wire tmp8711;
  wire tmp8712;
  wire tmp8713;
  wire tmp8714;
  wire tmp8715;
  wire tmp8716;
  wire tmp8717;
  wire tmp8718;
  wire tmp8719;
  wire tmp8720;
  wire tmp8721;
  wire tmp8722;
  wire tmp8723;
  wire tmp8724;
  wire tmp8725;
  wire tmp8726;
  wire tmp8727;
  wire tmp8728;
  wire tmp8729;
  wire tmp8730;
  wire tmp8731;
  wire tmp8732;
  wire tmp8733;
  wire tmp8734;
  wire tmp8735;
  wire tmp8736;
  wire tmp8737;
  wire tmp8738;
  wire tmp8739;
  wire tmp8740;
  wire tmp8741;
  wire tmp8742;
  wire tmp8743;
  wire tmp8744;
  wire tmp8745;
  wire tmp8746;
  wire tmp8747;
  wire tmp8748;
  wire tmp8749;
  wire tmp8750;
  wire tmp8751;
  wire tmp8752;
  wire tmp8753;
  wire tmp8754;
  wire tmp8755;
  wire tmp8756;
  wire tmp8757;
  wire tmp8758;
  wire tmp8759;
  wire tmp8760;
  wire tmp8761;
  wire tmp8762;
  wire tmp8763;
  wire tmp8764;
  wire tmp8765;
  wire tmp8766;
  wire tmp8767;
  wire tmp8768;
  wire tmp8769;
  wire tmp8770;
  wire tmp8771;
  wire tmp8772;
  wire tmp8773;
  wire tmp8774;
  wire tmp8775;
  wire tmp8776;
  wire tmp8777;
  wire tmp8778;
  wire tmp8779;
  wire tmp8780;
  wire tmp8781;
  wire tmp8782;
  wire tmp8783;
  wire tmp8784;
  wire tmp8785;
  wire tmp8786;
  wire tmp8787;
  wire tmp8788;
  wire tmp8789;
  wire tmp8790;
  wire tmp8791;
  wire tmp8792;
  wire tmp8793;
  wire tmp8794;
  wire tmp8795;
  wire tmp8796;
  wire tmp8797;
  wire tmp8798;
  wire tmp8799;
  wire tmp8800;
  wire tmp8801;
  wire tmp8802;
  wire tmp8803;
  wire tmp8804;
  wire tmp8805;
  wire tmp8806;
  wire tmp8807;
  wire tmp8808;
  wire tmp8809;
  wire tmp8810;
  wire tmp8811;
  wire tmp8812;
  wire tmp8813;
  wire tmp8814;
  wire tmp8815;
  wire tmp8816;
  wire tmp8817;
  wire tmp8818;
  wire tmp8819;
  wire tmp8820;
  wire tmp8821;
  wire tmp8822;
  wire tmp8823;
  wire tmp8824;
  wire tmp8825;
  wire tmp8826;
  wire tmp8827;
  wire tmp8828;
  wire tmp8829;
  wire tmp8830;
  wire tmp8831;
  wire tmp8832;
  wire tmp8833;
  wire tmp8834;
  wire tmp8835;
  wire tmp8836;
  wire tmp8837;
  wire tmp8838;
  wire tmp8839;
  wire tmp8840;
  wire tmp8841;
  wire tmp8842;
  wire tmp8843;
  wire tmp8844;
  wire tmp8845;
  wire tmp8846;
  wire tmp8847;
  wire tmp8848;
  wire tmp8849;
  wire tmp8850;
  wire tmp8851;
  wire tmp8852;
  wire tmp8853;
  wire tmp8854;
  wire tmp8855;
  wire tmp8856;
  wire tmp8857;
  wire tmp8858;
  wire tmp8859;
  wire tmp8860;
  wire tmp8861;
  wire tmp8862;
  wire tmp8863;
  wire tmp8864;
  wire tmp8865;
  wire tmp8866;
  wire tmp8867;
  wire tmp8868;
  wire tmp8869;
  wire tmp8870;
  wire tmp8871;
  wire tmp8872;
  wire tmp8873;
  wire tmp8874;
  wire tmp8875;
  wire tmp8876;
  wire tmp8877;
  wire tmp8878;
  wire tmp8879;
  wire tmp8880;
  wire tmp8881;
  wire tmp8882;
  wire tmp8883;
  wire tmp8884;
  wire tmp8885;
  wire tmp8886;
  wire tmp8887;
  wire tmp8888;
  wire tmp8889;
  wire tmp8890;
  wire tmp8891;
  wire tmp8892;
  wire tmp8893;
  wire tmp8894;
  wire tmp8895;
  wire tmp8896;
  wire tmp8897;
  wire tmp8898;
  wire tmp8899;
  wire tmp8900;
  wire tmp8901;
  wire tmp8902;
  wire tmp8903;
  wire tmp8904;
  wire tmp8905;
  wire tmp8906;
  wire tmp8907;
  wire tmp8908;
  wire tmp8909;
  wire tmp8910;
  wire tmp8911;
  wire tmp8912;
  wire tmp8913;
  wire tmp8914;
  wire tmp8915;
  wire tmp8916;
  wire tmp8917;
  wire tmp8918;
  wire tmp8919;
  wire tmp8920;
  wire tmp8921;
  wire tmp8922;
  wire tmp8923;
  wire tmp8924;
  wire tmp8925;
  wire tmp8926;
  wire tmp8927;
  wire tmp8928;
  wire tmp8929;
  wire tmp8930;
  wire tmp8931;
  wire tmp8932;
  wire tmp8933;
  wire tmp8934;
  wire tmp8935;
  wire tmp8936;
  wire tmp8937;
  wire tmp8938;
  wire tmp8939;
  wire tmp8940;
  wire tmp8941;
  wire tmp8942;
  wire tmp8943;
  wire tmp8944;
  wire tmp8945;
  wire tmp8946;
  wire tmp8947;
  wire tmp8948;
  wire tmp8949;
  wire tmp8950;
  wire tmp8951;
  wire tmp8952;
  wire tmp8953;
  wire tmp8954;
  wire tmp8955;
  wire tmp8956;
  wire tmp8957;
  wire tmp8958;
  wire tmp8959;
  wire tmp8960;
  wire tmp8961;
  wire tmp8962;
  wire tmp8963;
  wire tmp8964;
  wire tmp8965;
  wire tmp8966;
  wire tmp8967;
  wire tmp8968;
  wire tmp8969;
  wire tmp8970;
  wire tmp8971;
  wire tmp8972;
  wire tmp8973;
  wire tmp8974;
  wire tmp8975;
  wire tmp8976;
  wire tmp8977;
  wire tmp8978;
  wire tmp8979;
  wire tmp8980;
  wire tmp8981;
  wire tmp8982;
  wire tmp8983;
  wire tmp8984;
  wire tmp8985;
  wire tmp8986;
  wire tmp8987;
  wire tmp8988;
  wire tmp8989;
  wire tmp8990;
  wire tmp8991;

  reg s0;
  reg s1;
  reg s2;
  reg s3;
  reg s4;
  reg s5;
  reg s6;
  reg s7;
  reg s8;
  reg s9;
  reg s10;
  reg s11;
  reg s12;
  reg s13;
  reg s14;
  reg s15;
  reg s16;

  assign tmp9 = l3 ? 1 : 0;
  assign tmp8 = l1 ? tmp9 : 0;
  assign tmp12 = l1 ? 1 : 0;
  assign tmp11 = s0 ? tmp12 : tmp8;
  assign tmp10 = s1 ? tmp8 : tmp11;
  assign tmp7 = s2 ? tmp8 : tmp10;
  assign tmp16 = s1 ? tmp11 : 0;
  assign tmp17 = s0 ? tmp8 : 1;
  assign tmp15 = s2 ? tmp16 : tmp17;
  assign tmp19 = s1 ? 1 : 0;
  assign tmp20 = s1 ? tmp8 : tmp12;
  assign tmp18 = s2 ? tmp19 : tmp20;
  assign tmp14 = s3 ? tmp15 : tmp18;
  assign tmp24 = ~(l3 ? 1 : 0);
  assign tmp23 = s1 ? 1 : tmp24;
  assign tmp25 = ~(s1 ? tmp8 : tmp9);
  assign tmp22 = s2 ? tmp23 : tmp25;
  assign tmp26 = ~(l1 ? tmp9 : 0);
  assign tmp21 = ~(s3 ? tmp22 : tmp26);
  assign tmp13 = s4 ? tmp14 : tmp21;
  assign tmp6 = s5 ? tmp7 : tmp13;
  assign tmp29 = s6 ? 1 : tmp6;
  assign tmp34 = l2 ? 1 : tmp9;
  assign tmp35 = l2 ? 1 : 0;
  assign tmp33 = l1 ? tmp34 : tmp35;
  assign tmp38 = l1 ? 1 : tmp35;
  assign tmp37 = s0 ? tmp38 : tmp33;
  assign tmp36 = s1 ? tmp33 : tmp37;
  assign tmp32 = s2 ? tmp33 : tmp36;
  assign tmp42 = s1 ? tmp37 : tmp38;
  assign tmp43 = s0 ? tmp33 : 1;
  assign tmp41 = s2 ? tmp42 : tmp43;
  assign tmp46 = l1 ? tmp9 : tmp35;
  assign tmp45 = s1 ? tmp46 : tmp38;
  assign tmp44 = s2 ? tmp19 : tmp45;
  assign tmp40 = s3 ? tmp41 : tmp44;
  assign tmp49 = s1 ? tmp38 : tmp34;
  assign tmp50 = s1 ? tmp33 : tmp34;
  assign tmp48 = s2 ? tmp49 : tmp50;
  assign tmp47 = s3 ? tmp48 : tmp33;
  assign tmp39 = s4 ? tmp40 : tmp47;
  assign tmp31 = s5 ? tmp32 : tmp39;
  assign tmp30 = s6 ? tmp31 : 1;
  assign tmp28 = s7 ? tmp29 : tmp30;
  assign tmp51 = s7 ? tmp29 : tmp31;
  assign tmp27 = s8 ? tmp28 : tmp51;
  assign tmp5 = s9 ? tmp6 : tmp27;
  assign tmp55 = l1 ? 1 : tmp24;
  assign tmp57 = s0 ? tmp55 : tmp12;
  assign tmp56 = s1 ? tmp57 : tmp55;
  assign tmp54 = s2 ? tmp55 : tmp56;
  assign tmp61 = s1 ? tmp55 : 0;
  assign tmp63 = s0 ? tmp55 : 1;
  assign tmp62 = s1 ? tmp55 : tmp63;
  assign tmp60 = s2 ? tmp61 : tmp62;
  assign tmp65 = s1 ? tmp12 : tmp55;
  assign tmp64 = s2 ? tmp23 : tmp65;
  assign tmp59 = s3 ? tmp60 : tmp64;
  assign tmp67 = s2 ? 1 : tmp55;
  assign tmp66 = s3 ? tmp67 : tmp55;
  assign tmp58 = s4 ? tmp59 : tmp66;
  assign tmp53 = s5 ? tmp54 : tmp58;
  assign tmp71 = ~(s5 ? tmp54 : tmp58);
  assign tmp70 = s6 ? 1 : tmp71;
  assign tmp76 = l1 ? tmp35 : tmp34;
  assign tmp78 = l2 ? tmp9 : 0;
  assign tmp77 = l1 ? tmp78 : tmp34;
  assign tmp75 = s1 ? tmp76 : tmp77;
  assign tmp81 = l1 ? tmp35 : 1;
  assign tmp80 = s0 ? tmp77 : tmp81;
  assign tmp82 = s0 ? tmp76 : tmp77;
  assign tmp79 = s1 ? tmp80 : tmp82;
  assign tmp74 = s2 ? tmp75 : tmp79;
  assign tmp86 = s1 ? tmp77 : 1;
  assign tmp87 = s1 ? tmp76 : tmp80;
  assign tmp85 = s2 ? tmp86 : tmp87;
  assign tmp89 = s1 ? tmp12 : tmp24;
  assign tmp91 = ~(l1 ? tmp35 : tmp34);
  assign tmp90 = s1 ? tmp12 : tmp91;
  assign tmp88 = ~(s2 ? tmp89 : tmp90);
  assign tmp84 = s3 ? tmp85 : tmp88;
  assign tmp96 = ~(l2 ? 1 : 0);
  assign tmp95 = l1 ? 1 : tmp96;
  assign tmp94 = s1 ? tmp95 : 1;
  assign tmp97 = ~(l1 ? tmp78 : tmp34);
  assign tmp93 = s2 ? tmp94 : tmp97;
  assign tmp92 = ~(s3 ? tmp93 : tmp97);
  assign tmp83 = s4 ? tmp84 : tmp92;
  assign tmp73 = s5 ? tmp74 : tmp83;
  assign tmp72 = s6 ? tmp73 : 1;
  assign tmp69 = s7 ? tmp70 : tmp72;
  assign tmp100 = ~(s5 ? tmp74 : tmp83);
  assign tmp99 = ~(s6 ? tmp53 : tmp100);
  assign tmp98 = s7 ? tmp70 : tmp99;
  assign tmp68 = ~(s8 ? tmp69 : tmp98);
  assign tmp52 = ~(s9 ? tmp53 : tmp68);
  assign tmp4 = s11 ? tmp5 : tmp52;
  assign tmp105 = l1 ? tmp9 : 1;
  assign tmp107 = s0 ? 1 : tmp105;
  assign tmp106 = s1 ? tmp105 : tmp107;
  assign tmp104 = s2 ? tmp105 : tmp106;
  assign tmp111 = s1 ? tmp107 : 1;
  assign tmp112 = s0 ? tmp105 : 1;
  assign tmp110 = s2 ? tmp111 : tmp112;
  assign tmp115 = ~(l1 ? 1 : 0);
  assign tmp114 = s1 ? 1 : tmp115;
  assign tmp116 = s1 ? tmp105 : 1;
  assign tmp113 = s2 ? tmp114 : tmp116;
  assign tmp109 = s3 ? tmp110 : tmp113;
  assign tmp119 = s1 ? 1 : tmp105;
  assign tmp118 = s2 ? tmp119 : tmp105;
  assign tmp117 = s3 ? tmp118 : tmp105;
  assign tmp108 = s4 ? tmp109 : tmp117;
  assign tmp103 = s5 ? tmp104 : tmp108;
  assign tmp122 = s6 ? 1 : tmp103;
  assign tmp126 = l1 ? tmp34 : 1;
  assign tmp128 = s0 ? 1 : tmp126;
  assign tmp127 = s1 ? tmp126 : tmp128;
  assign tmp125 = s2 ? tmp126 : tmp127;
  assign tmp132 = s1 ? tmp128 : 1;
  assign tmp133 = s0 ? tmp126 : 1;
  assign tmp131 = s2 ? tmp132 : tmp133;
  assign tmp130 = s3 ? tmp131 : tmp113;
  assign tmp136 = s1 ? 1 : tmp126;
  assign tmp135 = s2 ? tmp136 : tmp126;
  assign tmp134 = s3 ? tmp135 : tmp126;
  assign tmp129 = s4 ? tmp130 : tmp134;
  assign tmp124 = s5 ? tmp125 : tmp129;
  assign tmp123 = s6 ? tmp124 : 1;
  assign tmp121 = s7 ? tmp122 : tmp123;
  assign tmp137 = s7 ? tmp122 : tmp124;
  assign tmp120 = s8 ? tmp121 : tmp137;
  assign tmp102 = s9 ? tmp103 : tmp120;
  assign tmp141 = l1 ? 1 : tmp9;
  assign tmp143 = s0 ? tmp141 : 1;
  assign tmp142 = s1 ? tmp143 : tmp141;
  assign tmp140 = s2 ? tmp141 : tmp142;
  assign tmp147 = s1 ? tmp141 : 1;
  assign tmp146 = s2 ? tmp147 : tmp143;
  assign tmp148 = s1 ? 1 : tmp141;
  assign tmp145 = s3 ? tmp146 : tmp148;
  assign tmp144 = s4 ? tmp145 : tmp141;
  assign tmp139 = s5 ? tmp140 : tmp144;
  assign tmp151 = s6 ? 1 : tmp139;
  assign tmp155 = l1 ? 1 : tmp34;
  assign tmp157 = s0 ? tmp155 : 1;
  assign tmp156 = s1 ? tmp157 : tmp155;
  assign tmp154 = s2 ? tmp155 : tmp156;
  assign tmp161 = s1 ? tmp155 : 1;
  assign tmp160 = s2 ? tmp161 : tmp157;
  assign tmp162 = s1 ? 1 : tmp155;
  assign tmp159 = s3 ? tmp160 : tmp162;
  assign tmp158 = s4 ? tmp159 : tmp155;
  assign tmp153 = s5 ? tmp154 : tmp158;
  assign tmp152 = s6 ? tmp153 : 1;
  assign tmp150 = s7 ? tmp151 : tmp152;
  assign tmp163 = s7 ? tmp151 : tmp153;
  assign tmp149 = s8 ? tmp150 : tmp163;
  assign tmp138 = s9 ? tmp139 : tmp149;
  assign tmp101 = s11 ? tmp102 : tmp138;
  assign tmp3 = s12 ? tmp4 : tmp101;
  assign tmp170 = s0 ? tmp9 : tmp141;
  assign tmp169 = s1 ? tmp141 : tmp170;
  assign tmp168 = s2 ? tmp141 : tmp169;
  assign tmp174 = s1 ? tmp170 : 1;
  assign tmp175 = s1 ? tmp141 : tmp143;
  assign tmp173 = s2 ? tmp174 : tmp175;
  assign tmp177 = s1 ? 1 : tmp9;
  assign tmp176 = s2 ? tmp148 : tmp177;
  assign tmp172 = s3 ? tmp173 : tmp176;
  assign tmp180 = ~(s1 ? tmp141 : tmp12);
  assign tmp179 = s2 ? tmp114 : tmp180;
  assign tmp181 = ~(l1 ? 1 : tmp9);
  assign tmp178 = ~(s3 ? tmp179 : tmp181);
  assign tmp171 = s4 ? tmp172 : tmp178;
  assign tmp167 = s5 ? tmp168 : tmp171;
  assign tmp185 = ~(s5 ? tmp168 : tmp171);
  assign tmp184 = s6 ? 1 : tmp185;
  assign tmp189 = l1 ? tmp35 : tmp24;
  assign tmp193 = l2 ? 1 : tmp24;
  assign tmp192 = l1 ? tmp35 : tmp193;
  assign tmp191 = s0 ? tmp189 : tmp192;
  assign tmp190 = s1 ? tmp189 : tmp191;
  assign tmp188 = s2 ? tmp189 : tmp190;
  assign tmp198 = s0 ? tmp193 : tmp189;
  assign tmp197 = s1 ? tmp198 : tmp12;
  assign tmp201 = l1 ? tmp35 : 0;
  assign tmp200 = s0 ? tmp189 : tmp201;
  assign tmp199 = s1 ? tmp189 : tmp200;
  assign tmp196 = s2 ? tmp197 : tmp199;
  assign tmp203 = s1 ? tmp81 : tmp181;
  assign tmp205 = ~(l2 ? 1 : tmp24);
  assign tmp204 = ~(s1 ? 1 : tmp205);
  assign tmp202 = s2 ? tmp203 : tmp204;
  assign tmp195 = s3 ? tmp196 : tmp202;
  assign tmp208 = s1 ? 1 : tmp81;
  assign tmp209 = s1 ? tmp189 : tmp81;
  assign tmp207 = s2 ? tmp208 : tmp209;
  assign tmp210 = s1 ? tmp189 : tmp192;
  assign tmp206 = s3 ? tmp207 : tmp210;
  assign tmp194 = s4 ? tmp195 : tmp206;
  assign tmp187 = s5 ? tmp188 : tmp194;
  assign tmp186 = s6 ? tmp187 : 1;
  assign tmp183 = s7 ? tmp184 : tmp186;
  assign tmp213 = ~(s5 ? tmp188 : tmp194);
  assign tmp212 = ~(s6 ? tmp167 : tmp213);
  assign tmp211 = s7 ? tmp184 : tmp212;
  assign tmp182 = ~(s8 ? tmp183 : tmp211);
  assign tmp166 = s9 ? tmp167 : tmp182;
  assign tmp214 = ~(s9 ? tmp6 : tmp27);
  assign tmp165 = s11 ? tmp166 : tmp214;
  assign tmp221 = s1 ? tmp8 : 0;
  assign tmp220 = s2 ? tmp221 : tmp8;
  assign tmp222 = s2 ? tmp19 : tmp8;
  assign tmp219 = s3 ? tmp220 : tmp222;
  assign tmp225 = s1 ? 1 : tmp26;
  assign tmp224 = s2 ? tmp225 : tmp26;
  assign tmp223 = ~(s3 ? tmp224 : tmp26);
  assign tmp218 = s4 ? tmp219 : tmp223;
  assign tmp217 = s5 ? tmp8 : tmp218;
  assign tmp229 = ~(s5 ? tmp8 : tmp218);
  assign tmp228 = s6 ? 1 : tmp229;
  assign tmp232 = l1 ? tmp193 : 1;
  assign tmp236 = s1 ? tmp232 : 1;
  assign tmp235 = s2 ? tmp236 : tmp232;
  assign tmp238 = s1 ? tmp81 : 1;
  assign tmp237 = s2 ? tmp238 : tmp232;
  assign tmp234 = s3 ? tmp235 : tmp237;
  assign tmp241 = s1 ? 1 : tmp232;
  assign tmp240 = s2 ? tmp241 : tmp232;
  assign tmp239 = s3 ? tmp240 : tmp232;
  assign tmp233 = s4 ? tmp234 : tmp239;
  assign tmp231 = s5 ? tmp232 : tmp233;
  assign tmp230 = s6 ? tmp231 : 1;
  assign tmp227 = s7 ? tmp228 : tmp230;
  assign tmp242 = s7 ? tmp228 : tmp231;
  assign tmp226 = ~(s8 ? tmp227 : tmp242);
  assign tmp216 = s9 ? tmp217 : tmp226;
  assign tmp247 = s2 ? tmp61 : tmp63;
  assign tmp249 = s1 ? 1 : tmp55;
  assign tmp248 = s2 ? tmp249 : tmp55;
  assign tmp246 = s3 ? tmp247 : tmp248;
  assign tmp252 = s1 ? tmp55 : 1;
  assign tmp251 = s2 ? 1 : tmp252;
  assign tmp250 = s3 ? tmp251 : tmp55;
  assign tmp245 = s4 ? tmp246 : tmp250;
  assign tmp244 = s5 ? tmp55 : tmp245;
  assign tmp255 = s6 ? 1 : tmp244;
  assign tmp258 = l1 ? 1 : tmp193;
  assign tmp262 = s1 ? tmp258 : tmp38;
  assign tmp263 = s0 ? tmp258 : 1;
  assign tmp261 = s2 ? tmp262 : tmp263;
  assign tmp264 = s2 ? tmp249 : tmp258;
  assign tmp260 = s3 ? tmp261 : tmp264;
  assign tmp267 = s1 ? tmp258 : 1;
  assign tmp266 = s2 ? 1 : tmp267;
  assign tmp265 = s3 ? tmp266 : tmp258;
  assign tmp259 = s4 ? tmp260 : tmp265;
  assign tmp257 = s5 ? tmp258 : tmp259;
  assign tmp256 = s6 ? tmp257 : 1;
  assign tmp254 = s7 ? tmp255 : tmp256;
  assign tmp268 = s7 ? tmp255 : tmp257;
  assign tmp253 = s8 ? tmp254 : tmp268;
  assign tmp243 = ~(s9 ? tmp244 : tmp253);
  assign tmp215 = s11 ? tmp216 : tmp243;
  assign tmp164 = ~(s12 ? tmp165 : tmp215);
  assign tmp2 = s13 ? tmp3 : tmp164;
  assign tmp281 = s1 ? tmp35 : tmp38;
  assign tmp283 = s0 ? tmp35 : tmp81;
  assign tmp282 = s1 ? tmp35 : tmp283;
  assign tmp280 = s2 ? tmp281 : tmp282;
  assign tmp285 = s1 ? tmp81 : 0;
  assign tmp286 = ~(s1 ? tmp95 : tmp96);
  assign tmp284 = s2 ? tmp285 : tmp286;
  assign tmp279 = s3 ? tmp280 : tmp284;
  assign tmp289 = s1 ? tmp38 : tmp201;
  assign tmp288 = s2 ? tmp289 : tmp35;
  assign tmp287 = s3 ? tmp288 : tmp35;
  assign tmp278 = s4 ? tmp279 : tmp287;
  assign tmp277 = s5 ? tmp35 : tmp278;
  assign tmp276 = s6 ? tmp277 : 1;
  assign tmp275 = s7 ? tmp29 : tmp276;
  assign tmp291 = ~(s6 ? tmp6 : tmp277);
  assign tmp290 = ~(s7 ? 1 : tmp291);
  assign tmp274 = ~(s8 ? tmp275 : tmp290);
  assign tmp273 = s9 ? 1 : tmp274;
  assign tmp299 = l1 ? tmp78 : tmp35;
  assign tmp298 = s1 ? tmp35 : tmp299;
  assign tmp301 = s0 ? tmp299 : tmp35;
  assign tmp302 = s0 ? tmp35 : tmp299;
  assign tmp300 = s1 ? tmp301 : tmp302;
  assign tmp297 = s2 ? tmp298 : tmp300;
  assign tmp306 = s1 ? tmp299 : tmp38;
  assign tmp308 = s0 ? tmp299 : tmp81;
  assign tmp307 = s1 ? tmp35 : tmp308;
  assign tmp305 = s2 ? tmp306 : tmp307;
  assign tmp310 = s1 ? tmp12 : 1;
  assign tmp311 = s1 ? tmp95 : tmp96;
  assign tmp309 = ~(s2 ? tmp310 : tmp311);
  assign tmp304 = s3 ? tmp305 : tmp309;
  assign tmp315 = ~(l1 ? 1 : tmp96);
  assign tmp314 = ~(s1 ? tmp299 : tmp315);
  assign tmp313 = s2 ? tmp94 : tmp314;
  assign tmp316 = ~(l1 ? tmp78 : tmp35);
  assign tmp312 = ~(s3 ? tmp313 : tmp316);
  assign tmp303 = s4 ? tmp304 : tmp312;
  assign tmp296 = s5 ? tmp297 : tmp303;
  assign tmp295 = s6 ? tmp296 : 1;
  assign tmp294 = s7 ? tmp70 : tmp295;
  assign tmp319 = ~(s5 ? tmp297 : tmp303);
  assign tmp318 = s6 ? tmp53 : tmp319;
  assign tmp317 = ~(s7 ? 1 : tmp318);
  assign tmp293 = ~(s8 ? tmp294 : tmp317);
  assign tmp292 = s9 ? 1 : tmp293;
  assign tmp272 = s11 ? tmp273 : tmp292;
  assign tmp323 = s7 ? tmp122 : tmp276;
  assign tmp325 = ~(s6 ? tmp103 : tmp277);
  assign tmp324 = ~(s7 ? 1 : tmp325);
  assign tmp322 = ~(s8 ? tmp323 : tmp324);
  assign tmp321 = s9 ? 1 : tmp322;
  assign tmp330 = s0 ? tmp105 : tmp9;
  assign tmp329 = s1 ? tmp330 : tmp105;
  assign tmp328 = s2 ? tmp105 : tmp329;
  assign tmp334 = s1 ? tmp105 : tmp112;
  assign tmp333 = s2 ? tmp116 : tmp334;
  assign tmp336 = s1 ? tmp9 : 1;
  assign tmp335 = s2 ? tmp114 : tmp336;
  assign tmp332 = s3 ? tmp333 : tmp335;
  assign tmp331 = s4 ? tmp332 : tmp117;
  assign tmp327 = s5 ? tmp328 : tmp331;
  assign tmp342 = l1 ? tmp193 : tmp35;
  assign tmp344 = s0 ? tmp342 : tmp193;
  assign tmp343 = s1 ? tmp344 : tmp342;
  assign tmp341 = s2 ? tmp342 : tmp343;
  assign tmp348 = s1 ? tmp342 : tmp38;
  assign tmp350 = s0 ? tmp342 : tmp81;
  assign tmp349 = s1 ? tmp342 : tmp350;
  assign tmp347 = s2 ? tmp348 : tmp349;
  assign tmp352 = s1 ? tmp81 : tmp12;
  assign tmp353 = s1 ? tmp193 : tmp35;
  assign tmp351 = s2 ? tmp352 : tmp353;
  assign tmp346 = s3 ? tmp347 : tmp351;
  assign tmp357 = l1 ? tmp193 : 0;
  assign tmp356 = s1 ? tmp38 : tmp357;
  assign tmp355 = s2 ? tmp356 : tmp342;
  assign tmp354 = s3 ? tmp355 : tmp342;
  assign tmp345 = s4 ? tmp346 : tmp354;
  assign tmp340 = s5 ? tmp341 : tmp345;
  assign tmp339 = s6 ? tmp340 : 1;
  assign tmp338 = s7 ? tmp151 : tmp339;
  assign tmp360 = ~(s5 ? tmp328 : tmp331);
  assign tmp359 = s6 ? 1 : tmp360;
  assign tmp361 = s6 ? tmp139 : tmp340;
  assign tmp358 = s7 ? tmp359 : tmp361;
  assign tmp337 = ~(s8 ? tmp338 : tmp358);
  assign tmp326 = s9 ? tmp327 : tmp337;
  assign tmp320 = s11 ? tmp321 : tmp326;
  assign tmp271 = s12 ? tmp272 : tmp320;
  assign tmp371 = ~(l2 ? tmp9 : 1);
  assign tmp370 = l1 ? tmp35 : tmp371;
  assign tmp373 = s0 ? tmp370 : tmp201;
  assign tmp374 = s0 ? tmp370 : tmp35;
  assign tmp372 = s1 ? tmp373 : tmp374;
  assign tmp369 = s2 ? tmp370 : tmp372;
  assign tmp379 = s0 ? tmp35 : tmp370;
  assign tmp378 = s1 ? tmp379 : tmp12;
  assign tmp380 = s1 ? tmp370 : tmp373;
  assign tmp377 = s2 ? tmp378 : tmp380;
  assign tmp382 = ~(s1 ? 1 : tmp96);
  assign tmp381 = s2 ? tmp285 : tmp382;
  assign tmp376 = s3 ? tmp377 : tmp381;
  assign tmp385 = s1 ? tmp370 : tmp35;
  assign tmp384 = s2 ? tmp289 : tmp385;
  assign tmp386 = s1 ? tmp201 : tmp35;
  assign tmp383 = s3 ? tmp384 : tmp386;
  assign tmp375 = s4 ? tmp376 : tmp383;
  assign tmp368 = s5 ? tmp369 : tmp375;
  assign tmp367 = s6 ? tmp368 : 1;
  assign tmp366 = s7 ? tmp184 : tmp367;
  assign tmp389 = ~(s5 ? tmp369 : tmp375);
  assign tmp388 = s6 ? tmp167 : tmp389;
  assign tmp387 = ~(s7 ? 1 : tmp388);
  assign tmp365 = ~(s8 ? tmp366 : tmp387);
  assign tmp364 = s9 ? 1 : tmp365;
  assign tmp363 = s11 ? tmp364 : tmp273;
  assign tmp393 = s7 ? tmp228 : tmp339;
  assign tmp396 = ~(s5 ? tmp341 : tmp345);
  assign tmp395 = ~(s6 ? tmp217 : tmp396);
  assign tmp394 = s7 ? tmp359 : tmp395;
  assign tmp392 = ~(s8 ? tmp393 : tmp394);
  assign tmp391 = s9 ? tmp327 : tmp392;
  assign tmp399 = s7 ? tmp255 : tmp339;
  assign tmp401 = s6 ? tmp244 : tmp340;
  assign tmp400 = s7 ? tmp359 : tmp401;
  assign tmp398 = ~(s8 ? tmp399 : tmp400);
  assign tmp397 = s9 ? tmp327 : tmp398;
  assign tmp390 = s11 ? tmp391 : tmp397;
  assign tmp362 = s12 ? tmp363 : tmp390;
  assign tmp270 = s13 ? tmp271 : tmp362;
  assign tmp402 = ~(s13 ? tmp3 : tmp164);
  assign tmp269 = ~(s15 ? tmp270 : tmp402);
  assign tmp1 = ~(s16 ? tmp2 : tmp269);
  assign recovery__1 = tmp1;

  assign tmp412 = l3 ? 1 : 0;
  assign tmp411 = l1 ? tmp412 : 0;
  assign tmp415 = l1 ? 1 : 0;
  assign tmp414 = s0 ? tmp415 : tmp411;
  assign tmp413 = s1 ? tmp411 : tmp414;
  assign tmp410 = s2 ? tmp411 : tmp413;
  assign tmp419 = s1 ? tmp414 : 0;
  assign tmp421 = s0 ? tmp411 : 0;
  assign tmp422 = s0 ? tmp411 : 1;
  assign tmp420 = s1 ? tmp421 : tmp422;
  assign tmp418 = s2 ? tmp419 : tmp420;
  assign tmp425 = s0 ? 1 : 0;
  assign tmp424 = s1 ? 1 : tmp425;
  assign tmp428 = ~(l1 ? tmp412 : 0);
  assign tmp427 = s0 ? 1 : tmp428;
  assign tmp429 = ~(s0 ? tmp411 : tmp415);
  assign tmp426 = ~(s1 ? tmp427 : tmp429);
  assign tmp423 = s2 ? tmp424 : tmp426;
  assign tmp417 = s3 ? tmp418 : tmp423;
  assign tmp433 = s0 ? tmp415 : 0;
  assign tmp435 = ~(l3 ? 1 : 0);
  assign tmp434 = ~(s0 ? 1 : tmp435);
  assign tmp432 = s1 ? tmp433 : tmp434;
  assign tmp437 = s0 ? tmp412 : tmp411;
  assign tmp438 = s0 ? 1 : tmp412;
  assign tmp436 = s1 ? tmp437 : tmp438;
  assign tmp431 = s2 ? tmp432 : tmp436;
  assign tmp441 = s0 ? 1 : tmp411;
  assign tmp440 = s1 ? tmp441 : tmp411;
  assign tmp439 = s2 ? tmp440 : tmp432;
  assign tmp430 = s3 ? tmp431 : tmp439;
  assign tmp416 = s4 ? tmp417 : tmp430;
  assign tmp409 = s5 ? tmp410 : tmp416;
  assign tmp445 = l2 ? 1 : tmp412;
  assign tmp446 = l2 ? 1 : 0;
  assign tmp444 = l1 ? tmp445 : tmp446;
  assign tmp449 = l1 ? 1 : tmp446;
  assign tmp448 = s0 ? tmp449 : tmp444;
  assign tmp447 = s1 ? tmp444 : tmp448;
  assign tmp443 = s2 ? tmp444 : tmp447;
  assign tmp453 = s1 ? tmp448 : tmp449;
  assign tmp455 = s0 ? tmp444 : tmp449;
  assign tmp456 = s0 ? tmp444 : 1;
  assign tmp454 = s1 ? tmp455 : tmp456;
  assign tmp452 = s2 ? tmp453 : tmp454;
  assign tmp460 = ~(l1 ? tmp412 : tmp446);
  assign tmp459 = s0 ? 1 : tmp460;
  assign tmp462 = l1 ? tmp412 : tmp446;
  assign tmp461 = ~(s0 ? tmp462 : tmp449);
  assign tmp458 = ~(s1 ? tmp459 : tmp461);
  assign tmp457 = s2 ? tmp424 : tmp458;
  assign tmp451 = s3 ? tmp452 : tmp457;
  assign tmp466 = s0 ? tmp449 : tmp445;
  assign tmp465 = s1 ? tmp449 : tmp466;
  assign tmp468 = s0 ? tmp445 : tmp444;
  assign tmp469 = s0 ? 1 : tmp445;
  assign tmp467 = s1 ? tmp468 : tmp469;
  assign tmp464 = s2 ? tmp465 : tmp467;
  assign tmp472 = s0 ? 1 : tmp444;
  assign tmp473 = s0 ? tmp462 : tmp444;
  assign tmp471 = s1 ? tmp472 : tmp473;
  assign tmp476 = ~(l2 ? 1 : tmp412);
  assign tmp475 = ~(s0 ? 1 : tmp476);
  assign tmp474 = s1 ? tmp449 : tmp475;
  assign tmp470 = s2 ? tmp471 : tmp474;
  assign tmp463 = s3 ? tmp464 : tmp470;
  assign tmp450 = s4 ? tmp451 : tmp463;
  assign tmp442 = s5 ? tmp443 : tmp450;
  assign tmp408 = s7 ? tmp409 : tmp442;
  assign tmp407 = s8 ? tmp408 : tmp409;
  assign tmp481 = l1 ? 1 : tmp435;
  assign tmp483 = s0 ? tmp481 : tmp415;
  assign tmp482 = s1 ? tmp483 : tmp481;
  assign tmp480 = s2 ? tmp481 : tmp482;
  assign tmp487 = s1 ? tmp481 : 0;
  assign tmp489 = s0 ? tmp481 : 0;
  assign tmp490 = s0 ? tmp481 : 1;
  assign tmp488 = s1 ? tmp489 : tmp490;
  assign tmp486 = s2 ? tmp487 : tmp488;
  assign tmp493 = s0 ? 1 : tmp435;
  assign tmp492 = s1 ? 1 : tmp493;
  assign tmp496 = ~(l1 ? 1 : 0);
  assign tmp495 = s0 ? tmp412 : tmp496;
  assign tmp497 = ~(s0 ? tmp415 : tmp481);
  assign tmp494 = ~(s1 ? tmp495 : tmp497);
  assign tmp491 = s2 ? tmp492 : tmp494;
  assign tmp485 = s3 ? tmp486 : tmp491;
  assign tmp500 = s1 ? tmp490 : 1;
  assign tmp501 = s1 ? tmp481 : 1;
  assign tmp499 = s2 ? tmp500 : tmp501;
  assign tmp504 = s0 ? 1 : tmp481;
  assign tmp505 = s0 ? tmp415 : tmp481;
  assign tmp503 = s1 ? tmp504 : tmp505;
  assign tmp507 = ~(s0 ? tmp412 : 0);
  assign tmp506 = s1 ? tmp490 : tmp507;
  assign tmp502 = s2 ? tmp503 : tmp506;
  assign tmp498 = s3 ? tmp499 : tmp502;
  assign tmp484 = s4 ? tmp485 : tmp498;
  assign tmp479 = s5 ? tmp480 : tmp484;
  assign tmp511 = l1 ? tmp446 : tmp445;
  assign tmp513 = l2 ? tmp412 : 0;
  assign tmp512 = l1 ? tmp513 : tmp445;
  assign tmp510 = s1 ? tmp511 : tmp512;
  assign tmp516 = l1 ? tmp446 : 1;
  assign tmp515 = s0 ? tmp512 : tmp516;
  assign tmp517 = s0 ? tmp511 : tmp512;
  assign tmp514 = s1 ? tmp515 : tmp517;
  assign tmp509 = s2 ? tmp510 : tmp514;
  assign tmp521 = s1 ? tmp512 : 1;
  assign tmp523 = s0 ? tmp511 : 1;
  assign tmp522 = s1 ? tmp523 : tmp515;
  assign tmp520 = s2 ? tmp521 : tmp522;
  assign tmp526 = s0 ? tmp516 : tmp496;
  assign tmp527 = ~(s0 ? tmp415 : tmp435);
  assign tmp525 = s1 ? tmp526 : tmp527;
  assign tmp530 = ~(l1 ? tmp446 : tmp445);
  assign tmp529 = ~(s0 ? tmp415 : tmp530);
  assign tmp528 = s1 ? tmp495 : tmp529;
  assign tmp524 = s2 ? tmp525 : tmp528;
  assign tmp519 = s3 ? tmp520 : tmp524;
  assign tmp536 = ~(l2 ? 1 : 0);
  assign tmp535 = ~(l1 ? 1 : tmp536);
  assign tmp534 = s0 ? tmp511 : tmp535;
  assign tmp538 = l1 ? 1 : tmp536;
  assign tmp537 = ~(s0 ? tmp538 : 1);
  assign tmp533 = s1 ? tmp534 : tmp537;
  assign tmp540 = s0 ? tmp516 : tmp535;
  assign tmp539 = s1 ? tmp512 : tmp540;
  assign tmp532 = s2 ? tmp533 : tmp539;
  assign tmp544 = l1 ? 1 : tmp476;
  assign tmp543 = s0 ? tmp415 : tmp544;
  assign tmp546 = ~(l1 ? tmp513 : tmp445);
  assign tmp545 = s0 ? tmp415 : tmp546;
  assign tmp542 = s1 ? tmp543 : tmp545;
  assign tmp548 = s0 ? tmp412 : 0;
  assign tmp547 = ~(s1 ? tmp534 : tmp548);
  assign tmp541 = ~(s2 ? tmp542 : tmp547);
  assign tmp531 = s3 ? tmp532 : tmp541;
  assign tmp518 = s4 ? tmp519 : tmp531;
  assign tmp508 = ~(s5 ? tmp509 : tmp518);
  assign tmp478 = s7 ? tmp479 : tmp508;
  assign tmp477 = ~(s8 ? tmp478 : tmp479);
  assign tmp406 = s11 ? tmp407 : tmp477;
  assign tmp554 = l1 ? tmp412 : 1;
  assign tmp556 = s0 ? 1 : tmp554;
  assign tmp555 = s1 ? tmp554 : tmp556;
  assign tmp553 = s2 ? tmp554 : tmp555;
  assign tmp560 = s1 ? tmp556 : 1;
  assign tmp561 = s0 ? tmp554 : 1;
  assign tmp559 = s2 ? tmp560 : tmp561;
  assign tmp564 = s0 ? 1 : tmp496;
  assign tmp563 = s1 ? 1 : tmp564;
  assign tmp565 = s1 ? tmp554 : tmp561;
  assign tmp562 = s2 ? tmp563 : tmp565;
  assign tmp558 = s3 ? tmp559 : tmp562;
  assign tmp568 = s1 ? 1 : tmp556;
  assign tmp567 = s2 ? tmp568 : tmp555;
  assign tmp570 = s1 ? tmp556 : tmp554;
  assign tmp571 = s1 ? 1 : tmp554;
  assign tmp569 = s2 ? tmp570 : tmp571;
  assign tmp566 = s3 ? tmp567 : tmp569;
  assign tmp557 = s4 ? tmp558 : tmp566;
  assign tmp552 = s5 ? tmp553 : tmp557;
  assign tmp574 = l1 ? tmp445 : 1;
  assign tmp576 = s0 ? 1 : tmp574;
  assign tmp575 = s1 ? tmp574 : tmp576;
  assign tmp573 = s2 ? tmp574 : tmp575;
  assign tmp580 = s1 ? tmp576 : 1;
  assign tmp581 = s0 ? tmp574 : 1;
  assign tmp579 = s2 ? tmp580 : tmp581;
  assign tmp578 = s3 ? tmp579 : tmp562;
  assign tmp584 = s1 ? 1 : tmp576;
  assign tmp583 = s2 ? tmp584 : tmp575;
  assign tmp586 = s1 ? tmp576 : tmp574;
  assign tmp587 = s1 ? 1 : tmp574;
  assign tmp585 = s2 ? tmp586 : tmp587;
  assign tmp582 = s3 ? tmp583 : tmp585;
  assign tmp577 = s4 ? tmp578 : tmp582;
  assign tmp572 = s5 ? tmp573 : tmp577;
  assign tmp551 = s7 ? tmp552 : tmp572;
  assign tmp550 = s8 ? tmp551 : tmp552;
  assign tmp592 = l1 ? 1 : tmp412;
  assign tmp594 = s0 ? tmp592 : 1;
  assign tmp593 = s1 ? tmp594 : tmp592;
  assign tmp591 = s2 ? tmp592 : tmp593;
  assign tmp598 = s1 ? tmp592 : 1;
  assign tmp597 = s2 ? tmp598 : tmp594;
  assign tmp601 = s0 ? 1 : tmp592;
  assign tmp600 = s1 ? 1 : tmp601;
  assign tmp602 = s1 ? tmp594 : tmp601;
  assign tmp599 = s2 ? tmp600 : tmp602;
  assign tmp596 = s3 ? tmp597 : tmp599;
  assign tmp606 = s0 ? 1 : tmp415;
  assign tmp605 = s1 ? tmp592 : tmp606;
  assign tmp604 = s2 ? tmp592 : tmp605;
  assign tmp607 = s2 ? tmp601 : tmp592;
  assign tmp603 = s3 ? tmp604 : tmp607;
  assign tmp595 = s4 ? tmp596 : tmp603;
  assign tmp590 = s5 ? tmp591 : tmp595;
  assign tmp610 = l1 ? 1 : tmp445;
  assign tmp612 = s0 ? tmp610 : 1;
  assign tmp611 = s1 ? tmp612 : tmp610;
  assign tmp609 = s2 ? tmp610 : tmp611;
  assign tmp616 = s1 ? tmp610 : 1;
  assign tmp615 = s2 ? tmp616 : tmp612;
  assign tmp619 = s0 ? 1 : tmp610;
  assign tmp618 = s1 ? tmp594 : tmp619;
  assign tmp617 = s2 ? tmp600 : tmp618;
  assign tmp614 = s3 ? tmp615 : tmp617;
  assign tmp623 = s0 ? 1 : tmp449;
  assign tmp622 = s1 ? tmp610 : tmp623;
  assign tmp621 = s2 ? tmp610 : tmp622;
  assign tmp624 = s2 ? tmp619 : tmp610;
  assign tmp620 = s3 ? tmp621 : tmp624;
  assign tmp613 = s4 ? tmp614 : tmp620;
  assign tmp608 = s5 ? tmp609 : tmp613;
  assign tmp589 = s7 ? tmp590 : tmp608;
  assign tmp588 = s8 ? tmp589 : tmp590;
  assign tmp549 = s11 ? tmp550 : tmp588;
  assign tmp405 = s12 ? tmp406 : tmp549;
  assign tmp632 = s0 ? tmp412 : tmp592;
  assign tmp631 = s1 ? tmp592 : tmp632;
  assign tmp630 = s2 ? tmp592 : tmp631;
  assign tmp636 = s1 ? tmp632 : 1;
  assign tmp635 = s2 ? tmp636 : tmp594;
  assign tmp638 = s1 ? tmp594 : tmp438;
  assign tmp637 = s2 ? tmp600 : tmp638;
  assign tmp634 = s3 ? tmp635 : tmp637;
  assign tmp642 = ~(s0 ? 1 : tmp496);
  assign tmp641 = s1 ? tmp548 : tmp642;
  assign tmp644 = s0 ? tmp415 : tmp592;
  assign tmp643 = s1 ? tmp644 : tmp606;
  assign tmp640 = s2 ? tmp641 : tmp643;
  assign tmp646 = s1 ? tmp601 : tmp592;
  assign tmp648 = s0 ? tmp592 : tmp415;
  assign tmp647 = s1 ? tmp548 : tmp648;
  assign tmp645 = s2 ? tmp646 : tmp647;
  assign tmp639 = s3 ? tmp640 : tmp645;
  assign tmp633 = s4 ? tmp634 : tmp639;
  assign tmp629 = s5 ? tmp630 : tmp633;
  assign tmp651 = l1 ? tmp446 : tmp435;
  assign tmp655 = l2 ? 1 : tmp435;
  assign tmp654 = l1 ? tmp446 : tmp655;
  assign tmp653 = s0 ? tmp651 : tmp654;
  assign tmp652 = s1 ? tmp651 : tmp653;
  assign tmp650 = s2 ? tmp651 : tmp652;
  assign tmp660 = s0 ? tmp655 : tmp651;
  assign tmp659 = s1 ? tmp660 : tmp415;
  assign tmp662 = s0 ? tmp651 : tmp415;
  assign tmp664 = l1 ? tmp446 : 0;
  assign tmp663 = s0 ? tmp651 : tmp664;
  assign tmp661 = s1 ? tmp662 : tmp663;
  assign tmp658 = s2 ? tmp659 : tmp661;
  assign tmp667 = s0 ? tmp664 : tmp516;
  assign tmp669 = ~(l1 ? 1 : tmp412);
  assign tmp668 = s0 ? tmp516 : tmp669;
  assign tmp666 = s1 ? tmp667 : tmp668;
  assign tmp672 = ~(l2 ? 1 : tmp435);
  assign tmp671 = s0 ? 1 : tmp672;
  assign tmp670 = ~(s1 ? tmp594 : tmp671);
  assign tmp665 = s2 ? tmp666 : tmp670;
  assign tmp657 = s3 ? tmp658 : tmp665;
  assign tmp676 = s0 ? tmp655 : 1;
  assign tmp677 = s0 ? 1 : tmp516;
  assign tmp675 = s1 ? tmp676 : tmp677;
  assign tmp679 = s0 ? tmp516 : tmp651;
  assign tmp678 = s1 ? tmp679 : tmp667;
  assign tmp674 = s2 ? tmp675 : tmp678;
  assign tmp683 = ~(l1 ? tmp446 : tmp655);
  assign tmp682 = ~(s0 ? 1 : tmp683);
  assign tmp681 = s1 ? tmp679 : tmp682;
  assign tmp686 = ~(l1 ? tmp446 : 1);
  assign tmp685 = ~(s0 ? tmp592 : tmp686);
  assign tmp684 = s1 ? tmp676 : tmp685;
  assign tmp680 = s2 ? tmp681 : tmp684;
  assign tmp673 = s3 ? tmp674 : tmp680;
  assign tmp656 = s4 ? tmp657 : tmp673;
  assign tmp649 = ~(s5 ? tmp650 : tmp656);
  assign tmp628 = s7 ? tmp629 : tmp649;
  assign tmp627 = s8 ? tmp628 : tmp629;
  assign tmp687 = ~(s8 ? tmp408 : tmp409);
  assign tmp626 = s11 ? tmp627 : tmp687;
  assign tmp695 = s1 ? tmp411 : 0;
  assign tmp696 = s1 ? tmp421 : tmp411;
  assign tmp694 = s2 ? tmp695 : tmp696;
  assign tmp698 = ~(s1 ? tmp427 : tmp428);
  assign tmp697 = s2 ? tmp424 : tmp698;
  assign tmp693 = s3 ? tmp694 : tmp697;
  assign tmp702 = ~(s0 ? 1 : tmp428);
  assign tmp701 = s1 ? tmp433 : tmp702;
  assign tmp700 = s2 ? tmp701 : tmp411;
  assign tmp703 = s2 ? tmp411 : tmp701;
  assign tmp699 = s3 ? tmp700 : tmp703;
  assign tmp692 = s4 ? tmp693 : tmp699;
  assign tmp691 = s5 ? tmp411 : tmp692;
  assign tmp705 = l1 ? tmp655 : 1;
  assign tmp709 = s1 ? tmp705 : 1;
  assign tmp711 = s0 ? tmp705 : 1;
  assign tmp710 = s1 ? tmp711 : tmp705;
  assign tmp708 = s2 ? tmp709 : tmp710;
  assign tmp714 = s0 ? tmp516 : 1;
  assign tmp713 = s1 ? tmp516 : tmp714;
  assign tmp715 = s1 ? tmp427 : tmp705;
  assign tmp712 = s2 ? tmp713 : tmp715;
  assign tmp707 = s3 ? tmp708 : tmp712;
  assign tmp719 = s0 ? 1 : tmp705;
  assign tmp718 = s1 ? tmp714 : tmp719;
  assign tmp717 = s2 ? tmp718 : tmp705;
  assign tmp720 = s2 ? tmp705 : tmp718;
  assign tmp716 = s3 ? tmp717 : tmp720;
  assign tmp706 = s4 ? tmp707 : tmp716;
  assign tmp704 = ~(s5 ? tmp705 : tmp706);
  assign tmp690 = s7 ? tmp691 : tmp704;
  assign tmp689 = s8 ? tmp690 : tmp691;
  assign tmp727 = s1 ? tmp481 : tmp490;
  assign tmp726 = s2 ? tmp481 : tmp727;
  assign tmp729 = s1 ? 1 : tmp504;
  assign tmp728 = s2 ? tmp729 : tmp481;
  assign tmp725 = s3 ? tmp726 : tmp728;
  assign tmp732 = s1 ? tmp504 : 1;
  assign tmp731 = s2 ? tmp500 : tmp732;
  assign tmp734 = s1 ? tmp504 : tmp481;
  assign tmp733 = s2 ? tmp734 : tmp490;
  assign tmp730 = s3 ? tmp731 : tmp733;
  assign tmp724 = s4 ? tmp725 : tmp730;
  assign tmp723 = s5 ? tmp481 : tmp724;
  assign tmp736 = l1 ? 1 : tmp655;
  assign tmp741 = s0 ? tmp736 : 1;
  assign tmp740 = s1 ? tmp736 : tmp741;
  assign tmp739 = s2 ? tmp736 : tmp740;
  assign tmp742 = s2 ? tmp729 : tmp736;
  assign tmp738 = s3 ? tmp739 : tmp742;
  assign tmp745 = s1 ? tmp741 : 1;
  assign tmp747 = s0 ? 1 : tmp736;
  assign tmp746 = s1 ? tmp747 : 1;
  assign tmp744 = s2 ? tmp745 : tmp746;
  assign tmp749 = s1 ? tmp747 : tmp736;
  assign tmp748 = s2 ? tmp749 : tmp741;
  assign tmp743 = s3 ? tmp744 : tmp748;
  assign tmp737 = s4 ? tmp738 : tmp743;
  assign tmp735 = s5 ? tmp736 : tmp737;
  assign tmp722 = s7 ? tmp723 : tmp735;
  assign tmp721 = ~(s8 ? tmp722 : tmp723);
  assign tmp688 = s11 ? tmp689 : tmp721;
  assign tmp625 = ~(s12 ? tmp626 : tmp688);
  assign tmp404 = s13 ? tmp405 : tmp625;
  assign tmp760 = s1 ? tmp446 : tmp449;
  assign tmp762 = s0 ? tmp446 : tmp449;
  assign tmp763 = s0 ? tmp446 : tmp516;
  assign tmp761 = s1 ? tmp762 : tmp763;
  assign tmp759 = s2 ? tmp760 : tmp761;
  assign tmp766 = s0 ? tmp516 : 0;
  assign tmp765 = s1 ? tmp516 : tmp766;
  assign tmp768 = s0 ? 1 : tmp538;
  assign tmp769 = s0 ? tmp538 : tmp536;
  assign tmp767 = ~(s1 ? tmp768 : tmp769);
  assign tmp764 = s2 ? tmp765 : tmp767;
  assign tmp758 = s3 ? tmp759 : tmp764;
  assign tmp773 = s0 ? tmp449 : tmp664;
  assign tmp772 = s1 ? tmp762 : tmp773;
  assign tmp775 = s0 ? tmp664 : tmp446;
  assign tmp776 = s0 ? tmp516 : tmp446;
  assign tmp774 = s1 ? tmp775 : tmp776;
  assign tmp771 = s2 ? tmp772 : tmp774;
  assign tmp779 = ~(s0 ? tmp538 : tmp536);
  assign tmp778 = s1 ? tmp776 : tmp779;
  assign tmp782 = ~(l1 ? tmp446 : 0);
  assign tmp781 = ~(s0 ? 1 : tmp782);
  assign tmp780 = s1 ? tmp762 : tmp781;
  assign tmp777 = s2 ? tmp778 : tmp780;
  assign tmp770 = s3 ? tmp771 : tmp777;
  assign tmp757 = s4 ? tmp758 : tmp770;
  assign tmp756 = s5 ? tmp446 : tmp757;
  assign tmp755 = s7 ? tmp409 : tmp756;
  assign tmp754 = s8 ? tmp755 : 0;
  assign tmp788 = l1 ? tmp513 : tmp446;
  assign tmp787 = s1 ? tmp446 : tmp788;
  assign tmp790 = s0 ? tmp788 : tmp446;
  assign tmp791 = s0 ? tmp446 : tmp788;
  assign tmp789 = s1 ? tmp790 : tmp791;
  assign tmp786 = s2 ? tmp787 : tmp789;
  assign tmp795 = s1 ? tmp788 : tmp449;
  assign tmp797 = s0 ? tmp788 : tmp516;
  assign tmp796 = s1 ? tmp762 : tmp797;
  assign tmp794 = s2 ? tmp795 : tmp796;
  assign tmp800 = ~(s0 ? tmp415 : 1);
  assign tmp799 = s1 ? tmp526 : tmp800;
  assign tmp798 = s2 ? tmp799 : tmp767;
  assign tmp793 = s3 ? tmp794 : tmp798;
  assign tmp804 = s0 ? tmp446 : tmp535;
  assign tmp803 = s1 ? tmp804 : tmp537;
  assign tmp807 = ~(l1 ? tmp513 : tmp446);
  assign tmp806 = s0 ? 1 : tmp807;
  assign tmp808 = ~(s0 ? tmp516 : tmp535);
  assign tmp805 = ~(s1 ? tmp806 : tmp808);
  assign tmp802 = s2 ? tmp803 : tmp805;
  assign tmp811 = s0 ? tmp415 : tmp538;
  assign tmp812 = s0 ? tmp538 : tmp807;
  assign tmp810 = s1 ? tmp811 : tmp812;
  assign tmp813 = ~(s1 ? tmp804 : 0);
  assign tmp809 = ~(s2 ? tmp810 : tmp813);
  assign tmp801 = s3 ? tmp802 : tmp809;
  assign tmp792 = s4 ? tmp793 : tmp801;
  assign tmp785 = ~(s5 ? tmp786 : tmp792);
  assign tmp784 = s7 ? tmp479 : tmp785;
  assign tmp783 = ~(s8 ? tmp784 : 1);
  assign tmp753 = s11 ? tmp754 : tmp783;
  assign tmp816 = s7 ? tmp552 : tmp756;
  assign tmp815 = s8 ? tmp816 : 0;
  assign tmp821 = l1 ? tmp655 : tmp446;
  assign tmp823 = s0 ? tmp821 : tmp655;
  assign tmp822 = s1 ? tmp823 : tmp821;
  assign tmp820 = s2 ? tmp821 : tmp822;
  assign tmp827 = s1 ? tmp821 : tmp449;
  assign tmp829 = s0 ? tmp821 : tmp449;
  assign tmp830 = s0 ? tmp821 : tmp516;
  assign tmp828 = s1 ? tmp829 : tmp830;
  assign tmp826 = s2 ? tmp827 : tmp828;
  assign tmp833 = s0 ? tmp516 : tmp415;
  assign tmp832 = s1 ? tmp516 : tmp833;
  assign tmp835 = s0 ? tmp415 : tmp655;
  assign tmp836 = s0 ? tmp655 : tmp446;
  assign tmp834 = s1 ? tmp835 : tmp836;
  assign tmp831 = s2 ? tmp832 : tmp834;
  assign tmp825 = s3 ? tmp826 : tmp831;
  assign tmp841 = l1 ? tmp655 : 0;
  assign tmp840 = s0 ? tmp449 : tmp841;
  assign tmp839 = s1 ? tmp762 : tmp840;
  assign tmp843 = s0 ? tmp841 : tmp821;
  assign tmp844 = s0 ? tmp516 : tmp821;
  assign tmp842 = s1 ? tmp843 : tmp844;
  assign tmp838 = s2 ? tmp839 : tmp842;
  assign tmp847 = s0 ? tmp655 : tmp821;
  assign tmp846 = s1 ? tmp844 : tmp847;
  assign tmp849 = s0 ? tmp415 : tmp841;
  assign tmp848 = s1 ? tmp762 : tmp849;
  assign tmp845 = s2 ? tmp846 : tmp848;
  assign tmp837 = s3 ? tmp838 : tmp845;
  assign tmp824 = s4 ? tmp825 : tmp837;
  assign tmp819 = s5 ? tmp820 : tmp824;
  assign tmp818 = s7 ? tmp590 : tmp819;
  assign tmp853 = s0 ? tmp554 : tmp412;
  assign tmp852 = s1 ? tmp853 : tmp554;
  assign tmp851 = s2 ? tmp554 : tmp852;
  assign tmp857 = s1 ? tmp554 : 1;
  assign tmp856 = s2 ? tmp857 : tmp561;
  assign tmp860 = s0 ? tmp415 : tmp435;
  assign tmp861 = ~(s0 ? tmp412 : 1);
  assign tmp859 = ~(s1 ? tmp860 : tmp861);
  assign tmp858 = s2 ? tmp563 : tmp859;
  assign tmp855 = s3 ? tmp856 : tmp858;
  assign tmp865 = s0 ? tmp412 : tmp554;
  assign tmp864 = s1 ? tmp556 : tmp865;
  assign tmp868 = ~(l1 ? tmp412 : 1);
  assign tmp867 = ~(s0 ? tmp415 : tmp868);
  assign tmp866 = s1 ? 1 : tmp867;
  assign tmp863 = s2 ? tmp864 : tmp866;
  assign tmp862 = s3 ? tmp567 : tmp863;
  assign tmp854 = s4 ? tmp855 : tmp862;
  assign tmp850 = ~(s5 ? tmp851 : tmp854);
  assign tmp817 = s8 ? tmp818 : tmp850;
  assign tmp814 = s11 ? tmp815 : tmp817;
  assign tmp752 = s12 ? tmp753 : tmp814;
  assign tmp876 = ~(l2 ? tmp412 : 1);
  assign tmp875 = l1 ? tmp446 : tmp876;
  assign tmp878 = s0 ? tmp875 : tmp664;
  assign tmp879 = s0 ? tmp875 : tmp446;
  assign tmp877 = s1 ? tmp878 : tmp879;
  assign tmp874 = s2 ? tmp875 : tmp877;
  assign tmp884 = s0 ? tmp446 : tmp875;
  assign tmp883 = s1 ? tmp884 : tmp415;
  assign tmp886 = s0 ? tmp875 : tmp415;
  assign tmp885 = s1 ? tmp886 : tmp878;
  assign tmp882 = s2 ? tmp883 : tmp885;
  assign tmp888 = s1 ? tmp667 : tmp766;
  assign tmp890 = s0 ? 1 : tmp536;
  assign tmp889 = ~(s1 ? 1 : tmp890);
  assign tmp887 = s2 ? tmp888 : tmp889;
  assign tmp881 = s3 ? tmp882 : tmp887;
  assign tmp894 = s0 ? tmp664 : tmp875;
  assign tmp893 = s1 ? tmp894 : tmp775;
  assign tmp892 = s2 ? tmp772 : tmp893;
  assign tmp897 = s0 ? tmp516 : tmp664;
  assign tmp898 = ~(s0 ? 1 : tmp536);
  assign tmp896 = s1 ? tmp897 : tmp898;
  assign tmp895 = s2 ? tmp896 : tmp780;
  assign tmp891 = s3 ? tmp892 : tmp895;
  assign tmp880 = s4 ? tmp881 : tmp891;
  assign tmp873 = ~(s5 ? tmp874 : tmp880);
  assign tmp872 = s7 ? tmp629 : tmp873;
  assign tmp871 = s8 ? tmp872 : 1;
  assign tmp899 = ~(s8 ? tmp755 : 0);
  assign tmp870 = s11 ? tmp871 : tmp899;
  assign tmp903 = ~(s5 ? tmp820 : tmp824);
  assign tmp902 = s7 ? tmp691 : tmp903;
  assign tmp904 = s5 ? tmp851 : tmp854;
  assign tmp901 = s8 ? tmp902 : tmp904;
  assign tmp906 = s7 ? tmp723 : tmp819;
  assign tmp905 = ~(s8 ? tmp906 : tmp850);
  assign tmp900 = s11 ? tmp901 : tmp905;
  assign tmp869 = ~(s12 ? tmp870 : tmp900);
  assign tmp751 = s13 ? tmp752 : tmp869;
  assign tmp750 = s15 ? tmp751 : tmp404;
  assign tmp403 = ~(s16 ? tmp404 : tmp750);
  assign recovery__2 = tmp403;

  assign tmp910 = s11 ? 1 : 0;
  assign tmp915 = l1 ? 1 : 0;
  assign tmp919 = s1 ? tmp915 : 0;
  assign tmp921 = s0 ? tmp915 : 0;
  assign tmp920 = s1 ? tmp921 : tmp915;
  assign tmp918 = s2 ? tmp919 : tmp920;
  assign tmp924 = s0 ? 1 : 0;
  assign tmp923 = s1 ? 1 : tmp924;
  assign tmp922 = s2 ? tmp923 : tmp915;
  assign tmp917 = s3 ? tmp918 : tmp922;
  assign tmp929 = ~(l1 ? 1 : 0);
  assign tmp928 = ~(s0 ? 1 : tmp929);
  assign tmp927 = s1 ? tmp921 : tmp928;
  assign tmp926 = s2 ? tmp927 : tmp915;
  assign tmp930 = s2 ? tmp915 : tmp921;
  assign tmp925 = s3 ? tmp926 : tmp930;
  assign tmp916 = s4 ? tmp917 : tmp925;
  assign tmp914 = s5 ? tmp915 : tmp916;
  assign tmp939 = s0 ? 1 : tmp929;
  assign tmp938 = ~(s1 ? tmp939 : tmp929);
  assign tmp937 = s2 ? tmp923 : tmp938;
  assign tmp936 = s3 ? tmp918 : tmp937;
  assign tmp941 = s2 ? tmp915 : tmp927;
  assign tmp940 = s3 ? tmp926 : tmp941;
  assign tmp935 = s4 ? tmp936 : tmp940;
  assign tmp934 = s5 ? tmp915 : tmp935;
  assign tmp933 = s6 ? tmp934 : tmp914;
  assign tmp946 = s2 ? tmp919 : tmp915;
  assign tmp948 = s1 ? 1 : 0;
  assign tmp947 = s2 ? tmp948 : tmp915;
  assign tmp945 = s3 ? tmp946 : tmp947;
  assign tmp951 = s1 ? 1 : tmp929;
  assign tmp950 = s2 ? tmp951 : tmp929;
  assign tmp949 = ~(s3 ? tmp950 : tmp929);
  assign tmp944 = s4 ? tmp945 : tmp949;
  assign tmp943 = s5 ? tmp915 : tmp944;
  assign tmp942 = s6 ? tmp943 : tmp934;
  assign tmp932 = s7 ? tmp933 : tmp942;
  assign tmp956 = s3 ? tmp946 : tmp922;
  assign tmp957 = s3 ? tmp926 : tmp915;
  assign tmp955 = s4 ? tmp956 : tmp957;
  assign tmp954 = s5 ? tmp915 : tmp955;
  assign tmp953 = s6 ? tmp934 : tmp954;
  assign tmp958 = s6 ? tmp954 : tmp943;
  assign tmp952 = s7 ? tmp953 : tmp958;
  assign tmp931 = s8 ? tmp932 : tmp952;
  assign tmp913 = s9 ? tmp914 : tmp931;
  assign tmp962 = s6 ? tmp914 : tmp943;
  assign tmp961 = s7 ? tmp933 : tmp962;
  assign tmp960 = s8 ? tmp932 : tmp961;
  assign tmp959 = s9 ? tmp914 : tmp960;
  assign tmp912 = s10 ? tmp913 : tmp959;
  assign tmp970 = s0 ? tmp915 : 1;
  assign tmp969 = s1 ? tmp921 : tmp970;
  assign tmp968 = s2 ? tmp919 : tmp969;
  assign tmp973 = s0 ? 1 : tmp915;
  assign tmp972 = s1 ? 1 : tmp973;
  assign tmp971 = s2 ? tmp972 : tmp915;
  assign tmp967 = s3 ? tmp968 : tmp971;
  assign tmp976 = s1 ? tmp915 : 1;
  assign tmp975 = s2 ? 1 : tmp976;
  assign tmp977 = s1 ? tmp973 : tmp915;
  assign tmp974 = s3 ? tmp975 : tmp977;
  assign tmp966 = s4 ? tmp967 : tmp974;
  assign tmp965 = s5 ? tmp915 : tmp966;
  assign tmp985 = s1 ? tmp970 : 1;
  assign tmp984 = s2 ? tmp985 : tmp976;
  assign tmp986 = s2 ? tmp977 : tmp970;
  assign tmp983 = s3 ? tmp984 : tmp986;
  assign tmp982 = s4 ? tmp967 : tmp983;
  assign tmp981 = s5 ? tmp915 : tmp982;
  assign tmp980 = s6 ? tmp981 : tmp965;
  assign tmp992 = s1 ? tmp915 : tmp970;
  assign tmp991 = s2 ? tmp919 : tmp992;
  assign tmp994 = s1 ? 1 : tmp915;
  assign tmp993 = s2 ? tmp994 : tmp915;
  assign tmp990 = s3 ? tmp991 : tmp993;
  assign tmp996 = s2 ? 1 : tmp915;
  assign tmp995 = s3 ? tmp996 : tmp915;
  assign tmp989 = s4 ? tmp990 : tmp995;
  assign tmp988 = s5 ? tmp915 : tmp989;
  assign tmp987 = s6 ? tmp988 : tmp981;
  assign tmp979 = s7 ? tmp980 : tmp987;
  assign tmp1002 = s2 ? tmp977 : tmp992;
  assign tmp1001 = s3 ? tmp976 : tmp1002;
  assign tmp1000 = s4 ? tmp967 : tmp1001;
  assign tmp999 = s5 ? tmp915 : tmp1000;
  assign tmp1005 = s3 ? tmp991 : tmp971;
  assign tmp1004 = s4 ? tmp1005 : tmp995;
  assign tmp1003 = s5 ? tmp915 : tmp1004;
  assign tmp998 = s6 ? tmp999 : tmp1003;
  assign tmp1006 = s6 ? tmp1003 : tmp988;
  assign tmp997 = s7 ? tmp998 : tmp1006;
  assign tmp978 = s8 ? tmp979 : tmp997;
  assign tmp964 = s9 ? tmp965 : tmp978;
  assign tmp1010 = s6 ? tmp999 : tmp965;
  assign tmp1011 = s6 ? tmp965 : tmp988;
  assign tmp1009 = s7 ? tmp1010 : tmp1011;
  assign tmp1008 = s8 ? tmp979 : tmp1009;
  assign tmp1007 = s9 ? tmp965 : tmp1008;
  assign tmp963 = s10 ? tmp964 : tmp1007;
  assign tmp911 = s11 ? tmp912 : tmp963;
  assign tmp909 = s12 ? tmp910 : tmp911;
  assign tmp1018 = s1 ? tmp915 : tmp928;
  assign tmp1017 = s2 ? tmp915 : tmp1018;
  assign tmp1022 = s1 ? tmp939 : 1;
  assign tmp1023 = ~(s0 ? tmp915 : 0);
  assign tmp1021 = s2 ? tmp1022 : tmp1023;
  assign tmp1024 = ~(s2 ? tmp915 : tmp919);
  assign tmp1020 = s3 ? tmp1021 : tmp1024;
  assign tmp1027 = s1 ? 1 : tmp939;
  assign tmp1026 = s2 ? tmp1027 : tmp929;
  assign tmp1029 = ~(s1 ? 1 : tmp929);
  assign tmp1028 = ~(s2 ? tmp915 : tmp1029);
  assign tmp1025 = s3 ? tmp1026 : tmp1028;
  assign tmp1019 = ~(s4 ? tmp1020 : tmp1025);
  assign tmp1016 = s5 ? tmp1017 : tmp1019;
  assign tmp1037 = ~(s1 ? tmp915 : tmp921);
  assign tmp1036 = s2 ? tmp1027 : tmp1037;
  assign tmp1035 = s3 ? tmp1021 : tmp1036;
  assign tmp1040 = ~(s1 ? tmp915 : tmp928);
  assign tmp1039 = s2 ? tmp1027 : tmp1040;
  assign tmp1042 = s1 ? tmp939 : tmp929;
  assign tmp1041 = s2 ? tmp1042 : tmp951;
  assign tmp1038 = s3 ? tmp1039 : tmp1041;
  assign tmp1034 = ~(s4 ? tmp1035 : tmp1038);
  assign tmp1033 = s5 ? tmp1017 : tmp1034;
  assign tmp1047 = ~(s1 ? tmp915 : 0);
  assign tmp1046 = s2 ? tmp951 : tmp1047;
  assign tmp1045 = s3 ? tmp1021 : tmp1046;
  assign tmp1044 = ~(s4 ? tmp1045 : tmp1025);
  assign tmp1043 = s5 ? tmp1017 : tmp1044;
  assign tmp1032 = s6 ? tmp1033 : tmp1043;
  assign tmp1052 = l2 ? 1 : 0;
  assign tmp1051 = l1 ? tmp1052 : 1;
  assign tmp1054 = s0 ? 1 : tmp1051;
  assign tmp1053 = s1 ? tmp1051 : tmp1054;
  assign tmp1050 = s2 ? tmp1051 : tmp1053;
  assign tmp1058 = s1 ? tmp1054 : 1;
  assign tmp1059 = s0 ? tmp1051 : 1;
  assign tmp1057 = s2 ? tmp1058 : tmp1059;
  assign tmp1056 = s3 ? tmp1057 : tmp1046;
  assign tmp1061 = s2 ? tmp951 : tmp1051;
  assign tmp1062 = s2 ? tmp1051 : tmp929;
  assign tmp1060 = s3 ? tmp1061 : tmp1062;
  assign tmp1055 = s4 ? tmp1056 : tmp1060;
  assign tmp1049 = s5 ? tmp1050 : tmp1055;
  assign tmp1065 = s3 ? tmp1057 : tmp1036;
  assign tmp1068 = s1 ? tmp1051 : tmp939;
  assign tmp1067 = s2 ? tmp1027 : tmp1068;
  assign tmp1070 = s1 ? tmp939 : tmp1051;
  assign tmp1069 = s2 ? tmp1070 : tmp951;
  assign tmp1066 = s3 ? tmp1067 : tmp1069;
  assign tmp1064 = s4 ? tmp1065 : tmp1066;
  assign tmp1063 = s5 ? tmp1050 : tmp1064;
  assign tmp1048 = ~(s6 ? tmp1049 : tmp1063);
  assign tmp1031 = s7 ? tmp1032 : tmp1048;
  assign tmp1077 = s1 ? tmp915 : tmp921;
  assign tmp1076 = ~(s2 ? tmp915 : tmp1077);
  assign tmp1075 = s3 ? tmp1021 : tmp1076;
  assign tmp1074 = ~(s4 ? tmp1075 : tmp1025);
  assign tmp1073 = s5 ? tmp1017 : tmp1074;
  assign tmp1081 = s2 ? tmp1022 : tmp929;
  assign tmp1080 = s3 ? tmp1081 : tmp1024;
  assign tmp1082 = s3 ? tmp1026 : tmp929;
  assign tmp1079 = ~(s4 ? tmp1080 : tmp1082);
  assign tmp1078 = s5 ? tmp1017 : tmp1079;
  assign tmp1072 = s6 ? tmp1073 : tmp1078;
  assign tmp1086 = s2 ? tmp1027 : tmp1051;
  assign tmp1085 = s3 ? tmp1086 : tmp1051;
  assign tmp1084 = s4 ? tmp1056 : tmp1085;
  assign tmp1083 = ~(s5 ? tmp1050 : tmp1084);
  assign tmp1071 = s7 ? tmp1072 : tmp1083;
  assign tmp1030 = s8 ? tmp1031 : tmp1071;
  assign tmp1015 = s9 ? tmp1016 : tmp1030;
  assign tmp1090 = s6 ? tmp1073 : tmp1016;
  assign tmp1094 = s2 ? tmp1051 : tmp951;
  assign tmp1093 = s3 ? tmp1086 : tmp1094;
  assign tmp1092 = s4 ? tmp1056 : tmp1093;
  assign tmp1091 = ~(s5 ? tmp1050 : tmp1092);
  assign tmp1089 = s7 ? tmp1090 : tmp1091;
  assign tmp1088 = s8 ? tmp1031 : tmp1089;
  assign tmp1087 = s9 ? tmp1016 : tmp1088;
  assign tmp1014 = s10 ? tmp1015 : tmp1087;
  assign tmp1100 = s2 ? tmp915 : tmp992;
  assign tmp1101 = s2 ? tmp972 : tmp994;
  assign tmp1099 = s3 ? tmp1100 : tmp1101;
  assign tmp1104 = ~(s1 ? tmp915 : tmp973);
  assign tmp1103 = s2 ? tmp1027 : tmp1104;
  assign tmp1105 = ~(s2 ? tmp977 : tmp1029);
  assign tmp1102 = ~(s3 ? tmp1103 : tmp1105);
  assign tmp1098 = s4 ? tmp1099 : tmp1102;
  assign tmp1097 = s5 ? tmp915 : tmp1098;
  assign tmp1112 = s2 ? tmp976 : tmp970;
  assign tmp1114 = s1 ? tmp970 : tmp973;
  assign tmp1113 = s2 ? tmp972 : tmp1114;
  assign tmp1111 = s3 ? tmp1112 : tmp1113;
  assign tmp1117 = s1 ? tmp915 : tmp973;
  assign tmp1116 = s2 ? tmp927 : tmp1117;
  assign tmp1118 = s2 ? tmp977 : tmp920;
  assign tmp1115 = s3 ? tmp1116 : tmp1118;
  assign tmp1110 = s4 ? tmp1111 : tmp1115;
  assign tmp1109 = s5 ? tmp915 : tmp1110;
  assign tmp1122 = s2 ? tmp976 : tmp992;
  assign tmp1121 = s3 ? tmp1122 : tmp1101;
  assign tmp1120 = s4 ? tmp1121 : tmp1102;
  assign tmp1119 = s5 ? tmp915 : tmp1120;
  assign tmp1108 = s6 ? tmp1109 : tmp1119;
  assign tmp1126 = l1 ? 1 : tmp1052;
  assign tmp1128 = s0 ? tmp1126 : tmp915;
  assign tmp1127 = s1 ? tmp1126 : tmp1128;
  assign tmp1125 = s2 ? tmp1126 : tmp1127;
  assign tmp1133 = s0 ? tmp915 : tmp1126;
  assign tmp1132 = s1 ? tmp1133 : 1;
  assign tmp1135 = s0 ? tmp1126 : 1;
  assign tmp1134 = s1 ? tmp1126 : tmp1135;
  assign tmp1131 = s2 ? tmp1132 : tmp1134;
  assign tmp1130 = s3 ? tmp1131 : tmp994;
  assign tmp1138 = ~(s1 ? tmp1126 : tmp915);
  assign tmp1137 = s2 ? tmp951 : tmp1138;
  assign tmp1136 = ~(s3 ? tmp1137 : tmp1138);
  assign tmp1129 = s4 ? tmp1130 : tmp1136;
  assign tmp1124 = s5 ? tmp1125 : tmp1129;
  assign tmp1142 = s2 ? tmp1132 : tmp1135;
  assign tmp1141 = s3 ? tmp1142 : tmp1113;
  assign tmp1145 = s1 ? tmp1133 : tmp973;
  assign tmp1144 = s2 ? tmp927 : tmp1145;
  assign tmp1148 = s0 ? 1 : tmp1126;
  assign tmp1147 = s1 ? tmp1148 : tmp973;
  assign tmp1146 = s2 ? tmp1147 : tmp920;
  assign tmp1143 = s3 ? tmp1144 : tmp1146;
  assign tmp1140 = s4 ? tmp1141 : tmp1143;
  assign tmp1139 = s5 ? tmp1125 : tmp1140;
  assign tmp1123 = s6 ? tmp1124 : tmp1139;
  assign tmp1107 = s7 ? tmp1108 : tmp1123;
  assign tmp1153 = s3 ? tmp1100 : tmp1113;
  assign tmp1152 = s4 ? tmp1153 : tmp1115;
  assign tmp1151 = s5 ? tmp915 : tmp1152;
  assign tmp1156 = ~(s3 ? tmp1026 : tmp929);
  assign tmp1155 = s4 ? tmp1099 : tmp1156;
  assign tmp1154 = s5 ? tmp915 : tmp1155;
  assign tmp1150 = s6 ? tmp1151 : tmp1154;
  assign tmp1159 = s4 ? tmp1121 : tmp1156;
  assign tmp1158 = s5 ? tmp915 : tmp1159;
  assign tmp1157 = s6 ? tmp1158 : tmp1124;
  assign tmp1149 = s7 ? tmp1150 : tmp1157;
  assign tmp1106 = s8 ? tmp1107 : tmp1149;
  assign tmp1096 = s9 ? tmp1097 : tmp1106;
  assign tmp1163 = s6 ? tmp1151 : tmp1097;
  assign tmp1164 = s6 ? tmp1119 : tmp1124;
  assign tmp1162 = s7 ? tmp1163 : tmp1164;
  assign tmp1161 = s8 ? tmp1107 : tmp1162;
  assign tmp1160 = s9 ? tmp1097 : tmp1161;
  assign tmp1095 = s10 ? tmp1096 : tmp1160;
  assign tmp1013 = ~(s11 ? tmp1014 : tmp1095);
  assign tmp1012 = ~(s12 ? tmp910 : tmp1013);
  assign tmp908 = s13 ? tmp909 : tmp1012;
  assign tmp1170 = s8 ? tmp933 : tmp954;
  assign tmp1171 = s8 ? tmp933 : tmp914;
  assign tmp1169 = s10 ? tmp1170 : tmp1171;
  assign tmp1175 = s7 ? tmp980 : 1;
  assign tmp1177 = s6 ? tmp1003 : 1;
  assign tmp1176 = s7 ? 1 : tmp1177;
  assign tmp1174 = s8 ? tmp1175 : tmp1176;
  assign tmp1173 = s9 ? 1 : tmp1174;
  assign tmp1181 = s6 ? tmp965 : 1;
  assign tmp1180 = s7 ? 1 : tmp1181;
  assign tmp1179 = s8 ? tmp1175 : tmp1180;
  assign tmp1178 = s9 ? 1 : tmp1179;
  assign tmp1172 = s10 ? tmp1173 : tmp1178;
  assign tmp1168 = s11 ? tmp1169 : tmp1172;
  assign tmp1167 = s12 ? tmp910 : tmp1168;
  assign tmp1193 = ~(s1 ? 1 : 0);
  assign tmp1192 = s2 ? tmp948 : tmp1193;
  assign tmp1191 = s3 ? tmp1057 : tmp1192;
  assign tmp1195 = s2 ? tmp948 : tmp1051;
  assign tmp1194 = s3 ? tmp1195 : tmp1051;
  assign tmp1190 = s4 ? tmp1191 : tmp1194;
  assign tmp1189 = s5 ? tmp1050 : tmp1190;
  assign tmp1200 = ~(s1 ? 1 : tmp924);
  assign tmp1199 = s2 ? tmp923 : tmp1200;
  assign tmp1198 = s3 ? tmp1057 : tmp1199;
  assign tmp1202 = s2 ? tmp923 : tmp1068;
  assign tmp1204 = s1 ? tmp924 : tmp1051;
  assign tmp1203 = s2 ? tmp1204 : tmp948;
  assign tmp1201 = s3 ? tmp1202 : tmp1203;
  assign tmp1197 = s4 ? tmp1198 : tmp1201;
  assign tmp1196 = s5 ? tmp1050 : tmp1197;
  assign tmp1188 = ~(s6 ? tmp1189 : tmp1196);
  assign tmp1187 = s7 ? tmp1032 : tmp1188;
  assign tmp1208 = ~(s4 ? tmp1045 : tmp1082);
  assign tmp1207 = s5 ? tmp1017 : tmp1208;
  assign tmp1209 = ~(s5 ? tmp1050 : tmp1190);
  assign tmp1206 = s6 ? tmp1207 : tmp1209;
  assign tmp1205 = s7 ? 1 : tmp1206;
  assign tmp1186 = s8 ? tmp1187 : tmp1205;
  assign tmp1185 = s9 ? 1 : tmp1186;
  assign tmp1213 = s6 ? tmp1043 : tmp1209;
  assign tmp1212 = s7 ? 1 : tmp1213;
  assign tmp1211 = s8 ? tmp1187 : tmp1212;
  assign tmp1210 = s9 ? 1 : tmp1211;
  assign tmp1184 = s10 ? tmp1185 : tmp1210;
  assign tmp1217 = s7 ? tmp1108 : 1;
  assign tmp1219 = s6 ? tmp1158 : 1;
  assign tmp1218 = s7 ? 1 : tmp1219;
  assign tmp1216 = s8 ? tmp1217 : tmp1218;
  assign tmp1215 = s9 ? 1 : tmp1216;
  assign tmp1223 = s6 ? tmp1119 : 1;
  assign tmp1222 = s7 ? 1 : tmp1223;
  assign tmp1221 = s8 ? tmp1217 : tmp1222;
  assign tmp1220 = s9 ? 1 : tmp1221;
  assign tmp1214 = s10 ? tmp1215 : tmp1220;
  assign tmp1183 = ~(s11 ? tmp1184 : tmp1214);
  assign tmp1182 = ~(s12 ? tmp910 : tmp1183);
  assign tmp1166 = s13 ? tmp1167 : tmp1182;
  assign tmp1235 = s2 ? tmp985 : 1;
  assign tmp1234 = s3 ? 1 : tmp1235;
  assign tmp1238 = s1 ? 1 : tmp970;
  assign tmp1237 = s2 ? 1 : tmp1238;
  assign tmp1236 = s3 ? tmp1237 : 1;
  assign tmp1233 = s4 ? tmp1234 : tmp1236;
  assign tmp1232 = s5 ? 1 : tmp1233;
  assign tmp1231 = s6 ? tmp1232 : 1;
  assign tmp1230 = s7 ? 1 : tmp1231;
  assign tmp1242 = s4 ? tmp1234 : 1;
  assign tmp1241 = s5 ? 1 : tmp1242;
  assign tmp1240 = s6 ? 1 : tmp1241;
  assign tmp1239 = s7 ? 1 : tmp1240;
  assign tmp1229 = s8 ? tmp1230 : tmp1239;
  assign tmp1228 = s9 ? 1 : tmp1229;
  assign tmp1246 = s6 ? 1 : tmp1232;
  assign tmp1245 = s7 ? 1 : tmp1246;
  assign tmp1244 = s8 ? tmp1230 : tmp1245;
  assign tmp1243 = s9 ? 1 : tmp1244;
  assign tmp1227 = s10 ? tmp1228 : tmp1243;
  assign tmp1255 = s2 ? tmp1027 : tmp1022;
  assign tmp1254 = s3 ? tmp1255 : 1;
  assign tmp1253 = s4 ? tmp1254 : 1;
  assign tmp1252 = s5 ? 1 : tmp1253;
  assign tmp1251 = s6 ? tmp1252 : 1;
  assign tmp1250 = s7 ? 1 : tmp1251;
  assign tmp1261 = s2 ? tmp1027 : 1;
  assign tmp1260 = s3 ? tmp1261 : 1;
  assign tmp1259 = s4 ? tmp1260 : 1;
  assign tmp1258 = s5 ? 1 : tmp1259;
  assign tmp1257 = s6 ? 1 : tmp1258;
  assign tmp1256 = s7 ? 1 : tmp1257;
  assign tmp1249 = s8 ? tmp1250 : tmp1256;
  assign tmp1248 = s9 ? 1 : tmp1249;
  assign tmp1265 = s6 ? 1 : tmp1252;
  assign tmp1264 = s7 ? 1 : tmp1265;
  assign tmp1263 = s8 ? tmp1250 : tmp1264;
  assign tmp1262 = s9 ? 1 : tmp1263;
  assign tmp1247 = ~(s10 ? tmp1248 : tmp1262);
  assign tmp1226 = s11 ? tmp1227 : tmp1247;
  assign tmp1275 = s2 ? tmp920 : tmp915;
  assign tmp1274 = s3 ? tmp1275 : tmp915;
  assign tmp1273 = s4 ? tmp945 : tmp1274;
  assign tmp1272 = s5 ? tmp915 : tmp1273;
  assign tmp1271 = s6 ? tmp1272 : tmp934;
  assign tmp1270 = s7 ? tmp933 : tmp1271;
  assign tmp1277 = s6 ? tmp954 : tmp1272;
  assign tmp1276 = s7 ? tmp953 : tmp1277;
  assign tmp1269 = s8 ? tmp1270 : tmp1276;
  assign tmp1268 = s9 ? tmp914 : tmp1269;
  assign tmp1281 = s6 ? tmp914 : tmp1272;
  assign tmp1280 = s7 ? tmp933 : tmp1281;
  assign tmp1279 = s8 ? tmp1270 : tmp1280;
  assign tmp1278 = s9 ? tmp914 : tmp1279;
  assign tmp1267 = s10 ? tmp1268 : tmp1278;
  assign tmp1266 = s11 ? tmp1267 : tmp963;
  assign tmp1225 = s12 ? tmp1226 : tmp1266;
  assign tmp1293 = s1 ? 1 : tmp1023;
  assign tmp1292 = s2 ? tmp1293 : 1;
  assign tmp1294 = s2 ? 1 : tmp929;
  assign tmp1291 = s3 ? tmp1292 : tmp1294;
  assign tmp1290 = s4 ? 1 : tmp1291;
  assign tmp1289 = s5 ? 1 : tmp1290;
  assign tmp1288 = s6 ? tmp1289 : 1;
  assign tmp1287 = s7 ? 1 : tmp1288;
  assign tmp1299 = s3 ? tmp1292 : 1;
  assign tmp1298 = s4 ? 1 : tmp1299;
  assign tmp1297 = s5 ? 1 : tmp1298;
  assign tmp1296 = s6 ? 1 : tmp1297;
  assign tmp1295 = s7 ? 1 : tmp1296;
  assign tmp1286 = s8 ? tmp1287 : tmp1295;
  assign tmp1285 = s9 ? 1 : tmp1286;
  assign tmp1303 = s6 ? 1 : tmp1289;
  assign tmp1302 = s7 ? 1 : tmp1303;
  assign tmp1301 = s8 ? tmp1287 : tmp1302;
  assign tmp1300 = s9 ? 1 : tmp1301;
  assign tmp1284 = s10 ? tmp1285 : tmp1300;
  assign tmp1312 = s2 ? tmp1238 : 1;
  assign tmp1311 = s3 ? 1 : tmp1312;
  assign tmp1313 = s3 ? 1 : tmp985;
  assign tmp1310 = s4 ? tmp1311 : tmp1313;
  assign tmp1309 = s5 ? 1 : tmp1310;
  assign tmp1308 = s6 ? tmp1309 : 1;
  assign tmp1307 = s7 ? 1 : tmp1308;
  assign tmp1317 = s4 ? tmp1311 : 1;
  assign tmp1316 = s5 ? 1 : tmp1317;
  assign tmp1315 = s6 ? 1 : tmp1316;
  assign tmp1314 = s7 ? 1 : tmp1315;
  assign tmp1306 = s8 ? tmp1307 : tmp1314;
  assign tmp1305 = s9 ? 1 : tmp1306;
  assign tmp1321 = s6 ? 1 : tmp1309;
  assign tmp1320 = s7 ? 1 : tmp1321;
  assign tmp1319 = s8 ? tmp1307 : tmp1320;
  assign tmp1318 = s9 ? 1 : tmp1319;
  assign tmp1304 = ~(s10 ? tmp1305 : tmp1318);
  assign tmp1283 = s11 ? tmp1284 : tmp1304;
  assign tmp1332 = ~(s1 ? tmp1133 : tmp915);
  assign tmp1331 = s2 ? tmp951 : tmp1332;
  assign tmp1334 = s1 ? tmp1126 : tmp915;
  assign tmp1333 = ~(s2 ? tmp1334 : tmp915);
  assign tmp1330 = ~(s3 ? tmp1331 : tmp1333);
  assign tmp1329 = s4 ? tmp1130 : tmp1330;
  assign tmp1328 = s5 ? tmp1125 : tmp1329;
  assign tmp1327 = s6 ? tmp1328 : tmp1139;
  assign tmp1326 = s7 ? tmp1108 : tmp1327;
  assign tmp1339 = ~(s3 ? tmp1331 : tmp1138);
  assign tmp1338 = s4 ? tmp1130 : tmp1339;
  assign tmp1337 = s5 ? tmp1125 : tmp1338;
  assign tmp1336 = s6 ? tmp1158 : tmp1337;
  assign tmp1335 = s7 ? tmp1150 : tmp1336;
  assign tmp1325 = s8 ? tmp1326 : tmp1335;
  assign tmp1324 = s9 ? tmp1097 : tmp1325;
  assign tmp1343 = s6 ? tmp1119 : tmp1328;
  assign tmp1342 = s7 ? tmp1163 : tmp1343;
  assign tmp1341 = s8 ? tmp1326 : tmp1342;
  assign tmp1340 = s9 ? tmp1097 : tmp1341;
  assign tmp1323 = s10 ? tmp1324 : tmp1340;
  assign tmp1322 = ~(s11 ? tmp1014 : tmp1323);
  assign tmp1282 = ~(s12 ? tmp1283 : tmp1322);
  assign tmp1224 = s13 ? tmp1225 : tmp1282;
  assign tmp1165 = s15 ? tmp1166 : tmp1224;
  assign tmp907 = s16 ? tmp908 : tmp1165;
  assign l1__1 = tmp907;

  assign tmp1361 = l2 ? 1 : 0;
  assign tmp1360 = l1 ? tmp1361 : 1;
  assign tmp1359 = s0 ? tmp1360 : 0;
  assign tmp1358 = s1 ? tmp1359 : 0;
  assign tmp1357 = ~(s2 ? tmp1358 : 0);
  assign tmp1356 = s3 ? 1 : tmp1357;
  assign tmp1365 = ~(s0 ? tmp1360 : 0);
  assign tmp1364 = s1 ? 1 : tmp1365;
  assign tmp1363 = s2 ? 1 : tmp1364;
  assign tmp1362 = s3 ? tmp1363 : 1;
  assign tmp1355 = s4 ? tmp1356 : tmp1362;
  assign tmp1354 = s5 ? 1 : tmp1355;
  assign tmp1353 = s6 ? tmp1354 : 1;
  assign tmp1352 = s7 ? 1 : tmp1353;
  assign tmp1369 = s4 ? tmp1356 : 1;
  assign tmp1368 = s5 ? 1 : tmp1369;
  assign tmp1367 = s6 ? 1 : tmp1368;
  assign tmp1366 = s7 ? 1 : tmp1367;
  assign tmp1351 = s8 ? tmp1352 : tmp1366;
  assign tmp1350 = s9 ? 1 : tmp1351;
  assign tmp1373 = s6 ? 1 : tmp1354;
  assign tmp1372 = s7 ? 1 : tmp1373;
  assign tmp1371 = s8 ? tmp1352 : tmp1372;
  assign tmp1370 = s9 ? 1 : tmp1371;
  assign tmp1349 = s10 ? tmp1350 : tmp1370;
  assign tmp1385 = ~(l1 ? 1 : tmp1361);
  assign tmp1384 = s0 ? 1 : tmp1385;
  assign tmp1383 = s1 ? 1 : tmp1384;
  assign tmp1386 = s1 ? tmp1384 : 1;
  assign tmp1382 = s2 ? tmp1383 : tmp1386;
  assign tmp1381 = s3 ? tmp1382 : 1;
  assign tmp1380 = s4 ? tmp1381 : 1;
  assign tmp1379 = s5 ? 1 : tmp1380;
  assign tmp1378 = s6 ? tmp1379 : 1;
  assign tmp1377 = s7 ? 1 : tmp1378;
  assign tmp1392 = s2 ? tmp1383 : 1;
  assign tmp1391 = s3 ? tmp1392 : 1;
  assign tmp1390 = s4 ? tmp1391 : 1;
  assign tmp1389 = s5 ? 1 : tmp1390;
  assign tmp1388 = s6 ? 1 : tmp1389;
  assign tmp1387 = s7 ? 1 : tmp1388;
  assign tmp1376 = s8 ? tmp1377 : tmp1387;
  assign tmp1375 = s9 ? 1 : tmp1376;
  assign tmp1396 = s6 ? 1 : tmp1379;
  assign tmp1395 = s7 ? 1 : tmp1396;
  assign tmp1394 = s8 ? tmp1377 : tmp1395;
  assign tmp1393 = s9 ? 1 : tmp1394;
  assign tmp1374 = s10 ? tmp1375 : tmp1393;
  assign tmp1348 = s11 ? tmp1349 : tmp1374;
  assign tmp1408 = s0 ? tmp1361 : 0;
  assign tmp1407 = s1 ? tmp1408 : 0;
  assign tmp1406 = s2 ? tmp1407 : 0;
  assign tmp1410 = ~(l2 ? 1 : 0);
  assign tmp1409 = ~(s2 ? 1 : tmp1410);
  assign tmp1405 = ~(s3 ? tmp1406 : tmp1409);
  assign tmp1404 = s4 ? 1 : tmp1405;
  assign tmp1403 = s5 ? 1 : tmp1404;
  assign tmp1402 = s6 ? tmp1403 : 1;
  assign tmp1401 = s7 ? 1 : tmp1402;
  assign tmp1415 = ~(s3 ? tmp1406 : 0);
  assign tmp1414 = s4 ? 1 : tmp1415;
  assign tmp1413 = s5 ? 1 : tmp1414;
  assign tmp1412 = s6 ? 1 : tmp1413;
  assign tmp1411 = s7 ? 1 : tmp1412;
  assign tmp1400 = s8 ? tmp1401 : tmp1411;
  assign tmp1399 = s9 ? 1 : tmp1400;
  assign tmp1419 = s6 ? 1 : tmp1403;
  assign tmp1418 = s7 ? 1 : tmp1419;
  assign tmp1417 = s8 ? tmp1401 : tmp1418;
  assign tmp1416 = s9 ? 1 : tmp1417;
  assign tmp1398 = s10 ? tmp1399 : tmp1416;
  assign tmp1431 = l1 ? 1 : tmp1410;
  assign tmp1430 = s0 ? tmp1431 : 1;
  assign tmp1429 = s1 ? 1 : tmp1430;
  assign tmp1428 = s2 ? 1 : tmp1429;
  assign tmp1427 = s3 ? 1 : tmp1428;
  assign tmp1432 = s3 ? 1 : tmp1429;
  assign tmp1426 = s4 ? tmp1427 : tmp1432;
  assign tmp1425 = s5 ? 1 : tmp1426;
  assign tmp1424 = s6 ? tmp1425 : 1;
  assign tmp1423 = s7 ? 1 : tmp1424;
  assign tmp1436 = s4 ? tmp1427 : 1;
  assign tmp1435 = s5 ? 1 : tmp1436;
  assign tmp1434 = s6 ? 1 : tmp1435;
  assign tmp1433 = s7 ? 1 : tmp1434;
  assign tmp1422 = s8 ? tmp1423 : tmp1433;
  assign tmp1421 = s9 ? 1 : tmp1422;
  assign tmp1440 = s6 ? 1 : tmp1425;
  assign tmp1439 = s7 ? 1 : tmp1440;
  assign tmp1438 = s8 ? tmp1423 : tmp1439;
  assign tmp1437 = s9 ? 1 : tmp1438;
  assign tmp1420 = s10 ? tmp1421 : tmp1437;
  assign tmp1397 = s11 ? tmp1398 : tmp1420;
  assign tmp1347 = s12 ? tmp1348 : tmp1397;
  assign tmp1454 = l1 ? 1 : tmp1361;
  assign tmp1453 = ~(s0 ? tmp1454 : 0);
  assign tmp1452 = s1 ? 1 : tmp1453;
  assign tmp1451 = s2 ? tmp1452 : 1;
  assign tmp1455 = s2 ? 1 : tmp1385;
  assign tmp1450 = s3 ? tmp1451 : tmp1455;
  assign tmp1449 = s4 ? 1 : tmp1450;
  assign tmp1448 = s5 ? 1 : tmp1449;
  assign tmp1447 = s6 ? tmp1448 : 1;
  assign tmp1446 = s7 ? 1 : tmp1447;
  assign tmp1460 = s3 ? tmp1451 : 1;
  assign tmp1459 = s4 ? 1 : tmp1460;
  assign tmp1458 = s5 ? 1 : tmp1459;
  assign tmp1457 = s6 ? 1 : tmp1458;
  assign tmp1456 = s7 ? 1 : tmp1457;
  assign tmp1445 = s8 ? tmp1446 : tmp1456;
  assign tmp1444 = s9 ? 1 : tmp1445;
  assign tmp1464 = s6 ? 1 : tmp1448;
  assign tmp1463 = s7 ? 1 : tmp1464;
  assign tmp1462 = s8 ? tmp1446 : tmp1463;
  assign tmp1461 = s9 ? 1 : tmp1462;
  assign tmp1443 = s10 ? tmp1444 : tmp1461;
  assign tmp1473 = s2 ? tmp1364 : 1;
  assign tmp1472 = s3 ? 1 : tmp1473;
  assign tmp1475 = ~(s1 ? tmp1359 : 0);
  assign tmp1474 = s3 ? 1 : tmp1475;
  assign tmp1471 = s4 ? tmp1472 : tmp1474;
  assign tmp1470 = s5 ? 1 : tmp1471;
  assign tmp1469 = s6 ? tmp1470 : 1;
  assign tmp1468 = s7 ? 1 : tmp1469;
  assign tmp1479 = s4 ? tmp1472 : 1;
  assign tmp1478 = s5 ? 1 : tmp1479;
  assign tmp1477 = s6 ? 1 : tmp1478;
  assign tmp1476 = s7 ? 1 : tmp1477;
  assign tmp1467 = s8 ? tmp1468 : tmp1476;
  assign tmp1466 = s9 ? 1 : tmp1467;
  assign tmp1483 = s6 ? 1 : tmp1470;
  assign tmp1482 = s7 ? 1 : tmp1483;
  assign tmp1481 = s8 ? tmp1468 : tmp1482;
  assign tmp1480 = s9 ? 1 : tmp1481;
  assign tmp1465 = s10 ? tmp1466 : tmp1480;
  assign tmp1442 = s11 ? tmp1443 : tmp1465;
  assign tmp1496 = l1 ? tmp1361 : 0;
  assign tmp1495 = s0 ? tmp1496 : 0;
  assign tmp1494 = ~(s1 ? tmp1495 : 0);
  assign tmp1493 = s2 ? 1 : tmp1494;
  assign tmp1498 = ~(l1 ? tmp1361 : 0);
  assign tmp1497 = s2 ? 1 : tmp1498;
  assign tmp1492 = s3 ? tmp1493 : tmp1497;
  assign tmp1491 = s4 ? 1 : tmp1492;
  assign tmp1490 = s5 ? 1 : tmp1491;
  assign tmp1489 = s6 ? tmp1490 : 1;
  assign tmp1488 = s7 ? 1 : tmp1489;
  assign tmp1503 = s3 ? tmp1493 : 1;
  assign tmp1502 = s4 ? 1 : tmp1503;
  assign tmp1501 = s5 ? 1 : tmp1502;
  assign tmp1500 = s6 ? 1 : tmp1501;
  assign tmp1499 = s7 ? 1 : tmp1500;
  assign tmp1487 = s8 ? tmp1488 : tmp1499;
  assign tmp1486 = s9 ? 1 : tmp1487;
  assign tmp1507 = s6 ? 1 : tmp1490;
  assign tmp1506 = s7 ? 1 : tmp1507;
  assign tmp1505 = s8 ? tmp1488 : tmp1506;
  assign tmp1504 = s9 ? 1 : tmp1505;
  assign tmp1485 = s10 ? tmp1486 : tmp1504;
  assign tmp1484 = s11 ? 1 : tmp1485;
  assign tmp1441 = s12 ? tmp1442 : tmp1484;
  assign tmp1346 = s13 ? tmp1347 : tmp1441;
  assign tmp1345 = s15 ? 1 : tmp1346;
  assign tmp1344 = ~(s16 ? 1 : tmp1345);
  assign l2__1 = tmp1344;

  assign tmp1516 = l3 ? 1 : 0;
  assign tmp1515 = l1 ? 1 : tmp1516;
  assign tmp1520 = s1 ? tmp1515 : 1;
  assign tmp1521 = s0 ? tmp1515 : 1;
  assign tmp1519 = s2 ? tmp1520 : tmp1521;
  assign tmp1524 = s0 ? 1 : tmp1516;
  assign tmp1523 = s1 ? 1 : tmp1524;
  assign tmp1522 = s2 ? tmp1523 : tmp1515;
  assign tmp1518 = s3 ? tmp1519 : tmp1522;
  assign tmp1528 = s0 ? tmp1515 : 0;
  assign tmp1530 = ~(l1 ? 1 : 0);
  assign tmp1529 = ~(s0 ? 1 : tmp1530);
  assign tmp1527 = s1 ? tmp1528 : tmp1529;
  assign tmp1532 = l1 ? 1 : 0;
  assign tmp1531 = s1 ? tmp1515 : tmp1532;
  assign tmp1526 = s2 ? tmp1527 : tmp1531;
  assign tmp1535 = s0 ? 1 : tmp1515;
  assign tmp1534 = s1 ? tmp1535 : tmp1515;
  assign tmp1533 = s2 ? tmp1534 : tmp1528;
  assign tmp1525 = s3 ? tmp1526 : tmp1533;
  assign tmp1517 = s4 ? tmp1518 : tmp1525;
  assign tmp1514 = s5 ? tmp1515 : tmp1517;
  assign tmp1544 = s0 ? tmp1516 : 1;
  assign tmp1543 = s1 ? tmp1544 : tmp1515;
  assign tmp1542 = s2 ? tmp1523 : tmp1543;
  assign tmp1541 = s3 ? tmp1519 : tmp1542;
  assign tmp1548 = s0 ? tmp1532 : tmp1515;
  assign tmp1547 = s1 ? tmp1548 : tmp1532;
  assign tmp1546 = s2 ? tmp1527 : tmp1547;
  assign tmp1551 = s0 ? tmp1516 : tmp1532;
  assign tmp1550 = s1 ? tmp1528 : tmp1551;
  assign tmp1549 = s2 ? tmp1534 : tmp1550;
  assign tmp1545 = s3 ? tmp1546 : tmp1549;
  assign tmp1540 = s4 ? tmp1541 : tmp1545;
  assign tmp1539 = s5 ? tmp1515 : tmp1540;
  assign tmp1538 = s6 ? tmp1539 : tmp1514;
  assign tmp1557 = s1 ? tmp1515 : tmp1521;
  assign tmp1556 = s2 ? tmp1520 : tmp1557;
  assign tmp1559 = s1 ? 1 : tmp1516;
  assign tmp1560 = s1 ? 1 : tmp1515;
  assign tmp1558 = s2 ? tmp1559 : tmp1560;
  assign tmp1555 = s3 ? tmp1556 : tmp1558;
  assign tmp1563 = s1 ? 1 : tmp1530;
  assign tmp1564 = ~(s1 ? tmp1515 : tmp1532);
  assign tmp1562 = s2 ? tmp1563 : tmp1564;
  assign tmp1565 = ~(l1 ? 1 : tmp1516);
  assign tmp1561 = ~(s3 ? tmp1562 : tmp1565);
  assign tmp1554 = s4 ? tmp1555 : tmp1561;
  assign tmp1553 = s5 ? tmp1515 : tmp1554;
  assign tmp1570 = s1 ? tmp1544 : tmp1535;
  assign tmp1569 = s2 ? tmp1523 : tmp1570;
  assign tmp1568 = s3 ? tmp1519 : tmp1569;
  assign tmp1574 = s0 ? 1 : tmp1532;
  assign tmp1573 = s1 ? tmp1548 : tmp1574;
  assign tmp1572 = s2 ? tmp1527 : tmp1573;
  assign tmp1575 = s2 ? tmp1535 : tmp1550;
  assign tmp1571 = s3 ? tmp1572 : tmp1575;
  assign tmp1567 = s4 ? tmp1568 : tmp1571;
  assign tmp1566 = s5 ? tmp1515 : tmp1567;
  assign tmp1552 = s6 ? tmp1553 : tmp1566;
  assign tmp1537 = s7 ? tmp1538 : tmp1552;
  assign tmp1580 = s3 ? tmp1556 : tmp1522;
  assign tmp1581 = s3 ? tmp1526 : tmp1515;
  assign tmp1579 = s4 ? tmp1580 : tmp1581;
  assign tmp1578 = s5 ? tmp1515 : tmp1579;
  assign tmp1577 = s6 ? tmp1539 : tmp1578;
  assign tmp1582 = s6 ? tmp1578 : tmp1553;
  assign tmp1576 = s7 ? tmp1577 : tmp1582;
  assign tmp1536 = s8 ? tmp1537 : tmp1576;
  assign tmp1513 = s9 ? tmp1514 : tmp1536;
  assign tmp1586 = s6 ? tmp1514 : tmp1553;
  assign tmp1585 = s7 ? tmp1538 : tmp1586;
  assign tmp1584 = s8 ? tmp1537 : tmp1585;
  assign tmp1583 = s9 ? tmp1514 : tmp1584;
  assign tmp1512 = s10 ? tmp1513 : tmp1583;
  assign tmp1590 = l1 ? tmp1516 : 1;
  assign tmp1594 = s1 ? tmp1590 : 1;
  assign tmp1595 = s0 ? tmp1590 : 1;
  assign tmp1593 = s2 ? tmp1594 : tmp1595;
  assign tmp1598 = s0 ? 1 : tmp1530;
  assign tmp1597 = s1 ? 1 : tmp1598;
  assign tmp1596 = s2 ? tmp1597 : tmp1590;
  assign tmp1592 = s3 ? tmp1593 : tmp1596;
  assign tmp1601 = s1 ? tmp1590 : tmp1516;
  assign tmp1600 = s2 ? tmp1516 : tmp1601;
  assign tmp1603 = s0 ? 1 : tmp1590;
  assign tmp1602 = s1 ? tmp1603 : tmp1590;
  assign tmp1599 = s3 ? tmp1600 : tmp1602;
  assign tmp1591 = s4 ? tmp1592 : tmp1599;
  assign tmp1589 = s5 ? tmp1590 : tmp1591;
  assign tmp1613 = ~(l1 ? tmp1516 : 1);
  assign tmp1612 = s0 ? tmp1532 : tmp1613;
  assign tmp1611 = ~(s1 ? tmp1612 : tmp1613);
  assign tmp1610 = s2 ? tmp1597 : tmp1611;
  assign tmp1609 = s3 ? tmp1593 : tmp1610;
  assign tmp1615 = s2 ? tmp1523 : tmp1601;
  assign tmp1619 = ~(l3 ? 1 : 0);
  assign tmp1618 = ~(s0 ? tmp1532 : tmp1619);
  assign tmp1617 = s1 ? 1 : tmp1618;
  assign tmp1616 = s2 ? tmp1602 : tmp1617;
  assign tmp1614 = s3 ? tmp1615 : tmp1616;
  assign tmp1608 = s4 ? tmp1609 : tmp1614;
  assign tmp1607 = s5 ? tmp1590 : tmp1608;
  assign tmp1623 = s2 ? tmp1559 : tmp1601;
  assign tmp1622 = s3 ? tmp1623 : tmp1602;
  assign tmp1621 = s4 ? tmp1592 : tmp1622;
  assign tmp1620 = s5 ? tmp1590 : tmp1621;
  assign tmp1606 = s6 ? tmp1607 : tmp1620;
  assign tmp1629 = s1 ? tmp1590 : tmp1595;
  assign tmp1628 = s2 ? tmp1594 : tmp1629;
  assign tmp1630 = s2 ? tmp1563 : tmp1594;
  assign tmp1627 = s3 ? tmp1628 : tmp1630;
  assign tmp1632 = s2 ? tmp1559 : tmp1590;
  assign tmp1631 = s3 ? tmp1632 : tmp1590;
  assign tmp1626 = s4 ? tmp1627 : tmp1631;
  assign tmp1625 = s5 ? tmp1590 : tmp1626;
  assign tmp1638 = ~(s0 ? tmp1590 : 1);
  assign tmp1637 = ~(s1 ? tmp1612 : tmp1638);
  assign tmp1636 = s2 ? tmp1597 : tmp1637;
  assign tmp1635 = s3 ? tmp1593 : tmp1636;
  assign tmp1641 = s1 ? tmp1590 : tmp1603;
  assign tmp1640 = s2 ? tmp1523 : tmp1641;
  assign tmp1639 = s3 ? tmp1640 : tmp1616;
  assign tmp1634 = s4 ? tmp1635 : tmp1639;
  assign tmp1633 = s5 ? tmp1590 : tmp1634;
  assign tmp1624 = s6 ? tmp1625 : tmp1633;
  assign tmp1605 = s7 ? tmp1606 : tmp1624;
  assign tmp1646 = s3 ? tmp1623 : tmp1616;
  assign tmp1645 = s4 ? tmp1609 : tmp1646;
  assign tmp1644 = s5 ? tmp1590 : tmp1645;
  assign tmp1649 = s3 ? tmp1628 : tmp1596;
  assign tmp1651 = s2 ? tmp1516 : tmp1590;
  assign tmp1650 = s3 ? tmp1651 : tmp1590;
  assign tmp1648 = s4 ? tmp1649 : tmp1650;
  assign tmp1647 = s5 ? tmp1590 : tmp1648;
  assign tmp1643 = s6 ? tmp1644 : tmp1647;
  assign tmp1654 = s4 ? tmp1649 : tmp1631;
  assign tmp1653 = s5 ? tmp1590 : tmp1654;
  assign tmp1652 = s6 ? tmp1653 : tmp1625;
  assign tmp1642 = s7 ? tmp1643 : tmp1652;
  assign tmp1604 = s8 ? tmp1605 : tmp1642;
  assign tmp1588 = s9 ? tmp1589 : tmp1604;
  assign tmp1658 = s6 ? tmp1644 : tmp1589;
  assign tmp1659 = s6 ? tmp1620 : tmp1625;
  assign tmp1657 = s7 ? tmp1658 : tmp1659;
  assign tmp1656 = s8 ? tmp1605 : tmp1657;
  assign tmp1655 = s9 ? tmp1589 : tmp1656;
  assign tmp1587 = s10 ? tmp1588 : tmp1655;
  assign tmp1511 = s11 ? tmp1512 : tmp1587;
  assign tmp1510 = s12 ? 1 : tmp1511;
  assign tmp1661 = s11 ? 1 : 0;
  assign tmp1666 = l1 ? 1 : tmp1619;
  assign tmp1670 = s1 ? 1 : tmp1666;
  assign tmp1671 = s1 ? tmp1666 : tmp1619;
  assign tmp1669 = s2 ? tmp1670 : tmp1671;
  assign tmp1668 = s3 ? tmp1666 : tmp1669;
  assign tmp1674 = s1 ? tmp1666 : 1;
  assign tmp1673 = s2 ? 1 : tmp1674;
  assign tmp1675 = s2 ? tmp1666 : tmp1670;
  assign tmp1672 = s3 ? tmp1673 : tmp1675;
  assign tmp1667 = s4 ? tmp1668 : tmp1672;
  assign tmp1665 = s5 ? tmp1666 : tmp1667;
  assign tmp1684 = s0 ? tmp1666 : 0;
  assign tmp1683 = s1 ? tmp1666 : tmp1684;
  assign tmp1682 = s2 ? tmp1666 : tmp1683;
  assign tmp1687 = s0 ? 1 : 0;
  assign tmp1688 = ~(s0 ? 1 : tmp1666);
  assign tmp1686 = s1 ? tmp1687 : tmp1688;
  assign tmp1689 = ~(l1 ? 1 : tmp1619);
  assign tmp1685 = ~(s2 ? tmp1686 : tmp1689);
  assign tmp1681 = s3 ? tmp1682 : tmp1685;
  assign tmp1693 = s0 ? tmp1516 : 0;
  assign tmp1692 = s1 ? tmp1693 : 0;
  assign tmp1695 = s0 ? 1 : tmp1666;
  assign tmp1696 = ~(s0 ? 1 : 0);
  assign tmp1694 = ~(s1 ? tmp1695 : tmp1696);
  assign tmp1691 = s2 ? tmp1692 : tmp1694;
  assign tmp1698 = s1 ? tmp1695 : tmp1666;
  assign tmp1699 = s0 ? tmp1666 : 1;
  assign tmp1697 = ~(s2 ? tmp1698 : tmp1699);
  assign tmp1690 = ~(s3 ? tmp1691 : tmp1697);
  assign tmp1680 = s4 ? tmp1681 : tmp1690;
  assign tmp1679 = s5 ? tmp1666 : tmp1680;
  assign tmp1702 = s3 ? tmp1682 : tmp1669;
  assign tmp1701 = s4 ? tmp1702 : tmp1672;
  assign tmp1700 = s5 ? tmp1666 : tmp1701;
  assign tmp1678 = s6 ? tmp1679 : tmp1700;
  assign tmp1707 = ~(s0 ? tmp1516 : tmp1689);
  assign tmp1706 = s1 ? tmp1666 : tmp1707;
  assign tmp1705 = s2 ? tmp1666 : tmp1706;
  assign tmp1711 = s1 ? tmp1666 : 0;
  assign tmp1710 = s2 ? tmp1711 : tmp1683;
  assign tmp1714 = s0 ? tmp1666 : tmp1532;
  assign tmp1713 = s1 ? tmp1714 : tmp1619;
  assign tmp1712 = s2 ? tmp1670 : tmp1713;
  assign tmp1709 = s3 ? tmp1710 : tmp1712;
  assign tmp1715 = s3 ? tmp1673 : tmp1666;
  assign tmp1708 = s4 ? tmp1709 : tmp1715;
  assign tmp1704 = s5 ? tmp1705 : tmp1708;
  assign tmp1721 = s0 ? tmp1532 : tmp1619;
  assign tmp1720 = ~(s1 ? tmp1714 : tmp1721);
  assign tmp1719 = ~(s2 ? tmp1686 : tmp1720);
  assign tmp1718 = s3 ? tmp1710 : tmp1719;
  assign tmp1725 = s0 ? tmp1532 : tmp1666;
  assign tmp1724 = s1 ? tmp1695 : tmp1725;
  assign tmp1723 = ~(s2 ? tmp1724 : tmp1699);
  assign tmp1722 = ~(s3 ? tmp1691 : tmp1723);
  assign tmp1717 = s4 ? tmp1718 : tmp1722;
  assign tmp1716 = s5 ? tmp1705 : tmp1717;
  assign tmp1703 = s6 ? tmp1704 : tmp1716;
  assign tmp1677 = s7 ? tmp1678 : tmp1703;
  assign tmp1732 = s1 ? 1 : tmp1695;
  assign tmp1731 = s2 ? tmp1732 : tmp1666;
  assign tmp1730 = s3 ? tmp1666 : tmp1731;
  assign tmp1735 = ~(s1 ? tmp1695 : 1);
  assign tmp1734 = s2 ? tmp1692 : tmp1735;
  assign tmp1733 = ~(s3 ? tmp1734 : tmp1697);
  assign tmp1729 = s4 ? tmp1730 : tmp1733;
  assign tmp1728 = s5 ? tmp1666 : tmp1729;
  assign tmp1739 = s2 ? tmp1666 : tmp1699;
  assign tmp1738 = s3 ? tmp1739 : tmp1669;
  assign tmp1737 = s4 ? tmp1738 : tmp1715;
  assign tmp1736 = s5 ? tmp1666 : tmp1737;
  assign tmp1727 = s6 ? tmp1728 : tmp1736;
  assign tmp1742 = s4 ? tmp1702 : tmp1715;
  assign tmp1741 = s5 ? tmp1666 : tmp1742;
  assign tmp1740 = s6 ? tmp1741 : tmp1704;
  assign tmp1726 = s7 ? tmp1727 : tmp1740;
  assign tmp1676 = s8 ? tmp1677 : tmp1726;
  assign tmp1664 = s9 ? tmp1665 : tmp1676;
  assign tmp1746 = s6 ? tmp1728 : tmp1665;
  assign tmp1747 = s6 ? tmp1700 : tmp1704;
  assign tmp1745 = s7 ? tmp1746 : tmp1747;
  assign tmp1744 = s8 ? tmp1677 : tmp1745;
  assign tmp1743 = s9 ? tmp1665 : tmp1744;
  assign tmp1663 = s10 ? tmp1664 : tmp1743;
  assign tmp1751 = l1 ? tmp1516 : 0;
  assign tmp1755 = s1 ? tmp1751 : 0;
  assign tmp1754 = s2 ? tmp1755 : tmp1751;
  assign tmp1757 = s1 ? 1 : tmp1687;
  assign tmp1756 = s2 ? tmp1757 : tmp1751;
  assign tmp1753 = s3 ? tmp1754 : tmp1756;
  assign tmp1762 = ~(l1 ? tmp1516 : 0);
  assign tmp1761 = s0 ? 1 : tmp1762;
  assign tmp1760 = s1 ? 1 : tmp1761;
  assign tmp1759 = s2 ? tmp1760 : tmp1762;
  assign tmp1764 = ~(s1 ? 1 : tmp1762);
  assign tmp1763 = ~(s2 ? tmp1751 : tmp1764);
  assign tmp1758 = ~(s3 ? tmp1759 : tmp1763);
  assign tmp1752 = s4 ? tmp1753 : tmp1758;
  assign tmp1750 = s5 ? tmp1751 : tmp1752;
  assign tmp1772 = s1 ? tmp1751 : 1;
  assign tmp1774 = s0 ? tmp1751 : 1;
  assign tmp1773 = s1 ? tmp1774 : tmp1751;
  assign tmp1771 = s2 ? tmp1772 : tmp1773;
  assign tmp1777 = s0 ? 1 : tmp1619;
  assign tmp1776 = ~(s1 ? tmp1777 : tmp1762);
  assign tmp1775 = s2 ? tmp1757 : tmp1776;
  assign tmp1770 = s3 ? tmp1771 : tmp1775;
  assign tmp1781 = s0 ? tmp1532 : 0;
  assign tmp1782 = ~(s0 ? 1 : tmp1762);
  assign tmp1780 = s1 ? tmp1781 : tmp1782;
  assign tmp1779 = s2 ? tmp1780 : tmp1751;
  assign tmp1783 = s2 ? tmp1751 : tmp1780;
  assign tmp1778 = s3 ? tmp1779 : tmp1783;
  assign tmp1769 = s4 ? tmp1770 : tmp1778;
  assign tmp1768 = s5 ? tmp1751 : tmp1769;
  assign tmp1787 = s2 ? tmp1772 : tmp1751;
  assign tmp1786 = s3 ? tmp1787 : tmp1756;
  assign tmp1785 = s4 ? tmp1786 : tmp1758;
  assign tmp1784 = s5 ? tmp1751 : tmp1785;
  assign tmp1767 = s6 ? tmp1768 : tmp1784;
  assign tmp1792 = l2 ? 1 : 0;
  assign tmp1791 = l1 ? tmp1516 : tmp1792;
  assign tmp1793 = s0 ? tmp1791 : tmp1751;
  assign tmp1790 = s2 ? tmp1791 : tmp1793;
  assign tmp1798 = s0 ? tmp1532 : tmp1791;
  assign tmp1797 = s1 ? tmp1798 : 1;
  assign tmp1800 = s0 ? tmp1791 : 1;
  assign tmp1799 = s1 ? tmp1791 : tmp1800;
  assign tmp1796 = s2 ? tmp1797 : tmp1799;
  assign tmp1802 = s1 ? 1 : 0;
  assign tmp1803 = s1 ? tmp1516 : tmp1532;
  assign tmp1801 = s2 ? tmp1802 : tmp1803;
  assign tmp1795 = s3 ? tmp1796 : tmp1801;
  assign tmp1806 = s1 ? 1 : tmp1762;
  assign tmp1807 = ~(s1 ? tmp1791 : tmp1751);
  assign tmp1805 = s2 ? tmp1806 : tmp1807;
  assign tmp1804 = ~(s3 ? tmp1805 : tmp1762);
  assign tmp1794 = s4 ? tmp1795 : tmp1804;
  assign tmp1789 = s5 ? tmp1790 : tmp1794;
  assign tmp1811 = s2 ? tmp1797 : tmp1800;
  assign tmp1814 = ~(s0 ? tmp1516 : tmp1532);
  assign tmp1813 = ~(s1 ? tmp1777 : tmp1814);
  assign tmp1812 = s2 ? tmp1757 : tmp1813;
  assign tmp1810 = s3 ? tmp1811 : tmp1812;
  assign tmp1818 = s0 ? tmp1751 : tmp1791;
  assign tmp1819 = s0 ? 1 : tmp1751;
  assign tmp1817 = s1 ? tmp1818 : tmp1819;
  assign tmp1816 = s2 ? tmp1780 : tmp1817;
  assign tmp1822 = s0 ? tmp1516 : tmp1751;
  assign tmp1821 = s1 ? tmp1819 : tmp1822;
  assign tmp1820 = s2 ? tmp1821 : tmp1780;
  assign tmp1815 = s3 ? tmp1816 : tmp1820;
  assign tmp1809 = s4 ? tmp1810 : tmp1815;
  assign tmp1808 = s5 ? tmp1790 : tmp1809;
  assign tmp1788 = s6 ? tmp1789 : tmp1808;
  assign tmp1766 = s7 ? tmp1767 : tmp1788;
  assign tmp1830 = s0 ? tmp1751 : 0;
  assign tmp1829 = s1 ? tmp1830 : tmp1751;
  assign tmp1828 = s2 ? tmp1755 : tmp1829;
  assign tmp1827 = s3 ? tmp1828 : tmp1775;
  assign tmp1826 = s4 ? tmp1827 : tmp1778;
  assign tmp1825 = s5 ? tmp1751 : tmp1826;
  assign tmp1833 = ~(s3 ? tmp1759 : tmp1762);
  assign tmp1832 = s4 ? tmp1753 : tmp1833;
  assign tmp1831 = s5 ? tmp1751 : tmp1832;
  assign tmp1824 = s6 ? tmp1825 : tmp1831;
  assign tmp1836 = s4 ? tmp1786 : tmp1833;
  assign tmp1835 = s5 ? tmp1751 : tmp1836;
  assign tmp1834 = s6 ? tmp1835 : tmp1789;
  assign tmp1823 = s7 ? tmp1824 : tmp1834;
  assign tmp1765 = s8 ? tmp1766 : tmp1823;
  assign tmp1749 = s9 ? tmp1750 : tmp1765;
  assign tmp1840 = s6 ? tmp1825 : tmp1750;
  assign tmp1841 = s6 ? tmp1784 : tmp1789;
  assign tmp1839 = s7 ? tmp1840 : tmp1841;
  assign tmp1838 = s8 ? tmp1766 : tmp1839;
  assign tmp1837 = s9 ? tmp1750 : tmp1838;
  assign tmp1748 = ~(s10 ? tmp1749 : tmp1837);
  assign tmp1662 = s11 ? tmp1663 : tmp1748;
  assign tmp1660 = ~(s12 ? tmp1661 : tmp1662);
  assign tmp1509 = s13 ? tmp1510 : tmp1660;
  assign tmp1854 = s2 ? tmp1802 : 0;
  assign tmp1853 = ~(s3 ? tmp1854 : 0);
  assign tmp1852 = s4 ? 1 : tmp1853;
  assign tmp1851 = s5 ? 1 : tmp1852;
  assign tmp1859 = s1 ? tmp1687 : tmp1696;
  assign tmp1858 = s2 ? tmp1859 : 1;
  assign tmp1860 = s2 ? 1 : tmp1687;
  assign tmp1857 = s3 ? tmp1858 : tmp1860;
  assign tmp1856 = s4 ? 1 : tmp1857;
  assign tmp1855 = s5 ? 1 : tmp1856;
  assign tmp1850 = s6 ? tmp1851 : tmp1855;
  assign tmp1849 = s7 ? tmp1538 : tmp1850;
  assign tmp1862 = s6 ? tmp1578 : tmp1851;
  assign tmp1861 = s7 ? 1 : tmp1862;
  assign tmp1848 = s8 ? tmp1849 : tmp1861;
  assign tmp1847 = s9 ? 1 : tmp1848;
  assign tmp1866 = s6 ? tmp1514 : tmp1851;
  assign tmp1865 = s7 ? 1 : tmp1866;
  assign tmp1864 = s8 ? tmp1849 : tmp1865;
  assign tmp1863 = s9 ? 1 : tmp1864;
  assign tmp1846 = s10 ? tmp1847 : tmp1863;
  assign tmp1874 = l1 ? tmp1792 : 1;
  assign tmp1876 = s0 ? tmp1874 : tmp1792;
  assign tmp1875 = s1 ? tmp1876 : tmp1874;
  assign tmp1873 = s2 ? tmp1874 : tmp1875;
  assign tmp1880 = s1 ? tmp1874 : 1;
  assign tmp1882 = s0 ? tmp1874 : 1;
  assign tmp1881 = s1 ? tmp1874 : tmp1882;
  assign tmp1879 = s2 ? tmp1880 : tmp1881;
  assign tmp1884 = ~(s1 ? 1 : 0);
  assign tmp1883 = s2 ? tmp1802 : tmp1884;
  assign tmp1878 = s3 ? tmp1879 : tmp1883;
  assign tmp1887 = s1 ? tmp1874 : tmp1530;
  assign tmp1886 = s2 ? tmp1802 : tmp1887;
  assign tmp1889 = ~(l1 ? tmp1792 : 1);
  assign tmp1888 = ~(s1 ? 1 : tmp1889);
  assign tmp1885 = s3 ? tmp1886 : tmp1888;
  assign tmp1877 = s4 ? tmp1878 : tmp1885;
  assign tmp1872 = s5 ? tmp1873 : tmp1877;
  assign tmp1893 = s2 ? tmp1880 : tmp1882;
  assign tmp1895 = ~(s1 ? 1 : tmp1687);
  assign tmp1894 = s2 ? tmp1757 : tmp1895;
  assign tmp1892 = s3 ? tmp1893 : tmp1894;
  assign tmp1899 = s0 ? 1 : tmp1889;
  assign tmp1898 = ~(s1 ? tmp1899 : tmp1529);
  assign tmp1897 = s2 ? tmp1757 : tmp1898;
  assign tmp1902 = ~(s0 ? 1 : tmp1889);
  assign tmp1901 = s1 ? tmp1687 : tmp1902;
  assign tmp1900 = s2 ? tmp1901 : tmp1802;
  assign tmp1896 = s3 ? tmp1897 : tmp1900;
  assign tmp1891 = s4 ? tmp1892 : tmp1896;
  assign tmp1890 = s5 ? tmp1873 : tmp1891;
  assign tmp1871 = s6 ? tmp1872 : tmp1890;
  assign tmp1870 = s7 ? tmp1606 : tmp1871;
  assign tmp1904 = ~(s6 ? tmp1653 : tmp1872);
  assign tmp1903 = ~(s7 ? 1 : tmp1904);
  assign tmp1869 = ~(s8 ? tmp1870 : tmp1903);
  assign tmp1868 = s9 ? 1 : tmp1869;
  assign tmp1908 = ~(s6 ? tmp1620 : tmp1872);
  assign tmp1907 = ~(s7 ? 1 : tmp1908);
  assign tmp1906 = ~(s8 ? tmp1870 : tmp1907);
  assign tmp1905 = s9 ? 1 : tmp1906;
  assign tmp1867 = ~(s10 ? tmp1868 : tmp1905);
  assign tmp1845 = s11 ? tmp1846 : tmp1867;
  assign tmp1844 = s12 ? 1 : tmp1845;
  assign tmp1918 = s1 ? tmp1532 : tmp1696;
  assign tmp1917 = s2 ? tmp1532 : tmp1918;
  assign tmp1922 = s1 ? tmp1574 : 0;
  assign tmp1921 = s2 ? tmp1922 : tmp1532;
  assign tmp1920 = s3 ? tmp1921 : 1;
  assign tmp1925 = s1 ? tmp1532 : 1;
  assign tmp1924 = s2 ? 1 : tmp1925;
  assign tmp1923 = s3 ? tmp1924 : tmp1925;
  assign tmp1919 = s4 ? tmp1920 : tmp1923;
  assign tmp1916 = s5 ? tmp1917 : tmp1919;
  assign tmp1930 = s1 ? tmp1687 : 0;
  assign tmp1929 = ~(s2 ? tmp1930 : 0);
  assign tmp1928 = s3 ? tmp1921 : tmp1929;
  assign tmp1933 = s1 ? tmp1574 : tmp1696;
  assign tmp1932 = s2 ? 1 : tmp1933;
  assign tmp1936 = s0 ? tmp1532 : 1;
  assign tmp1935 = s1 ? 1 : tmp1936;
  assign tmp1934 = s2 ? tmp1935 : 1;
  assign tmp1931 = s3 ? tmp1932 : tmp1934;
  assign tmp1927 = s4 ? tmp1928 : tmp1931;
  assign tmp1926 = s5 ? tmp1917 : tmp1927;
  assign tmp1915 = s6 ? tmp1916 : tmp1926;
  assign tmp1914 = s7 ? tmp1678 : tmp1915;
  assign tmp1938 = s6 ? tmp1741 : tmp1916;
  assign tmp1937 = s7 ? 1 : tmp1938;
  assign tmp1913 = s8 ? tmp1914 : tmp1937;
  assign tmp1912 = s9 ? 1 : tmp1913;
  assign tmp1942 = s6 ? tmp1700 : tmp1916;
  assign tmp1941 = s7 ? 1 : tmp1942;
  assign tmp1940 = s8 ? tmp1914 : tmp1941;
  assign tmp1939 = s9 ? 1 : tmp1940;
  assign tmp1911 = s10 ? tmp1912 : tmp1939;
  assign tmp1946 = s7 ? tmp1767 : tmp1871;
  assign tmp1948 = ~(s6 ? tmp1835 : tmp1872);
  assign tmp1947 = ~(s7 ? 1 : tmp1948);
  assign tmp1945 = ~(s8 ? tmp1946 : tmp1947);
  assign tmp1944 = s9 ? 1 : tmp1945;
  assign tmp1952 = ~(s6 ? tmp1784 : tmp1872);
  assign tmp1951 = ~(s7 ? 1 : tmp1952);
  assign tmp1950 = ~(s8 ? tmp1946 : tmp1951);
  assign tmp1949 = s9 ? 1 : tmp1950;
  assign tmp1943 = s10 ? tmp1944 : tmp1949;
  assign tmp1910 = s11 ? tmp1911 : tmp1943;
  assign tmp1909 = ~(s12 ? tmp1661 : tmp1910);
  assign tmp1843 = s13 ? tmp1844 : tmp1909;
  assign tmp1968 = ~(l2 ? 1 : tmp1619);
  assign tmp1967 = l1 ? 1 : tmp1968;
  assign tmp1966 = s0 ? tmp1967 : 0;
  assign tmp1965 = s1 ? tmp1966 : tmp1532;
  assign tmp1964 = s2 ? tmp1965 : tmp1531;
  assign tmp1969 = s2 ? tmp1515 : tmp1967;
  assign tmp1963 = s3 ? tmp1964 : tmp1969;
  assign tmp1962 = s4 ? tmp1555 : tmp1963;
  assign tmp1961 = s5 ? tmp1515 : tmp1962;
  assign tmp1960 = s6 ? tmp1961 : tmp1566;
  assign tmp1959 = s7 ? tmp1538 : tmp1960;
  assign tmp1974 = s3 ? tmp1964 : tmp1515;
  assign tmp1973 = s4 ? tmp1555 : tmp1974;
  assign tmp1972 = s5 ? tmp1515 : tmp1973;
  assign tmp1971 = s6 ? tmp1578 : tmp1972;
  assign tmp1970 = s7 ? tmp1577 : tmp1971;
  assign tmp1958 = s8 ? tmp1959 : tmp1970;
  assign tmp1957 = s9 ? tmp1514 : tmp1958;
  assign tmp1978 = s6 ? tmp1514 : tmp1961;
  assign tmp1977 = s7 ? tmp1538 : tmp1978;
  assign tmp1976 = s8 ? tmp1959 : tmp1977;
  assign tmp1975 = s9 ? tmp1514 : tmp1976;
  assign tmp1956 = s10 ? tmp1957 : tmp1975;
  assign tmp1987 = s2 ? tmp1563 : tmp1629;
  assign tmp1986 = s3 ? tmp1628 : tmp1987;
  assign tmp1985 = s4 ? tmp1986 : tmp1631;
  assign tmp1984 = s5 ? tmp1590 : tmp1985;
  assign tmp1983 = s6 ? tmp1984 : tmp1633;
  assign tmp1982 = s7 ? tmp1606 : tmp1983;
  assign tmp1989 = s6 ? tmp1653 : tmp1984;
  assign tmp1988 = s7 ? tmp1643 : tmp1989;
  assign tmp1981 = s8 ? tmp1982 : tmp1988;
  assign tmp1980 = s9 ? tmp1589 : tmp1981;
  assign tmp1993 = s6 ? tmp1620 : tmp1984;
  assign tmp1992 = s7 ? tmp1658 : tmp1993;
  assign tmp1991 = s8 ? tmp1982 : tmp1992;
  assign tmp1990 = s9 ? tmp1589 : tmp1991;
  assign tmp1979 = s10 ? tmp1980 : tmp1990;
  assign tmp1955 = s11 ? tmp1956 : tmp1979;
  assign tmp1954 = s12 ? 1 : tmp1955;
  assign tmp2006 = ~(s0 ? tmp1874 : 0);
  assign tmp2005 = s1 ? 1 : tmp2006;
  assign tmp2004 = s2 ? tmp2005 : 1;
  assign tmp2003 = s3 ? 1 : tmp2004;
  assign tmp2009 = s0 ? tmp1874 : 0;
  assign tmp2008 = ~(s1 ? tmp2009 : 0);
  assign tmp2007 = s3 ? 1 : tmp2008;
  assign tmp2002 = s4 ? tmp2003 : tmp2007;
  assign tmp2001 = s5 ? 1 : tmp2002;
  assign tmp2000 = s6 ? tmp2001 : 1;
  assign tmp1999 = s7 ? 1 : tmp2000;
  assign tmp2013 = s4 ? tmp2003 : 1;
  assign tmp2012 = s5 ? 1 : tmp2013;
  assign tmp2011 = s6 ? 1 : tmp2012;
  assign tmp2010 = s7 ? 1 : tmp2011;
  assign tmp1998 = s8 ? tmp1999 : tmp2010;
  assign tmp1997 = s9 ? 1 : tmp1998;
  assign tmp2017 = s6 ? 1 : tmp2001;
  assign tmp2016 = s7 ? 1 : tmp2017;
  assign tmp2015 = s8 ? tmp1999 : tmp2016;
  assign tmp2014 = s9 ? 1 : tmp2015;
  assign tmp1996 = ~(s10 ? tmp1997 : tmp2014);
  assign tmp1995 = s11 ? 1 : tmp1996;
  assign tmp2031 = l2 ? 1 : tmp1619;
  assign tmp2030 = l1 ? tmp2031 : 1;
  assign tmp2032 = ~(l1 ? tmp1516 : tmp1792);
  assign tmp2029 = s0 ? tmp2030 : tmp2032;
  assign tmp2028 = s1 ? tmp2029 : tmp1762;
  assign tmp2027 = s2 ? tmp1806 : tmp2028;
  assign tmp2034 = ~(l1 ? tmp2031 : 1);
  assign tmp2033 = ~(s2 ? tmp1751 : tmp2034);
  assign tmp2026 = ~(s3 ? tmp2027 : tmp2033);
  assign tmp2025 = s4 ? tmp1795 : tmp2026;
  assign tmp2024 = s5 ? tmp1790 : tmp2025;
  assign tmp2023 = s6 ? tmp2024 : tmp1808;
  assign tmp2022 = s7 ? tmp1767 : tmp2023;
  assign tmp2039 = ~(s3 ? tmp2027 : tmp1762);
  assign tmp2038 = s4 ? tmp1795 : tmp2039;
  assign tmp2037 = s5 ? tmp1790 : tmp2038;
  assign tmp2036 = s6 ? tmp1835 : tmp2037;
  assign tmp2035 = s7 ? tmp1824 : tmp2036;
  assign tmp2021 = s8 ? tmp2022 : tmp2035;
  assign tmp2020 = s9 ? tmp1750 : tmp2021;
  assign tmp2043 = s6 ? tmp1784 : tmp2024;
  assign tmp2042 = s7 ? tmp1840 : tmp2043;
  assign tmp2041 = s8 ? tmp2022 : tmp2042;
  assign tmp2040 = s9 ? tmp1750 : tmp2041;
  assign tmp2019 = ~(s10 ? tmp2020 : tmp2040);
  assign tmp2018 = s11 ? tmp1663 : tmp2019;
  assign tmp1994 = ~(s12 ? tmp1995 : tmp2018);
  assign tmp1953 = s13 ? tmp1954 : tmp1994;
  assign tmp1842 = s15 ? tmp1843 : tmp1953;
  assign tmp1508 = s16 ? tmp1509 : tmp1842;
  assign l3__1 = tmp1508;

  assign tmp2045 = ~(s15 ? 1 : 0);
  assign tmp2044 = ~(s16 ? 1 : tmp2045);
  assign s16n = tmp2044;

  assign tmp2063 = l2 ? 1 : 0;
  assign tmp2062 = l1 ? tmp2063 : 1;
  assign tmp2061 = s0 ? tmp2062 : 0;
  assign tmp2060 = s1 ? tmp2061 : 0;
  assign tmp2059 = ~(s2 ? tmp2060 : 0);
  assign tmp2058 = s3 ? 1 : tmp2059;
  assign tmp2067 = ~(s0 ? tmp2062 : 0);
  assign tmp2066 = s1 ? 1 : tmp2067;
  assign tmp2065 = s2 ? 1 : tmp2066;
  assign tmp2064 = s3 ? tmp2065 : 1;
  assign tmp2057 = s4 ? tmp2058 : tmp2064;
  assign tmp2056 = s5 ? 1 : tmp2057;
  assign tmp2055 = s6 ? tmp2056 : 1;
  assign tmp2054 = s7 ? 1 : tmp2055;
  assign tmp2071 = s4 ? tmp2058 : 1;
  assign tmp2070 = s5 ? 1 : tmp2071;
  assign tmp2069 = s6 ? 1 : tmp2070;
  assign tmp2068 = s7 ? 1 : tmp2069;
  assign tmp2053 = s8 ? tmp2054 : tmp2068;
  assign tmp2052 = s9 ? 1 : tmp2053;
  assign tmp2075 = s6 ? 1 : tmp2056;
  assign tmp2074 = s7 ? 1 : tmp2075;
  assign tmp2073 = s8 ? tmp2054 : tmp2074;
  assign tmp2072 = s9 ? 1 : tmp2073;
  assign tmp2051 = s10 ? tmp2052 : tmp2072;
  assign tmp2087 = ~(l1 ? 1 : tmp2063);
  assign tmp2086 = s0 ? 1 : tmp2087;
  assign tmp2085 = s1 ? 1 : tmp2086;
  assign tmp2088 = s1 ? tmp2086 : 1;
  assign tmp2084 = s2 ? tmp2085 : tmp2088;
  assign tmp2083 = s3 ? tmp2084 : 1;
  assign tmp2082 = s4 ? tmp2083 : 1;
  assign tmp2081 = s5 ? 1 : tmp2082;
  assign tmp2080 = s6 ? tmp2081 : 1;
  assign tmp2079 = s7 ? 1 : tmp2080;
  assign tmp2094 = s2 ? tmp2085 : 1;
  assign tmp2093 = s3 ? tmp2094 : 1;
  assign tmp2092 = s4 ? tmp2093 : 1;
  assign tmp2091 = s5 ? 1 : tmp2092;
  assign tmp2090 = s6 ? 1 : tmp2091;
  assign tmp2089 = s7 ? 1 : tmp2090;
  assign tmp2078 = s8 ? tmp2079 : tmp2089;
  assign tmp2077 = s9 ? 1 : tmp2078;
  assign tmp2098 = s6 ? 1 : tmp2081;
  assign tmp2097 = s7 ? 1 : tmp2098;
  assign tmp2096 = s8 ? tmp2079 : tmp2097;
  assign tmp2095 = s9 ? 1 : tmp2096;
  assign tmp2076 = s10 ? tmp2077 : tmp2095;
  assign tmp2050 = s11 ? tmp2051 : tmp2076;
  assign tmp2110 = s0 ? tmp2063 : 0;
  assign tmp2109 = s1 ? tmp2110 : 0;
  assign tmp2108 = s2 ? tmp2109 : 0;
  assign tmp2112 = ~(l2 ? 1 : 0);
  assign tmp2111 = ~(s2 ? 1 : tmp2112);
  assign tmp2107 = ~(s3 ? tmp2108 : tmp2111);
  assign tmp2106 = s4 ? 1 : tmp2107;
  assign tmp2105 = s5 ? 1 : tmp2106;
  assign tmp2104 = s6 ? tmp2105 : 1;
  assign tmp2103 = s7 ? 1 : tmp2104;
  assign tmp2117 = ~(s3 ? tmp2108 : 0);
  assign tmp2116 = s4 ? 1 : tmp2117;
  assign tmp2115 = s5 ? 1 : tmp2116;
  assign tmp2114 = s6 ? 1 : tmp2115;
  assign tmp2113 = s7 ? 1 : tmp2114;
  assign tmp2102 = s8 ? tmp2103 : tmp2113;
  assign tmp2101 = s9 ? 1 : tmp2102;
  assign tmp2121 = s6 ? 1 : tmp2105;
  assign tmp2120 = s7 ? 1 : tmp2121;
  assign tmp2119 = s8 ? tmp2103 : tmp2120;
  assign tmp2118 = s9 ? 1 : tmp2119;
  assign tmp2100 = s10 ? tmp2101 : tmp2118;
  assign tmp2133 = l1 ? 1 : tmp2112;
  assign tmp2132 = s0 ? tmp2133 : 1;
  assign tmp2131 = s1 ? 1 : tmp2132;
  assign tmp2130 = s2 ? 1 : tmp2131;
  assign tmp2129 = s3 ? 1 : tmp2130;
  assign tmp2134 = s3 ? 1 : tmp2131;
  assign tmp2128 = s4 ? tmp2129 : tmp2134;
  assign tmp2127 = s5 ? 1 : tmp2128;
  assign tmp2126 = s6 ? tmp2127 : 1;
  assign tmp2125 = s7 ? 1 : tmp2126;
  assign tmp2138 = s4 ? tmp2129 : 1;
  assign tmp2137 = s5 ? 1 : tmp2138;
  assign tmp2136 = s6 ? 1 : tmp2137;
  assign tmp2135 = s7 ? 1 : tmp2136;
  assign tmp2124 = s8 ? tmp2125 : tmp2135;
  assign tmp2123 = s9 ? 1 : tmp2124;
  assign tmp2142 = s6 ? 1 : tmp2127;
  assign tmp2141 = s7 ? 1 : tmp2142;
  assign tmp2140 = s8 ? tmp2125 : tmp2141;
  assign tmp2139 = s9 ? 1 : tmp2140;
  assign tmp2122 = s10 ? tmp2123 : tmp2139;
  assign tmp2099 = s11 ? tmp2100 : tmp2122;
  assign tmp2049 = s12 ? tmp2050 : tmp2099;
  assign tmp2156 = l1 ? 1 : tmp2063;
  assign tmp2155 = ~(s0 ? tmp2156 : 0);
  assign tmp2154 = s1 ? 1 : tmp2155;
  assign tmp2153 = s2 ? tmp2154 : 1;
  assign tmp2157 = s2 ? 1 : tmp2087;
  assign tmp2152 = s3 ? tmp2153 : tmp2157;
  assign tmp2151 = s4 ? 1 : tmp2152;
  assign tmp2150 = s5 ? 1 : tmp2151;
  assign tmp2149 = s6 ? tmp2150 : 1;
  assign tmp2148 = s7 ? 1 : tmp2149;
  assign tmp2162 = s3 ? tmp2153 : 1;
  assign tmp2161 = s4 ? 1 : tmp2162;
  assign tmp2160 = s5 ? 1 : tmp2161;
  assign tmp2159 = s6 ? 1 : tmp2160;
  assign tmp2158 = s7 ? 1 : tmp2159;
  assign tmp2147 = s8 ? tmp2148 : tmp2158;
  assign tmp2146 = s9 ? 1 : tmp2147;
  assign tmp2166 = s6 ? 1 : tmp2150;
  assign tmp2165 = s7 ? 1 : tmp2166;
  assign tmp2164 = s8 ? tmp2148 : tmp2165;
  assign tmp2163 = s9 ? 1 : tmp2164;
  assign tmp2145 = s10 ? tmp2146 : tmp2163;
  assign tmp2175 = s2 ? tmp2066 : 1;
  assign tmp2174 = s3 ? 1 : tmp2175;
  assign tmp2177 = ~(s1 ? tmp2061 : 0);
  assign tmp2176 = s3 ? 1 : tmp2177;
  assign tmp2173 = s4 ? tmp2174 : tmp2176;
  assign tmp2172 = s5 ? 1 : tmp2173;
  assign tmp2171 = s6 ? tmp2172 : 1;
  assign tmp2170 = s7 ? 1 : tmp2171;
  assign tmp2181 = s4 ? tmp2174 : 1;
  assign tmp2180 = s5 ? 1 : tmp2181;
  assign tmp2179 = s6 ? 1 : tmp2180;
  assign tmp2178 = s7 ? 1 : tmp2179;
  assign tmp2169 = s8 ? tmp2170 : tmp2178;
  assign tmp2168 = s9 ? 1 : tmp2169;
  assign tmp2185 = s6 ? 1 : tmp2172;
  assign tmp2184 = s7 ? 1 : tmp2185;
  assign tmp2183 = s8 ? tmp2170 : tmp2184;
  assign tmp2182 = s9 ? 1 : tmp2183;
  assign tmp2167 = s10 ? tmp2168 : tmp2182;
  assign tmp2144 = s11 ? tmp2145 : tmp2167;
  assign tmp2198 = l1 ? tmp2063 : 0;
  assign tmp2197 = s0 ? tmp2198 : 0;
  assign tmp2196 = ~(s1 ? tmp2197 : 0);
  assign tmp2195 = s2 ? 1 : tmp2196;
  assign tmp2200 = ~(l1 ? tmp2063 : 0);
  assign tmp2199 = s2 ? 1 : tmp2200;
  assign tmp2194 = s3 ? tmp2195 : tmp2199;
  assign tmp2193 = s4 ? 1 : tmp2194;
  assign tmp2192 = s5 ? 1 : tmp2193;
  assign tmp2191 = s6 ? tmp2192 : 1;
  assign tmp2190 = s7 ? 1 : tmp2191;
  assign tmp2205 = s3 ? tmp2195 : 1;
  assign tmp2204 = s4 ? 1 : tmp2205;
  assign tmp2203 = s5 ? 1 : tmp2204;
  assign tmp2202 = s6 ? 1 : tmp2203;
  assign tmp2201 = s7 ? 1 : tmp2202;
  assign tmp2189 = s8 ? tmp2190 : tmp2201;
  assign tmp2188 = s9 ? 1 : tmp2189;
  assign tmp2209 = s6 ? 1 : tmp2192;
  assign tmp2208 = s7 ? 1 : tmp2209;
  assign tmp2207 = s8 ? tmp2190 : tmp2208;
  assign tmp2206 = s9 ? 1 : tmp2207;
  assign tmp2187 = s10 ? tmp2188 : tmp2206;
  assign tmp2186 = s11 ? 1 : tmp2187;
  assign tmp2143 = s12 ? tmp2144 : tmp2186;
  assign tmp2048 = s13 ? tmp2049 : tmp2143;
  assign tmp2047 = s15 ? 1 : tmp2048;
  assign tmp2046 = ~(s16 ? 1 : tmp2047);
  assign s15n = tmp2046;

  assign s14n = 0;

  assign tmp2218 = l3 ? 1 : 0;
  assign tmp2217 = l1 ? 1 : tmp2218;
  assign tmp2222 = s1 ? tmp2217 : 1;
  assign tmp2223 = s0 ? tmp2217 : 1;
  assign tmp2221 = s2 ? tmp2222 : tmp2223;
  assign tmp2226 = s0 ? 1 : tmp2218;
  assign tmp2225 = s1 ? 1 : tmp2226;
  assign tmp2224 = s2 ? tmp2225 : tmp2217;
  assign tmp2220 = s3 ? tmp2221 : tmp2224;
  assign tmp2230 = s0 ? tmp2217 : 0;
  assign tmp2232 = ~(l1 ? 1 : 0);
  assign tmp2231 = ~(s0 ? 1 : tmp2232);
  assign tmp2229 = s1 ? tmp2230 : tmp2231;
  assign tmp2234 = l1 ? 1 : 0;
  assign tmp2233 = s1 ? tmp2217 : tmp2234;
  assign tmp2228 = s2 ? tmp2229 : tmp2233;
  assign tmp2237 = s0 ? 1 : tmp2217;
  assign tmp2236 = s1 ? tmp2237 : tmp2217;
  assign tmp2235 = s2 ? tmp2236 : tmp2230;
  assign tmp2227 = s3 ? tmp2228 : tmp2235;
  assign tmp2219 = s4 ? tmp2220 : tmp2227;
  assign tmp2216 = s5 ? tmp2217 : tmp2219;
  assign tmp2246 = s0 ? tmp2218 : 1;
  assign tmp2245 = s1 ? tmp2246 : tmp2217;
  assign tmp2244 = s2 ? tmp2225 : tmp2245;
  assign tmp2243 = s3 ? tmp2221 : tmp2244;
  assign tmp2250 = s0 ? tmp2234 : tmp2217;
  assign tmp2249 = s1 ? tmp2250 : tmp2234;
  assign tmp2248 = s2 ? tmp2229 : tmp2249;
  assign tmp2253 = s0 ? tmp2218 : tmp2234;
  assign tmp2252 = s1 ? tmp2230 : tmp2253;
  assign tmp2251 = s2 ? tmp2236 : tmp2252;
  assign tmp2247 = s3 ? tmp2248 : tmp2251;
  assign tmp2242 = s4 ? tmp2243 : tmp2247;
  assign tmp2241 = s5 ? tmp2217 : tmp2242;
  assign tmp2240 = s6 ? tmp2241 : tmp2216;
  assign tmp2259 = s1 ? tmp2217 : tmp2223;
  assign tmp2258 = s2 ? tmp2222 : tmp2259;
  assign tmp2261 = s1 ? 1 : tmp2218;
  assign tmp2262 = s1 ? 1 : tmp2217;
  assign tmp2260 = s2 ? tmp2261 : tmp2262;
  assign tmp2257 = s3 ? tmp2258 : tmp2260;
  assign tmp2265 = s1 ? 1 : tmp2232;
  assign tmp2266 = ~(s1 ? tmp2217 : tmp2234);
  assign tmp2264 = s2 ? tmp2265 : tmp2266;
  assign tmp2267 = ~(l1 ? 1 : tmp2218);
  assign tmp2263 = ~(s3 ? tmp2264 : tmp2267);
  assign tmp2256 = s4 ? tmp2257 : tmp2263;
  assign tmp2255 = s5 ? tmp2217 : tmp2256;
  assign tmp2272 = s1 ? tmp2246 : tmp2237;
  assign tmp2271 = s2 ? tmp2225 : tmp2272;
  assign tmp2270 = s3 ? tmp2221 : tmp2271;
  assign tmp2276 = s0 ? 1 : tmp2234;
  assign tmp2275 = s1 ? tmp2250 : tmp2276;
  assign tmp2274 = s2 ? tmp2229 : tmp2275;
  assign tmp2277 = s2 ? tmp2237 : tmp2252;
  assign tmp2273 = s3 ? tmp2274 : tmp2277;
  assign tmp2269 = s4 ? tmp2270 : tmp2273;
  assign tmp2268 = s5 ? tmp2217 : tmp2269;
  assign tmp2254 = s6 ? tmp2255 : tmp2268;
  assign tmp2239 = s7 ? tmp2240 : tmp2254;
  assign tmp2282 = s3 ? tmp2258 : tmp2224;
  assign tmp2283 = s3 ? tmp2228 : tmp2217;
  assign tmp2281 = s4 ? tmp2282 : tmp2283;
  assign tmp2280 = s5 ? tmp2217 : tmp2281;
  assign tmp2279 = s6 ? tmp2241 : tmp2280;
  assign tmp2284 = s6 ? tmp2280 : tmp2255;
  assign tmp2278 = s7 ? tmp2279 : tmp2284;
  assign tmp2238 = s8 ? tmp2239 : tmp2278;
  assign tmp2215 = s9 ? tmp2216 : tmp2238;
  assign tmp2288 = s6 ? tmp2216 : tmp2255;
  assign tmp2287 = s7 ? tmp2240 : tmp2288;
  assign tmp2286 = s8 ? tmp2239 : tmp2287;
  assign tmp2285 = s9 ? tmp2216 : tmp2286;
  assign tmp2214 = s10 ? tmp2215 : tmp2285;
  assign tmp2292 = l1 ? tmp2218 : 1;
  assign tmp2296 = s1 ? tmp2292 : 1;
  assign tmp2297 = s0 ? tmp2292 : 1;
  assign tmp2295 = s2 ? tmp2296 : tmp2297;
  assign tmp2300 = s0 ? 1 : tmp2232;
  assign tmp2299 = s1 ? 1 : tmp2300;
  assign tmp2298 = s2 ? tmp2299 : tmp2292;
  assign tmp2294 = s3 ? tmp2295 : tmp2298;
  assign tmp2303 = s1 ? tmp2292 : tmp2218;
  assign tmp2302 = s2 ? tmp2218 : tmp2303;
  assign tmp2305 = s0 ? 1 : tmp2292;
  assign tmp2304 = s1 ? tmp2305 : tmp2292;
  assign tmp2301 = s3 ? tmp2302 : tmp2304;
  assign tmp2293 = s4 ? tmp2294 : tmp2301;
  assign tmp2291 = s5 ? tmp2292 : tmp2293;
  assign tmp2315 = ~(l1 ? tmp2218 : 1);
  assign tmp2314 = s0 ? tmp2234 : tmp2315;
  assign tmp2313 = ~(s1 ? tmp2314 : tmp2315);
  assign tmp2312 = s2 ? tmp2299 : tmp2313;
  assign tmp2311 = s3 ? tmp2295 : tmp2312;
  assign tmp2317 = s2 ? tmp2225 : tmp2303;
  assign tmp2321 = ~(l3 ? 1 : 0);
  assign tmp2320 = ~(s0 ? tmp2234 : tmp2321);
  assign tmp2319 = s1 ? 1 : tmp2320;
  assign tmp2318 = s2 ? tmp2304 : tmp2319;
  assign tmp2316 = s3 ? tmp2317 : tmp2318;
  assign tmp2310 = s4 ? tmp2311 : tmp2316;
  assign tmp2309 = s5 ? tmp2292 : tmp2310;
  assign tmp2325 = s2 ? tmp2261 : tmp2303;
  assign tmp2324 = s3 ? tmp2325 : tmp2304;
  assign tmp2323 = s4 ? tmp2294 : tmp2324;
  assign tmp2322 = s5 ? tmp2292 : tmp2323;
  assign tmp2308 = s6 ? tmp2309 : tmp2322;
  assign tmp2331 = s1 ? tmp2292 : tmp2297;
  assign tmp2330 = s2 ? tmp2296 : tmp2331;
  assign tmp2332 = s2 ? tmp2265 : tmp2296;
  assign tmp2329 = s3 ? tmp2330 : tmp2332;
  assign tmp2334 = s2 ? tmp2261 : tmp2292;
  assign tmp2333 = s3 ? tmp2334 : tmp2292;
  assign tmp2328 = s4 ? tmp2329 : tmp2333;
  assign tmp2327 = s5 ? tmp2292 : tmp2328;
  assign tmp2340 = ~(s0 ? tmp2292 : 1);
  assign tmp2339 = ~(s1 ? tmp2314 : tmp2340);
  assign tmp2338 = s2 ? tmp2299 : tmp2339;
  assign tmp2337 = s3 ? tmp2295 : tmp2338;
  assign tmp2343 = s1 ? tmp2292 : tmp2305;
  assign tmp2342 = s2 ? tmp2225 : tmp2343;
  assign tmp2341 = s3 ? tmp2342 : tmp2318;
  assign tmp2336 = s4 ? tmp2337 : tmp2341;
  assign tmp2335 = s5 ? tmp2292 : tmp2336;
  assign tmp2326 = s6 ? tmp2327 : tmp2335;
  assign tmp2307 = s7 ? tmp2308 : tmp2326;
  assign tmp2348 = s3 ? tmp2325 : tmp2318;
  assign tmp2347 = s4 ? tmp2311 : tmp2348;
  assign tmp2346 = s5 ? tmp2292 : tmp2347;
  assign tmp2351 = s3 ? tmp2330 : tmp2298;
  assign tmp2353 = s2 ? tmp2218 : tmp2292;
  assign tmp2352 = s3 ? tmp2353 : tmp2292;
  assign tmp2350 = s4 ? tmp2351 : tmp2352;
  assign tmp2349 = s5 ? tmp2292 : tmp2350;
  assign tmp2345 = s6 ? tmp2346 : tmp2349;
  assign tmp2356 = s4 ? tmp2351 : tmp2333;
  assign tmp2355 = s5 ? tmp2292 : tmp2356;
  assign tmp2354 = s6 ? tmp2355 : tmp2327;
  assign tmp2344 = s7 ? tmp2345 : tmp2354;
  assign tmp2306 = s8 ? tmp2307 : tmp2344;
  assign tmp2290 = s9 ? tmp2291 : tmp2306;
  assign tmp2360 = s6 ? tmp2346 : tmp2291;
  assign tmp2361 = s6 ? tmp2322 : tmp2327;
  assign tmp2359 = s7 ? tmp2360 : tmp2361;
  assign tmp2358 = s8 ? tmp2307 : tmp2359;
  assign tmp2357 = s9 ? tmp2291 : tmp2358;
  assign tmp2289 = s10 ? tmp2290 : tmp2357;
  assign tmp2213 = s11 ? tmp2214 : tmp2289;
  assign tmp2212 = s12 ? 1 : tmp2213;
  assign tmp2363 = s11 ? 1 : 0;
  assign tmp2368 = l1 ? 1 : tmp2321;
  assign tmp2372 = s1 ? 1 : tmp2368;
  assign tmp2373 = s1 ? tmp2368 : tmp2321;
  assign tmp2371 = s2 ? tmp2372 : tmp2373;
  assign tmp2370 = s3 ? tmp2368 : tmp2371;
  assign tmp2376 = s1 ? tmp2368 : 1;
  assign tmp2375 = s2 ? 1 : tmp2376;
  assign tmp2377 = s2 ? tmp2368 : tmp2372;
  assign tmp2374 = s3 ? tmp2375 : tmp2377;
  assign tmp2369 = s4 ? tmp2370 : tmp2374;
  assign tmp2367 = s5 ? tmp2368 : tmp2369;
  assign tmp2386 = s0 ? tmp2368 : 0;
  assign tmp2385 = s1 ? tmp2368 : tmp2386;
  assign tmp2384 = s2 ? tmp2368 : tmp2385;
  assign tmp2389 = s0 ? 1 : 0;
  assign tmp2390 = ~(s0 ? 1 : tmp2368);
  assign tmp2388 = s1 ? tmp2389 : tmp2390;
  assign tmp2391 = ~(l1 ? 1 : tmp2321);
  assign tmp2387 = ~(s2 ? tmp2388 : tmp2391);
  assign tmp2383 = s3 ? tmp2384 : tmp2387;
  assign tmp2395 = s0 ? tmp2218 : 0;
  assign tmp2394 = s1 ? tmp2395 : 0;
  assign tmp2397 = s0 ? 1 : tmp2368;
  assign tmp2398 = ~(s0 ? 1 : 0);
  assign tmp2396 = ~(s1 ? tmp2397 : tmp2398);
  assign tmp2393 = s2 ? tmp2394 : tmp2396;
  assign tmp2400 = s1 ? tmp2397 : tmp2368;
  assign tmp2401 = s0 ? tmp2368 : 1;
  assign tmp2399 = ~(s2 ? tmp2400 : tmp2401);
  assign tmp2392 = ~(s3 ? tmp2393 : tmp2399);
  assign tmp2382 = s4 ? tmp2383 : tmp2392;
  assign tmp2381 = s5 ? tmp2368 : tmp2382;
  assign tmp2404 = s3 ? tmp2384 : tmp2371;
  assign tmp2403 = s4 ? tmp2404 : tmp2374;
  assign tmp2402 = s5 ? tmp2368 : tmp2403;
  assign tmp2380 = s6 ? tmp2381 : tmp2402;
  assign tmp2409 = ~(s0 ? tmp2218 : tmp2391);
  assign tmp2408 = s1 ? tmp2368 : tmp2409;
  assign tmp2407 = s2 ? tmp2368 : tmp2408;
  assign tmp2413 = s1 ? tmp2368 : 0;
  assign tmp2412 = s2 ? tmp2413 : tmp2385;
  assign tmp2416 = s0 ? tmp2368 : tmp2234;
  assign tmp2415 = s1 ? tmp2416 : tmp2321;
  assign tmp2414 = s2 ? tmp2372 : tmp2415;
  assign tmp2411 = s3 ? tmp2412 : tmp2414;
  assign tmp2417 = s3 ? tmp2375 : tmp2368;
  assign tmp2410 = s4 ? tmp2411 : tmp2417;
  assign tmp2406 = s5 ? tmp2407 : tmp2410;
  assign tmp2423 = s0 ? tmp2234 : tmp2321;
  assign tmp2422 = ~(s1 ? tmp2416 : tmp2423);
  assign tmp2421 = ~(s2 ? tmp2388 : tmp2422);
  assign tmp2420 = s3 ? tmp2412 : tmp2421;
  assign tmp2427 = s0 ? tmp2234 : tmp2368;
  assign tmp2426 = s1 ? tmp2397 : tmp2427;
  assign tmp2425 = ~(s2 ? tmp2426 : tmp2401);
  assign tmp2424 = ~(s3 ? tmp2393 : tmp2425);
  assign tmp2419 = s4 ? tmp2420 : tmp2424;
  assign tmp2418 = s5 ? tmp2407 : tmp2419;
  assign tmp2405 = s6 ? tmp2406 : tmp2418;
  assign tmp2379 = s7 ? tmp2380 : tmp2405;
  assign tmp2434 = s1 ? 1 : tmp2397;
  assign tmp2433 = s2 ? tmp2434 : tmp2368;
  assign tmp2432 = s3 ? tmp2368 : tmp2433;
  assign tmp2437 = ~(s1 ? tmp2397 : 1);
  assign tmp2436 = s2 ? tmp2394 : tmp2437;
  assign tmp2435 = ~(s3 ? tmp2436 : tmp2399);
  assign tmp2431 = s4 ? tmp2432 : tmp2435;
  assign tmp2430 = s5 ? tmp2368 : tmp2431;
  assign tmp2441 = s2 ? tmp2368 : tmp2401;
  assign tmp2440 = s3 ? tmp2441 : tmp2371;
  assign tmp2439 = s4 ? tmp2440 : tmp2417;
  assign tmp2438 = s5 ? tmp2368 : tmp2439;
  assign tmp2429 = s6 ? tmp2430 : tmp2438;
  assign tmp2444 = s4 ? tmp2404 : tmp2417;
  assign tmp2443 = s5 ? tmp2368 : tmp2444;
  assign tmp2442 = s6 ? tmp2443 : tmp2406;
  assign tmp2428 = s7 ? tmp2429 : tmp2442;
  assign tmp2378 = s8 ? tmp2379 : tmp2428;
  assign tmp2366 = s9 ? tmp2367 : tmp2378;
  assign tmp2448 = s6 ? tmp2430 : tmp2367;
  assign tmp2449 = s6 ? tmp2402 : tmp2406;
  assign tmp2447 = s7 ? tmp2448 : tmp2449;
  assign tmp2446 = s8 ? tmp2379 : tmp2447;
  assign tmp2445 = s9 ? tmp2367 : tmp2446;
  assign tmp2365 = s10 ? tmp2366 : tmp2445;
  assign tmp2453 = l1 ? tmp2218 : 0;
  assign tmp2457 = s1 ? tmp2453 : 0;
  assign tmp2456 = s2 ? tmp2457 : tmp2453;
  assign tmp2459 = s1 ? 1 : tmp2389;
  assign tmp2458 = s2 ? tmp2459 : tmp2453;
  assign tmp2455 = s3 ? tmp2456 : tmp2458;
  assign tmp2464 = ~(l1 ? tmp2218 : 0);
  assign tmp2463 = s0 ? 1 : tmp2464;
  assign tmp2462 = s1 ? 1 : tmp2463;
  assign tmp2461 = s2 ? tmp2462 : tmp2464;
  assign tmp2466 = ~(s1 ? 1 : tmp2464);
  assign tmp2465 = ~(s2 ? tmp2453 : tmp2466);
  assign tmp2460 = ~(s3 ? tmp2461 : tmp2465);
  assign tmp2454 = s4 ? tmp2455 : tmp2460;
  assign tmp2452 = s5 ? tmp2453 : tmp2454;
  assign tmp2474 = s1 ? tmp2453 : 1;
  assign tmp2476 = s0 ? tmp2453 : 1;
  assign tmp2475 = s1 ? tmp2476 : tmp2453;
  assign tmp2473 = s2 ? tmp2474 : tmp2475;
  assign tmp2479 = s0 ? 1 : tmp2321;
  assign tmp2478 = ~(s1 ? tmp2479 : tmp2464);
  assign tmp2477 = s2 ? tmp2459 : tmp2478;
  assign tmp2472 = s3 ? tmp2473 : tmp2477;
  assign tmp2483 = s0 ? tmp2234 : 0;
  assign tmp2484 = ~(s0 ? 1 : tmp2464);
  assign tmp2482 = s1 ? tmp2483 : tmp2484;
  assign tmp2481 = s2 ? tmp2482 : tmp2453;
  assign tmp2485 = s2 ? tmp2453 : tmp2482;
  assign tmp2480 = s3 ? tmp2481 : tmp2485;
  assign tmp2471 = s4 ? tmp2472 : tmp2480;
  assign tmp2470 = s5 ? tmp2453 : tmp2471;
  assign tmp2489 = s2 ? tmp2474 : tmp2453;
  assign tmp2488 = s3 ? tmp2489 : tmp2458;
  assign tmp2487 = s4 ? tmp2488 : tmp2460;
  assign tmp2486 = s5 ? tmp2453 : tmp2487;
  assign tmp2469 = s6 ? tmp2470 : tmp2486;
  assign tmp2494 = l2 ? 1 : 0;
  assign tmp2493 = l1 ? tmp2218 : tmp2494;
  assign tmp2495 = s0 ? tmp2493 : tmp2453;
  assign tmp2492 = s2 ? tmp2493 : tmp2495;
  assign tmp2500 = s0 ? tmp2234 : tmp2493;
  assign tmp2499 = s1 ? tmp2500 : 1;
  assign tmp2502 = s0 ? tmp2493 : 1;
  assign tmp2501 = s1 ? tmp2493 : tmp2502;
  assign tmp2498 = s2 ? tmp2499 : tmp2501;
  assign tmp2504 = s1 ? 1 : 0;
  assign tmp2505 = s1 ? tmp2218 : tmp2234;
  assign tmp2503 = s2 ? tmp2504 : tmp2505;
  assign tmp2497 = s3 ? tmp2498 : tmp2503;
  assign tmp2508 = s1 ? 1 : tmp2464;
  assign tmp2509 = ~(s1 ? tmp2493 : tmp2453);
  assign tmp2507 = s2 ? tmp2508 : tmp2509;
  assign tmp2506 = ~(s3 ? tmp2507 : tmp2464);
  assign tmp2496 = s4 ? tmp2497 : tmp2506;
  assign tmp2491 = s5 ? tmp2492 : tmp2496;
  assign tmp2513 = s2 ? tmp2499 : tmp2502;
  assign tmp2516 = ~(s0 ? tmp2218 : tmp2234);
  assign tmp2515 = ~(s1 ? tmp2479 : tmp2516);
  assign tmp2514 = s2 ? tmp2459 : tmp2515;
  assign tmp2512 = s3 ? tmp2513 : tmp2514;
  assign tmp2520 = s0 ? tmp2453 : tmp2493;
  assign tmp2521 = s0 ? 1 : tmp2453;
  assign tmp2519 = s1 ? tmp2520 : tmp2521;
  assign tmp2518 = s2 ? tmp2482 : tmp2519;
  assign tmp2524 = s0 ? tmp2218 : tmp2453;
  assign tmp2523 = s1 ? tmp2521 : tmp2524;
  assign tmp2522 = s2 ? tmp2523 : tmp2482;
  assign tmp2517 = s3 ? tmp2518 : tmp2522;
  assign tmp2511 = s4 ? tmp2512 : tmp2517;
  assign tmp2510 = s5 ? tmp2492 : tmp2511;
  assign tmp2490 = s6 ? tmp2491 : tmp2510;
  assign tmp2468 = s7 ? tmp2469 : tmp2490;
  assign tmp2532 = s0 ? tmp2453 : 0;
  assign tmp2531 = s1 ? tmp2532 : tmp2453;
  assign tmp2530 = s2 ? tmp2457 : tmp2531;
  assign tmp2529 = s3 ? tmp2530 : tmp2477;
  assign tmp2528 = s4 ? tmp2529 : tmp2480;
  assign tmp2527 = s5 ? tmp2453 : tmp2528;
  assign tmp2535 = ~(s3 ? tmp2461 : tmp2464);
  assign tmp2534 = s4 ? tmp2455 : tmp2535;
  assign tmp2533 = s5 ? tmp2453 : tmp2534;
  assign tmp2526 = s6 ? tmp2527 : tmp2533;
  assign tmp2538 = s4 ? tmp2488 : tmp2535;
  assign tmp2537 = s5 ? tmp2453 : tmp2538;
  assign tmp2536 = s6 ? tmp2537 : tmp2491;
  assign tmp2525 = s7 ? tmp2526 : tmp2536;
  assign tmp2467 = s8 ? tmp2468 : tmp2525;
  assign tmp2451 = s9 ? tmp2452 : tmp2467;
  assign tmp2542 = s6 ? tmp2527 : tmp2452;
  assign tmp2543 = s6 ? tmp2486 : tmp2491;
  assign tmp2541 = s7 ? tmp2542 : tmp2543;
  assign tmp2540 = s8 ? tmp2468 : tmp2541;
  assign tmp2539 = s9 ? tmp2452 : tmp2540;
  assign tmp2450 = ~(s10 ? tmp2451 : tmp2539);
  assign tmp2364 = s11 ? tmp2365 : tmp2450;
  assign tmp2362 = ~(s12 ? tmp2363 : tmp2364);
  assign tmp2211 = s13 ? tmp2212 : tmp2362;
  assign tmp2556 = s2 ? tmp2504 : 0;
  assign tmp2555 = ~(s3 ? tmp2556 : 0);
  assign tmp2554 = s4 ? 1 : tmp2555;
  assign tmp2553 = s5 ? 1 : tmp2554;
  assign tmp2561 = s1 ? tmp2389 : tmp2398;
  assign tmp2560 = s2 ? tmp2561 : 1;
  assign tmp2562 = s2 ? 1 : tmp2389;
  assign tmp2559 = s3 ? tmp2560 : tmp2562;
  assign tmp2558 = s4 ? 1 : tmp2559;
  assign tmp2557 = s5 ? 1 : tmp2558;
  assign tmp2552 = s6 ? tmp2553 : tmp2557;
  assign tmp2551 = s7 ? tmp2240 : tmp2552;
  assign tmp2564 = s6 ? tmp2280 : tmp2553;
  assign tmp2563 = s7 ? 1 : tmp2564;
  assign tmp2550 = s8 ? tmp2551 : tmp2563;
  assign tmp2549 = s9 ? 1 : tmp2550;
  assign tmp2568 = s6 ? tmp2216 : tmp2553;
  assign tmp2567 = s7 ? 1 : tmp2568;
  assign tmp2566 = s8 ? tmp2551 : tmp2567;
  assign tmp2565 = s9 ? 1 : tmp2566;
  assign tmp2548 = s10 ? tmp2549 : tmp2565;
  assign tmp2576 = l1 ? tmp2494 : 1;
  assign tmp2578 = s0 ? tmp2576 : tmp2494;
  assign tmp2577 = s1 ? tmp2578 : tmp2576;
  assign tmp2575 = s2 ? tmp2576 : tmp2577;
  assign tmp2582 = s1 ? tmp2576 : 1;
  assign tmp2584 = s0 ? tmp2576 : 1;
  assign tmp2583 = s1 ? tmp2576 : tmp2584;
  assign tmp2581 = s2 ? tmp2582 : tmp2583;
  assign tmp2586 = ~(s1 ? 1 : 0);
  assign tmp2585 = s2 ? tmp2504 : tmp2586;
  assign tmp2580 = s3 ? tmp2581 : tmp2585;
  assign tmp2589 = s1 ? tmp2576 : tmp2232;
  assign tmp2588 = s2 ? tmp2504 : tmp2589;
  assign tmp2591 = ~(l1 ? tmp2494 : 1);
  assign tmp2590 = ~(s1 ? 1 : tmp2591);
  assign tmp2587 = s3 ? tmp2588 : tmp2590;
  assign tmp2579 = s4 ? tmp2580 : tmp2587;
  assign tmp2574 = s5 ? tmp2575 : tmp2579;
  assign tmp2595 = s2 ? tmp2582 : tmp2584;
  assign tmp2597 = ~(s1 ? 1 : tmp2389);
  assign tmp2596 = s2 ? tmp2459 : tmp2597;
  assign tmp2594 = s3 ? tmp2595 : tmp2596;
  assign tmp2601 = s0 ? 1 : tmp2591;
  assign tmp2600 = ~(s1 ? tmp2601 : tmp2231);
  assign tmp2599 = s2 ? tmp2459 : tmp2600;
  assign tmp2604 = ~(s0 ? 1 : tmp2591);
  assign tmp2603 = s1 ? tmp2389 : tmp2604;
  assign tmp2602 = s2 ? tmp2603 : tmp2504;
  assign tmp2598 = s3 ? tmp2599 : tmp2602;
  assign tmp2593 = s4 ? tmp2594 : tmp2598;
  assign tmp2592 = s5 ? tmp2575 : tmp2593;
  assign tmp2573 = s6 ? tmp2574 : tmp2592;
  assign tmp2572 = s7 ? tmp2308 : tmp2573;
  assign tmp2606 = ~(s6 ? tmp2355 : tmp2574);
  assign tmp2605 = ~(s7 ? 1 : tmp2606);
  assign tmp2571 = ~(s8 ? tmp2572 : tmp2605);
  assign tmp2570 = s9 ? 1 : tmp2571;
  assign tmp2610 = ~(s6 ? tmp2322 : tmp2574);
  assign tmp2609 = ~(s7 ? 1 : tmp2610);
  assign tmp2608 = ~(s8 ? tmp2572 : tmp2609);
  assign tmp2607 = s9 ? 1 : tmp2608;
  assign tmp2569 = ~(s10 ? tmp2570 : tmp2607);
  assign tmp2547 = s11 ? tmp2548 : tmp2569;
  assign tmp2546 = s12 ? 1 : tmp2547;
  assign tmp2620 = s1 ? tmp2234 : tmp2398;
  assign tmp2619 = s2 ? tmp2234 : tmp2620;
  assign tmp2624 = s1 ? tmp2276 : 0;
  assign tmp2623 = s2 ? tmp2624 : tmp2234;
  assign tmp2622 = s3 ? tmp2623 : 1;
  assign tmp2627 = s1 ? tmp2234 : 1;
  assign tmp2626 = s2 ? 1 : tmp2627;
  assign tmp2625 = s3 ? tmp2626 : tmp2627;
  assign tmp2621 = s4 ? tmp2622 : tmp2625;
  assign tmp2618 = s5 ? tmp2619 : tmp2621;
  assign tmp2632 = s1 ? tmp2389 : 0;
  assign tmp2631 = ~(s2 ? tmp2632 : 0);
  assign tmp2630 = s3 ? tmp2623 : tmp2631;
  assign tmp2635 = s1 ? tmp2276 : tmp2398;
  assign tmp2634 = s2 ? 1 : tmp2635;
  assign tmp2638 = s0 ? tmp2234 : 1;
  assign tmp2637 = s1 ? 1 : tmp2638;
  assign tmp2636 = s2 ? tmp2637 : 1;
  assign tmp2633 = s3 ? tmp2634 : tmp2636;
  assign tmp2629 = s4 ? tmp2630 : tmp2633;
  assign tmp2628 = s5 ? tmp2619 : tmp2629;
  assign tmp2617 = s6 ? tmp2618 : tmp2628;
  assign tmp2616 = s7 ? tmp2380 : tmp2617;
  assign tmp2640 = s6 ? tmp2443 : tmp2618;
  assign tmp2639 = s7 ? 1 : tmp2640;
  assign tmp2615 = s8 ? tmp2616 : tmp2639;
  assign tmp2614 = s9 ? 1 : tmp2615;
  assign tmp2644 = s6 ? tmp2402 : tmp2618;
  assign tmp2643 = s7 ? 1 : tmp2644;
  assign tmp2642 = s8 ? tmp2616 : tmp2643;
  assign tmp2641 = s9 ? 1 : tmp2642;
  assign tmp2613 = s10 ? tmp2614 : tmp2641;
  assign tmp2648 = s7 ? tmp2469 : tmp2573;
  assign tmp2650 = ~(s6 ? tmp2537 : tmp2574);
  assign tmp2649 = ~(s7 ? 1 : tmp2650);
  assign tmp2647 = ~(s8 ? tmp2648 : tmp2649);
  assign tmp2646 = s9 ? 1 : tmp2647;
  assign tmp2654 = ~(s6 ? tmp2486 : tmp2574);
  assign tmp2653 = ~(s7 ? 1 : tmp2654);
  assign tmp2652 = ~(s8 ? tmp2648 : tmp2653);
  assign tmp2651 = s9 ? 1 : tmp2652;
  assign tmp2645 = s10 ? tmp2646 : tmp2651;
  assign tmp2612 = s11 ? tmp2613 : tmp2645;
  assign tmp2611 = ~(s12 ? tmp2363 : tmp2612);
  assign tmp2545 = s13 ? tmp2546 : tmp2611;
  assign tmp2670 = ~(l2 ? 1 : tmp2321);
  assign tmp2669 = l1 ? 1 : tmp2670;
  assign tmp2668 = s0 ? tmp2669 : 0;
  assign tmp2667 = s1 ? tmp2668 : tmp2234;
  assign tmp2666 = s2 ? tmp2667 : tmp2233;
  assign tmp2671 = s2 ? tmp2217 : tmp2669;
  assign tmp2665 = s3 ? tmp2666 : tmp2671;
  assign tmp2664 = s4 ? tmp2257 : tmp2665;
  assign tmp2663 = s5 ? tmp2217 : tmp2664;
  assign tmp2662 = s6 ? tmp2663 : tmp2268;
  assign tmp2661 = s7 ? tmp2240 : tmp2662;
  assign tmp2676 = s3 ? tmp2666 : tmp2217;
  assign tmp2675 = s4 ? tmp2257 : tmp2676;
  assign tmp2674 = s5 ? tmp2217 : tmp2675;
  assign tmp2673 = s6 ? tmp2280 : tmp2674;
  assign tmp2672 = s7 ? tmp2279 : tmp2673;
  assign tmp2660 = s8 ? tmp2661 : tmp2672;
  assign tmp2659 = s9 ? tmp2216 : tmp2660;
  assign tmp2680 = s6 ? tmp2216 : tmp2663;
  assign tmp2679 = s7 ? tmp2240 : tmp2680;
  assign tmp2678 = s8 ? tmp2661 : tmp2679;
  assign tmp2677 = s9 ? tmp2216 : tmp2678;
  assign tmp2658 = s10 ? tmp2659 : tmp2677;
  assign tmp2689 = s2 ? tmp2265 : tmp2331;
  assign tmp2688 = s3 ? tmp2330 : tmp2689;
  assign tmp2687 = s4 ? tmp2688 : tmp2333;
  assign tmp2686 = s5 ? tmp2292 : tmp2687;
  assign tmp2685 = s6 ? tmp2686 : tmp2335;
  assign tmp2684 = s7 ? tmp2308 : tmp2685;
  assign tmp2691 = s6 ? tmp2355 : tmp2686;
  assign tmp2690 = s7 ? tmp2345 : tmp2691;
  assign tmp2683 = s8 ? tmp2684 : tmp2690;
  assign tmp2682 = s9 ? tmp2291 : tmp2683;
  assign tmp2695 = s6 ? tmp2322 : tmp2686;
  assign tmp2694 = s7 ? tmp2360 : tmp2695;
  assign tmp2693 = s8 ? tmp2684 : tmp2694;
  assign tmp2692 = s9 ? tmp2291 : tmp2693;
  assign tmp2681 = s10 ? tmp2682 : tmp2692;
  assign tmp2657 = s11 ? tmp2658 : tmp2681;
  assign tmp2656 = s12 ? 1 : tmp2657;
  assign tmp2708 = ~(s0 ? tmp2576 : 0);
  assign tmp2707 = s1 ? 1 : tmp2708;
  assign tmp2706 = s2 ? tmp2707 : 1;
  assign tmp2705 = s3 ? 1 : tmp2706;
  assign tmp2711 = s0 ? tmp2576 : 0;
  assign tmp2710 = ~(s1 ? tmp2711 : 0);
  assign tmp2709 = s3 ? 1 : tmp2710;
  assign tmp2704 = s4 ? tmp2705 : tmp2709;
  assign tmp2703 = s5 ? 1 : tmp2704;
  assign tmp2702 = s6 ? tmp2703 : 1;
  assign tmp2701 = s7 ? 1 : tmp2702;
  assign tmp2715 = s4 ? tmp2705 : 1;
  assign tmp2714 = s5 ? 1 : tmp2715;
  assign tmp2713 = s6 ? 1 : tmp2714;
  assign tmp2712 = s7 ? 1 : tmp2713;
  assign tmp2700 = s8 ? tmp2701 : tmp2712;
  assign tmp2699 = s9 ? 1 : tmp2700;
  assign tmp2719 = s6 ? 1 : tmp2703;
  assign tmp2718 = s7 ? 1 : tmp2719;
  assign tmp2717 = s8 ? tmp2701 : tmp2718;
  assign tmp2716 = s9 ? 1 : tmp2717;
  assign tmp2698 = ~(s10 ? tmp2699 : tmp2716);
  assign tmp2697 = s11 ? 1 : tmp2698;
  assign tmp2733 = l2 ? 1 : tmp2321;
  assign tmp2732 = l1 ? tmp2733 : 1;
  assign tmp2734 = ~(l1 ? tmp2218 : tmp2494);
  assign tmp2731 = s0 ? tmp2732 : tmp2734;
  assign tmp2730 = s1 ? tmp2731 : tmp2464;
  assign tmp2729 = s2 ? tmp2508 : tmp2730;
  assign tmp2736 = ~(l1 ? tmp2733 : 1);
  assign tmp2735 = ~(s2 ? tmp2453 : tmp2736);
  assign tmp2728 = ~(s3 ? tmp2729 : tmp2735);
  assign tmp2727 = s4 ? tmp2497 : tmp2728;
  assign tmp2726 = s5 ? tmp2492 : tmp2727;
  assign tmp2725 = s6 ? tmp2726 : tmp2510;
  assign tmp2724 = s7 ? tmp2469 : tmp2725;
  assign tmp2741 = ~(s3 ? tmp2729 : tmp2464);
  assign tmp2740 = s4 ? tmp2497 : tmp2741;
  assign tmp2739 = s5 ? tmp2492 : tmp2740;
  assign tmp2738 = s6 ? tmp2537 : tmp2739;
  assign tmp2737 = s7 ? tmp2526 : tmp2738;
  assign tmp2723 = s8 ? tmp2724 : tmp2737;
  assign tmp2722 = s9 ? tmp2452 : tmp2723;
  assign tmp2745 = s6 ? tmp2486 : tmp2726;
  assign tmp2744 = s7 ? tmp2542 : tmp2745;
  assign tmp2743 = s8 ? tmp2724 : tmp2744;
  assign tmp2742 = s9 ? tmp2452 : tmp2743;
  assign tmp2721 = ~(s10 ? tmp2722 : tmp2742);
  assign tmp2720 = s11 ? tmp2365 : tmp2721;
  assign tmp2696 = ~(s12 ? tmp2697 : tmp2720);
  assign tmp2655 = s13 ? tmp2656 : tmp2696;
  assign tmp2544 = s15 ? tmp2545 : tmp2655;
  assign tmp2210 = s16 ? tmp2211 : tmp2544;
  assign s13n = tmp2210;

  assign tmp2763 = l2 ? 1 : 0;
  assign tmp2762 = l1 ? tmp2763 : 1;
  assign tmp2761 = s0 ? tmp2762 : 0;
  assign tmp2760 = s1 ? tmp2761 : 0;
  assign tmp2759 = ~(s2 ? tmp2760 : 0);
  assign tmp2758 = s3 ? 1 : tmp2759;
  assign tmp2767 = ~(s0 ? tmp2762 : 0);
  assign tmp2766 = s1 ? 1 : tmp2767;
  assign tmp2765 = s2 ? 1 : tmp2766;
  assign tmp2764 = s3 ? tmp2765 : 1;
  assign tmp2757 = s4 ? tmp2758 : tmp2764;
  assign tmp2756 = s5 ? 1 : tmp2757;
  assign tmp2755 = s6 ? tmp2756 : 1;
  assign tmp2754 = s7 ? 1 : tmp2755;
  assign tmp2771 = s4 ? tmp2758 : 1;
  assign tmp2770 = s5 ? 1 : tmp2771;
  assign tmp2769 = s6 ? 1 : tmp2770;
  assign tmp2768 = s7 ? 1 : tmp2769;
  assign tmp2753 = s8 ? tmp2754 : tmp2768;
  assign tmp2752 = s9 ? 1 : tmp2753;
  assign tmp2775 = s6 ? 1 : tmp2756;
  assign tmp2774 = s7 ? 1 : tmp2775;
  assign tmp2773 = s8 ? tmp2754 : tmp2774;
  assign tmp2772 = s9 ? 1 : tmp2773;
  assign tmp2751 = s10 ? tmp2752 : tmp2772;
  assign tmp2787 = ~(l1 ? 1 : tmp2763);
  assign tmp2786 = s0 ? 1 : tmp2787;
  assign tmp2785 = s1 ? 1 : tmp2786;
  assign tmp2788 = s1 ? tmp2786 : 1;
  assign tmp2784 = s2 ? tmp2785 : tmp2788;
  assign tmp2783 = s3 ? tmp2784 : 1;
  assign tmp2782 = s4 ? tmp2783 : 1;
  assign tmp2781 = s5 ? 1 : tmp2782;
  assign tmp2780 = s6 ? tmp2781 : 1;
  assign tmp2779 = s7 ? 1 : tmp2780;
  assign tmp2794 = s2 ? tmp2785 : 1;
  assign tmp2793 = s3 ? tmp2794 : 1;
  assign tmp2792 = s4 ? tmp2793 : 1;
  assign tmp2791 = s5 ? 1 : tmp2792;
  assign tmp2790 = s6 ? 1 : tmp2791;
  assign tmp2789 = s7 ? 1 : tmp2790;
  assign tmp2778 = s8 ? tmp2779 : tmp2789;
  assign tmp2777 = s9 ? 1 : tmp2778;
  assign tmp2798 = s6 ? 1 : tmp2781;
  assign tmp2797 = s7 ? 1 : tmp2798;
  assign tmp2796 = s8 ? tmp2779 : tmp2797;
  assign tmp2795 = s9 ? 1 : tmp2796;
  assign tmp2776 = s10 ? tmp2777 : tmp2795;
  assign tmp2750 = s11 ? tmp2751 : tmp2776;
  assign tmp2810 = s0 ? tmp2763 : 0;
  assign tmp2809 = s1 ? tmp2810 : 0;
  assign tmp2808 = s2 ? tmp2809 : 0;
  assign tmp2812 = ~(l2 ? 1 : 0);
  assign tmp2811 = ~(s2 ? 1 : tmp2812);
  assign tmp2807 = ~(s3 ? tmp2808 : tmp2811);
  assign tmp2806 = s4 ? 1 : tmp2807;
  assign tmp2805 = s5 ? 1 : tmp2806;
  assign tmp2804 = s6 ? tmp2805 : 1;
  assign tmp2803 = s7 ? 1 : tmp2804;
  assign tmp2817 = ~(s3 ? tmp2808 : 0);
  assign tmp2816 = s4 ? 1 : tmp2817;
  assign tmp2815 = s5 ? 1 : tmp2816;
  assign tmp2814 = s6 ? 1 : tmp2815;
  assign tmp2813 = s7 ? 1 : tmp2814;
  assign tmp2802 = s8 ? tmp2803 : tmp2813;
  assign tmp2801 = s9 ? 1 : tmp2802;
  assign tmp2821 = s6 ? 1 : tmp2805;
  assign tmp2820 = s7 ? 1 : tmp2821;
  assign tmp2819 = s8 ? tmp2803 : tmp2820;
  assign tmp2818 = s9 ? 1 : tmp2819;
  assign tmp2800 = s10 ? tmp2801 : tmp2818;
  assign tmp2833 = l1 ? 1 : tmp2812;
  assign tmp2832 = s0 ? tmp2833 : 1;
  assign tmp2831 = s1 ? 1 : tmp2832;
  assign tmp2830 = s2 ? 1 : tmp2831;
  assign tmp2829 = s3 ? 1 : tmp2830;
  assign tmp2834 = s3 ? 1 : tmp2831;
  assign tmp2828 = s4 ? tmp2829 : tmp2834;
  assign tmp2827 = s5 ? 1 : tmp2828;
  assign tmp2826 = s6 ? tmp2827 : 1;
  assign tmp2825 = s7 ? 1 : tmp2826;
  assign tmp2838 = s4 ? tmp2829 : 1;
  assign tmp2837 = s5 ? 1 : tmp2838;
  assign tmp2836 = s6 ? 1 : tmp2837;
  assign tmp2835 = s7 ? 1 : tmp2836;
  assign tmp2824 = s8 ? tmp2825 : tmp2835;
  assign tmp2823 = s9 ? 1 : tmp2824;
  assign tmp2842 = s6 ? 1 : tmp2827;
  assign tmp2841 = s7 ? 1 : tmp2842;
  assign tmp2840 = s8 ? tmp2825 : tmp2841;
  assign tmp2839 = s9 ? 1 : tmp2840;
  assign tmp2822 = s10 ? tmp2823 : tmp2839;
  assign tmp2799 = s11 ? tmp2800 : tmp2822;
  assign tmp2749 = s12 ? tmp2750 : tmp2799;
  assign tmp2856 = l1 ? 1 : tmp2763;
  assign tmp2855 = ~(s0 ? tmp2856 : 0);
  assign tmp2854 = s1 ? 1 : tmp2855;
  assign tmp2853 = s2 ? tmp2854 : 1;
  assign tmp2857 = s2 ? 1 : tmp2787;
  assign tmp2852 = s3 ? tmp2853 : tmp2857;
  assign tmp2851 = s4 ? 1 : tmp2852;
  assign tmp2850 = s5 ? 1 : tmp2851;
  assign tmp2849 = s6 ? tmp2850 : 1;
  assign tmp2848 = s7 ? 1 : tmp2849;
  assign tmp2862 = s3 ? tmp2853 : 1;
  assign tmp2861 = s4 ? 1 : tmp2862;
  assign tmp2860 = s5 ? 1 : tmp2861;
  assign tmp2859 = s6 ? 1 : tmp2860;
  assign tmp2858 = s7 ? 1 : tmp2859;
  assign tmp2847 = s8 ? tmp2848 : tmp2858;
  assign tmp2846 = s9 ? 1 : tmp2847;
  assign tmp2866 = s6 ? 1 : tmp2850;
  assign tmp2865 = s7 ? 1 : tmp2866;
  assign tmp2864 = s8 ? tmp2848 : tmp2865;
  assign tmp2863 = s9 ? 1 : tmp2864;
  assign tmp2845 = s10 ? tmp2846 : tmp2863;
  assign tmp2875 = s2 ? tmp2766 : 1;
  assign tmp2874 = s3 ? 1 : tmp2875;
  assign tmp2877 = ~(s1 ? tmp2761 : 0);
  assign tmp2876 = s3 ? 1 : tmp2877;
  assign tmp2873 = s4 ? tmp2874 : tmp2876;
  assign tmp2872 = s5 ? 1 : tmp2873;
  assign tmp2871 = s6 ? tmp2872 : 1;
  assign tmp2870 = s7 ? 1 : tmp2871;
  assign tmp2881 = s4 ? tmp2874 : 1;
  assign tmp2880 = s5 ? 1 : tmp2881;
  assign tmp2879 = s6 ? 1 : tmp2880;
  assign tmp2878 = s7 ? 1 : tmp2879;
  assign tmp2869 = s8 ? tmp2870 : tmp2878;
  assign tmp2868 = s9 ? 1 : tmp2869;
  assign tmp2885 = s6 ? 1 : tmp2872;
  assign tmp2884 = s7 ? 1 : tmp2885;
  assign tmp2883 = s8 ? tmp2870 : tmp2884;
  assign tmp2882 = s9 ? 1 : tmp2883;
  assign tmp2867 = s10 ? tmp2868 : tmp2882;
  assign tmp2844 = s11 ? tmp2845 : tmp2867;
  assign tmp2898 = l1 ? tmp2763 : 0;
  assign tmp2897 = s0 ? tmp2898 : 0;
  assign tmp2896 = ~(s1 ? tmp2897 : 0);
  assign tmp2895 = s2 ? 1 : tmp2896;
  assign tmp2900 = ~(l1 ? tmp2763 : 0);
  assign tmp2899 = s2 ? 1 : tmp2900;
  assign tmp2894 = s3 ? tmp2895 : tmp2899;
  assign tmp2893 = s4 ? 1 : tmp2894;
  assign tmp2892 = s5 ? 1 : tmp2893;
  assign tmp2891 = s6 ? tmp2892 : 1;
  assign tmp2890 = s7 ? 1 : tmp2891;
  assign tmp2905 = s3 ? tmp2895 : 1;
  assign tmp2904 = s4 ? 1 : tmp2905;
  assign tmp2903 = s5 ? 1 : tmp2904;
  assign tmp2902 = s6 ? 1 : tmp2903;
  assign tmp2901 = s7 ? 1 : tmp2902;
  assign tmp2889 = s8 ? tmp2890 : tmp2901;
  assign tmp2888 = s9 ? 1 : tmp2889;
  assign tmp2909 = s6 ? 1 : tmp2892;
  assign tmp2908 = s7 ? 1 : tmp2909;
  assign tmp2907 = s8 ? tmp2890 : tmp2908;
  assign tmp2906 = s9 ? 1 : tmp2907;
  assign tmp2887 = s10 ? tmp2888 : tmp2906;
  assign tmp2886 = s11 ? 1 : tmp2887;
  assign tmp2843 = s12 ? tmp2844 : tmp2886;
  assign tmp2748 = s13 ? tmp2749 : tmp2843;
  assign tmp2747 = s15 ? 1 : tmp2748;
  assign tmp2746 = ~(s16 ? 1 : tmp2747);
  assign s12n = tmp2746;

  assign tmp2913 = s11 ? 1 : 0;
  assign tmp2918 = l1 ? 1 : 0;
  assign tmp2922 = s1 ? tmp2918 : 0;
  assign tmp2924 = s0 ? tmp2918 : 0;
  assign tmp2923 = s1 ? tmp2924 : tmp2918;
  assign tmp2921 = s2 ? tmp2922 : tmp2923;
  assign tmp2927 = s0 ? 1 : 0;
  assign tmp2926 = s1 ? 1 : tmp2927;
  assign tmp2925 = s2 ? tmp2926 : tmp2918;
  assign tmp2920 = s3 ? tmp2921 : tmp2925;
  assign tmp2932 = ~(l1 ? 1 : 0);
  assign tmp2931 = ~(s0 ? 1 : tmp2932);
  assign tmp2930 = s1 ? tmp2924 : tmp2931;
  assign tmp2929 = s2 ? tmp2930 : tmp2918;
  assign tmp2933 = s2 ? tmp2918 : tmp2924;
  assign tmp2928 = s3 ? tmp2929 : tmp2933;
  assign tmp2919 = s4 ? tmp2920 : tmp2928;
  assign tmp2917 = s5 ? tmp2918 : tmp2919;
  assign tmp2942 = s0 ? 1 : tmp2932;
  assign tmp2941 = ~(s1 ? tmp2942 : tmp2932);
  assign tmp2940 = s2 ? tmp2926 : tmp2941;
  assign tmp2939 = s3 ? tmp2921 : tmp2940;
  assign tmp2944 = s2 ? tmp2918 : tmp2930;
  assign tmp2943 = s3 ? tmp2929 : tmp2944;
  assign tmp2938 = s4 ? tmp2939 : tmp2943;
  assign tmp2937 = s5 ? tmp2918 : tmp2938;
  assign tmp2936 = s6 ? tmp2937 : tmp2917;
  assign tmp2949 = s2 ? tmp2922 : tmp2918;
  assign tmp2951 = s1 ? 1 : 0;
  assign tmp2950 = s2 ? tmp2951 : tmp2918;
  assign tmp2948 = s3 ? tmp2949 : tmp2950;
  assign tmp2954 = s1 ? 1 : tmp2932;
  assign tmp2953 = s2 ? tmp2954 : tmp2932;
  assign tmp2952 = ~(s3 ? tmp2953 : tmp2932);
  assign tmp2947 = s4 ? tmp2948 : tmp2952;
  assign tmp2946 = s5 ? tmp2918 : tmp2947;
  assign tmp2945 = s6 ? tmp2946 : tmp2937;
  assign tmp2935 = s7 ? tmp2936 : tmp2945;
  assign tmp2959 = s3 ? tmp2949 : tmp2925;
  assign tmp2960 = s3 ? tmp2929 : tmp2918;
  assign tmp2958 = s4 ? tmp2959 : tmp2960;
  assign tmp2957 = s5 ? tmp2918 : tmp2958;
  assign tmp2956 = s6 ? tmp2937 : tmp2957;
  assign tmp2961 = s6 ? tmp2957 : tmp2946;
  assign tmp2955 = s7 ? tmp2956 : tmp2961;
  assign tmp2934 = s8 ? tmp2935 : tmp2955;
  assign tmp2916 = s9 ? tmp2917 : tmp2934;
  assign tmp2965 = s6 ? tmp2917 : tmp2946;
  assign tmp2964 = s7 ? tmp2936 : tmp2965;
  assign tmp2963 = s8 ? tmp2935 : tmp2964;
  assign tmp2962 = s9 ? tmp2917 : tmp2963;
  assign tmp2915 = s10 ? tmp2916 : tmp2962;
  assign tmp2973 = s0 ? tmp2918 : 1;
  assign tmp2972 = s1 ? tmp2924 : tmp2973;
  assign tmp2971 = s2 ? tmp2922 : tmp2972;
  assign tmp2976 = s0 ? 1 : tmp2918;
  assign tmp2975 = s1 ? 1 : tmp2976;
  assign tmp2974 = s2 ? tmp2975 : tmp2918;
  assign tmp2970 = s3 ? tmp2971 : tmp2974;
  assign tmp2979 = s1 ? tmp2918 : 1;
  assign tmp2978 = s2 ? 1 : tmp2979;
  assign tmp2980 = s1 ? tmp2976 : tmp2918;
  assign tmp2977 = s3 ? tmp2978 : tmp2980;
  assign tmp2969 = s4 ? tmp2970 : tmp2977;
  assign tmp2968 = s5 ? tmp2918 : tmp2969;
  assign tmp2988 = s1 ? tmp2973 : 1;
  assign tmp2987 = s2 ? tmp2988 : tmp2979;
  assign tmp2989 = s2 ? tmp2980 : tmp2973;
  assign tmp2986 = s3 ? tmp2987 : tmp2989;
  assign tmp2985 = s4 ? tmp2970 : tmp2986;
  assign tmp2984 = s5 ? tmp2918 : tmp2985;
  assign tmp2983 = s6 ? tmp2984 : tmp2968;
  assign tmp2995 = s1 ? tmp2918 : tmp2973;
  assign tmp2994 = s2 ? tmp2922 : tmp2995;
  assign tmp2997 = s1 ? 1 : tmp2918;
  assign tmp2996 = s2 ? tmp2997 : tmp2918;
  assign tmp2993 = s3 ? tmp2994 : tmp2996;
  assign tmp2999 = s2 ? 1 : tmp2918;
  assign tmp2998 = s3 ? tmp2999 : tmp2918;
  assign tmp2992 = s4 ? tmp2993 : tmp2998;
  assign tmp2991 = s5 ? tmp2918 : tmp2992;
  assign tmp2990 = s6 ? tmp2991 : tmp2984;
  assign tmp2982 = s7 ? tmp2983 : tmp2990;
  assign tmp3005 = s2 ? tmp2980 : tmp2995;
  assign tmp3004 = s3 ? tmp2979 : tmp3005;
  assign tmp3003 = s4 ? tmp2970 : tmp3004;
  assign tmp3002 = s5 ? tmp2918 : tmp3003;
  assign tmp3008 = s3 ? tmp2994 : tmp2974;
  assign tmp3007 = s4 ? tmp3008 : tmp2998;
  assign tmp3006 = s5 ? tmp2918 : tmp3007;
  assign tmp3001 = s6 ? tmp3002 : tmp3006;
  assign tmp3009 = s6 ? tmp3006 : tmp2991;
  assign tmp3000 = s7 ? tmp3001 : tmp3009;
  assign tmp2981 = s8 ? tmp2982 : tmp3000;
  assign tmp2967 = s9 ? tmp2968 : tmp2981;
  assign tmp3013 = s6 ? tmp3002 : tmp2968;
  assign tmp3014 = s6 ? tmp2968 : tmp2991;
  assign tmp3012 = s7 ? tmp3013 : tmp3014;
  assign tmp3011 = s8 ? tmp2982 : tmp3012;
  assign tmp3010 = s9 ? tmp2968 : tmp3011;
  assign tmp2966 = s10 ? tmp2967 : tmp3010;
  assign tmp2914 = s11 ? tmp2915 : tmp2966;
  assign tmp2912 = s12 ? tmp2913 : tmp2914;
  assign tmp3021 = s1 ? tmp2918 : tmp2931;
  assign tmp3020 = s2 ? tmp2918 : tmp3021;
  assign tmp3025 = s1 ? tmp2942 : 1;
  assign tmp3026 = ~(s0 ? tmp2918 : 0);
  assign tmp3024 = s2 ? tmp3025 : tmp3026;
  assign tmp3027 = ~(s2 ? tmp2918 : tmp2922);
  assign tmp3023 = s3 ? tmp3024 : tmp3027;
  assign tmp3030 = s1 ? 1 : tmp2942;
  assign tmp3029 = s2 ? tmp3030 : tmp2932;
  assign tmp3032 = ~(s1 ? 1 : tmp2932);
  assign tmp3031 = ~(s2 ? tmp2918 : tmp3032);
  assign tmp3028 = s3 ? tmp3029 : tmp3031;
  assign tmp3022 = ~(s4 ? tmp3023 : tmp3028);
  assign tmp3019 = s5 ? tmp3020 : tmp3022;
  assign tmp3040 = ~(s1 ? tmp2918 : tmp2924);
  assign tmp3039 = s2 ? tmp3030 : tmp3040;
  assign tmp3038 = s3 ? tmp3024 : tmp3039;
  assign tmp3043 = ~(s1 ? tmp2918 : tmp2931);
  assign tmp3042 = s2 ? tmp3030 : tmp3043;
  assign tmp3045 = s1 ? tmp2942 : tmp2932;
  assign tmp3044 = s2 ? tmp3045 : tmp2954;
  assign tmp3041 = s3 ? tmp3042 : tmp3044;
  assign tmp3037 = ~(s4 ? tmp3038 : tmp3041);
  assign tmp3036 = s5 ? tmp3020 : tmp3037;
  assign tmp3050 = ~(s1 ? tmp2918 : 0);
  assign tmp3049 = s2 ? tmp2954 : tmp3050;
  assign tmp3048 = s3 ? tmp3024 : tmp3049;
  assign tmp3047 = ~(s4 ? tmp3048 : tmp3028);
  assign tmp3046 = s5 ? tmp3020 : tmp3047;
  assign tmp3035 = s6 ? tmp3036 : tmp3046;
  assign tmp3055 = l2 ? 1 : 0;
  assign tmp3054 = l1 ? tmp3055 : 1;
  assign tmp3057 = s0 ? 1 : tmp3054;
  assign tmp3056 = s1 ? tmp3054 : tmp3057;
  assign tmp3053 = s2 ? tmp3054 : tmp3056;
  assign tmp3061 = s1 ? tmp3057 : 1;
  assign tmp3062 = s0 ? tmp3054 : 1;
  assign tmp3060 = s2 ? tmp3061 : tmp3062;
  assign tmp3059 = s3 ? tmp3060 : tmp3049;
  assign tmp3064 = s2 ? tmp2954 : tmp3054;
  assign tmp3065 = s2 ? tmp3054 : tmp2932;
  assign tmp3063 = s3 ? tmp3064 : tmp3065;
  assign tmp3058 = s4 ? tmp3059 : tmp3063;
  assign tmp3052 = s5 ? tmp3053 : tmp3058;
  assign tmp3068 = s3 ? tmp3060 : tmp3039;
  assign tmp3071 = s1 ? tmp3054 : tmp2942;
  assign tmp3070 = s2 ? tmp3030 : tmp3071;
  assign tmp3073 = s1 ? tmp2942 : tmp3054;
  assign tmp3072 = s2 ? tmp3073 : tmp2954;
  assign tmp3069 = s3 ? tmp3070 : tmp3072;
  assign tmp3067 = s4 ? tmp3068 : tmp3069;
  assign tmp3066 = s5 ? tmp3053 : tmp3067;
  assign tmp3051 = ~(s6 ? tmp3052 : tmp3066);
  assign tmp3034 = s7 ? tmp3035 : tmp3051;
  assign tmp3080 = s1 ? tmp2918 : tmp2924;
  assign tmp3079 = ~(s2 ? tmp2918 : tmp3080);
  assign tmp3078 = s3 ? tmp3024 : tmp3079;
  assign tmp3077 = ~(s4 ? tmp3078 : tmp3028);
  assign tmp3076 = s5 ? tmp3020 : tmp3077;
  assign tmp3084 = s2 ? tmp3025 : tmp2932;
  assign tmp3083 = s3 ? tmp3084 : tmp3027;
  assign tmp3085 = s3 ? tmp3029 : tmp2932;
  assign tmp3082 = ~(s4 ? tmp3083 : tmp3085);
  assign tmp3081 = s5 ? tmp3020 : tmp3082;
  assign tmp3075 = s6 ? tmp3076 : tmp3081;
  assign tmp3089 = s2 ? tmp3030 : tmp3054;
  assign tmp3088 = s3 ? tmp3089 : tmp3054;
  assign tmp3087 = s4 ? tmp3059 : tmp3088;
  assign tmp3086 = ~(s5 ? tmp3053 : tmp3087);
  assign tmp3074 = s7 ? tmp3075 : tmp3086;
  assign tmp3033 = s8 ? tmp3034 : tmp3074;
  assign tmp3018 = s9 ? tmp3019 : tmp3033;
  assign tmp3093 = s6 ? tmp3076 : tmp3019;
  assign tmp3097 = s2 ? tmp3054 : tmp2954;
  assign tmp3096 = s3 ? tmp3089 : tmp3097;
  assign tmp3095 = s4 ? tmp3059 : tmp3096;
  assign tmp3094 = ~(s5 ? tmp3053 : tmp3095);
  assign tmp3092 = s7 ? tmp3093 : tmp3094;
  assign tmp3091 = s8 ? tmp3034 : tmp3092;
  assign tmp3090 = s9 ? tmp3019 : tmp3091;
  assign tmp3017 = s10 ? tmp3018 : tmp3090;
  assign tmp3103 = s2 ? tmp2918 : tmp2995;
  assign tmp3104 = s2 ? tmp2975 : tmp2997;
  assign tmp3102 = s3 ? tmp3103 : tmp3104;
  assign tmp3107 = ~(s1 ? tmp2918 : tmp2976);
  assign tmp3106 = s2 ? tmp3030 : tmp3107;
  assign tmp3108 = ~(s2 ? tmp2980 : tmp3032);
  assign tmp3105 = ~(s3 ? tmp3106 : tmp3108);
  assign tmp3101 = s4 ? tmp3102 : tmp3105;
  assign tmp3100 = s5 ? tmp2918 : tmp3101;
  assign tmp3115 = s2 ? tmp2979 : tmp2973;
  assign tmp3117 = s1 ? tmp2973 : tmp2976;
  assign tmp3116 = s2 ? tmp2975 : tmp3117;
  assign tmp3114 = s3 ? tmp3115 : tmp3116;
  assign tmp3120 = s1 ? tmp2918 : tmp2976;
  assign tmp3119 = s2 ? tmp2930 : tmp3120;
  assign tmp3121 = s2 ? tmp2980 : tmp2923;
  assign tmp3118 = s3 ? tmp3119 : tmp3121;
  assign tmp3113 = s4 ? tmp3114 : tmp3118;
  assign tmp3112 = s5 ? tmp2918 : tmp3113;
  assign tmp3125 = s2 ? tmp2979 : tmp2995;
  assign tmp3124 = s3 ? tmp3125 : tmp3104;
  assign tmp3123 = s4 ? tmp3124 : tmp3105;
  assign tmp3122 = s5 ? tmp2918 : tmp3123;
  assign tmp3111 = s6 ? tmp3112 : tmp3122;
  assign tmp3129 = l1 ? 1 : tmp3055;
  assign tmp3131 = s0 ? tmp3129 : tmp2918;
  assign tmp3130 = s1 ? tmp3129 : tmp3131;
  assign tmp3128 = s2 ? tmp3129 : tmp3130;
  assign tmp3136 = s0 ? tmp2918 : tmp3129;
  assign tmp3135 = s1 ? tmp3136 : 1;
  assign tmp3138 = s0 ? tmp3129 : 1;
  assign tmp3137 = s1 ? tmp3129 : tmp3138;
  assign tmp3134 = s2 ? tmp3135 : tmp3137;
  assign tmp3133 = s3 ? tmp3134 : tmp2997;
  assign tmp3141 = ~(s1 ? tmp3129 : tmp2918);
  assign tmp3140 = s2 ? tmp2954 : tmp3141;
  assign tmp3139 = ~(s3 ? tmp3140 : tmp3141);
  assign tmp3132 = s4 ? tmp3133 : tmp3139;
  assign tmp3127 = s5 ? tmp3128 : tmp3132;
  assign tmp3145 = s2 ? tmp3135 : tmp3138;
  assign tmp3144 = s3 ? tmp3145 : tmp3116;
  assign tmp3148 = s1 ? tmp3136 : tmp2976;
  assign tmp3147 = s2 ? tmp2930 : tmp3148;
  assign tmp3151 = s0 ? 1 : tmp3129;
  assign tmp3150 = s1 ? tmp3151 : tmp2976;
  assign tmp3149 = s2 ? tmp3150 : tmp2923;
  assign tmp3146 = s3 ? tmp3147 : tmp3149;
  assign tmp3143 = s4 ? tmp3144 : tmp3146;
  assign tmp3142 = s5 ? tmp3128 : tmp3143;
  assign tmp3126 = s6 ? tmp3127 : tmp3142;
  assign tmp3110 = s7 ? tmp3111 : tmp3126;
  assign tmp3156 = s3 ? tmp3103 : tmp3116;
  assign tmp3155 = s4 ? tmp3156 : tmp3118;
  assign tmp3154 = s5 ? tmp2918 : tmp3155;
  assign tmp3159 = ~(s3 ? tmp3029 : tmp2932);
  assign tmp3158 = s4 ? tmp3102 : tmp3159;
  assign tmp3157 = s5 ? tmp2918 : tmp3158;
  assign tmp3153 = s6 ? tmp3154 : tmp3157;
  assign tmp3162 = s4 ? tmp3124 : tmp3159;
  assign tmp3161 = s5 ? tmp2918 : tmp3162;
  assign tmp3160 = s6 ? tmp3161 : tmp3127;
  assign tmp3152 = s7 ? tmp3153 : tmp3160;
  assign tmp3109 = s8 ? tmp3110 : tmp3152;
  assign tmp3099 = s9 ? tmp3100 : tmp3109;
  assign tmp3166 = s6 ? tmp3154 : tmp3100;
  assign tmp3167 = s6 ? tmp3122 : tmp3127;
  assign tmp3165 = s7 ? tmp3166 : tmp3167;
  assign tmp3164 = s8 ? tmp3110 : tmp3165;
  assign tmp3163 = s9 ? tmp3100 : tmp3164;
  assign tmp3098 = s10 ? tmp3099 : tmp3163;
  assign tmp3016 = ~(s11 ? tmp3017 : tmp3098);
  assign tmp3015 = ~(s12 ? tmp2913 : tmp3016);
  assign tmp2911 = s13 ? tmp2912 : tmp3015;
  assign tmp3176 = s6 ? tmp2946 : tmp2917;
  assign tmp3175 = s7 ? tmp2936 : tmp3176;
  assign tmp3174 = s8 ? tmp3175 : tmp2961;
  assign tmp3173 = s9 ? tmp2946 : tmp3174;
  assign tmp3178 = s8 ? tmp3175 : tmp2965;
  assign tmp3177 = s9 ? tmp2946 : tmp3178;
  assign tmp3172 = s10 ? tmp3173 : tmp3177;
  assign tmp3182 = s7 ? tmp2983 : 1;
  assign tmp3184 = s6 ? tmp3006 : 1;
  assign tmp3183 = s7 ? 1 : tmp3184;
  assign tmp3181 = s8 ? tmp3182 : tmp3183;
  assign tmp3180 = s9 ? 1 : tmp3181;
  assign tmp3188 = s6 ? tmp2968 : 1;
  assign tmp3187 = s7 ? 1 : tmp3188;
  assign tmp3186 = s8 ? tmp3182 : tmp3187;
  assign tmp3185 = s9 ? 1 : tmp3186;
  assign tmp3179 = s10 ? tmp3180 : tmp3185;
  assign tmp3171 = s11 ? tmp3172 : tmp3179;
  assign tmp3170 = s12 ? tmp2913 : tmp3171;
  assign tmp3200 = ~(s1 ? 1 : 0);
  assign tmp3199 = s2 ? tmp2951 : tmp3200;
  assign tmp3198 = s3 ? tmp3060 : tmp3199;
  assign tmp3202 = s2 ? tmp2951 : tmp3054;
  assign tmp3201 = s3 ? tmp3202 : tmp3054;
  assign tmp3197 = s4 ? tmp3198 : tmp3201;
  assign tmp3196 = s5 ? tmp3053 : tmp3197;
  assign tmp3207 = ~(s1 ? 1 : tmp2927);
  assign tmp3206 = s2 ? tmp2926 : tmp3207;
  assign tmp3205 = s3 ? tmp3060 : tmp3206;
  assign tmp3209 = s2 ? tmp2926 : tmp3071;
  assign tmp3211 = s1 ? tmp2927 : tmp3054;
  assign tmp3210 = s2 ? tmp3211 : tmp2951;
  assign tmp3208 = s3 ? tmp3209 : tmp3210;
  assign tmp3204 = s4 ? tmp3205 : tmp3208;
  assign tmp3203 = s5 ? tmp3053 : tmp3204;
  assign tmp3195 = ~(s6 ? tmp3196 : tmp3203);
  assign tmp3194 = s7 ? tmp3035 : tmp3195;
  assign tmp3215 = ~(s4 ? tmp3048 : tmp3085);
  assign tmp3214 = s5 ? tmp3020 : tmp3215;
  assign tmp3216 = ~(s5 ? tmp3053 : tmp3197);
  assign tmp3213 = s6 ? tmp3214 : tmp3216;
  assign tmp3212 = s7 ? 1 : tmp3213;
  assign tmp3193 = s8 ? tmp3194 : tmp3212;
  assign tmp3192 = s9 ? 1 : tmp3193;
  assign tmp3220 = s6 ? tmp3046 : tmp3216;
  assign tmp3219 = s7 ? 1 : tmp3220;
  assign tmp3218 = s8 ? tmp3194 : tmp3219;
  assign tmp3217 = s9 ? 1 : tmp3218;
  assign tmp3191 = s10 ? tmp3192 : tmp3217;
  assign tmp3224 = s7 ? tmp3111 : 1;
  assign tmp3226 = s6 ? tmp3161 : 1;
  assign tmp3225 = s7 ? 1 : tmp3226;
  assign tmp3223 = s8 ? tmp3224 : tmp3225;
  assign tmp3222 = s9 ? 1 : tmp3223;
  assign tmp3230 = s6 ? tmp3122 : 1;
  assign tmp3229 = s7 ? 1 : tmp3230;
  assign tmp3228 = s8 ? tmp3224 : tmp3229;
  assign tmp3227 = s9 ? 1 : tmp3228;
  assign tmp3221 = s10 ? tmp3222 : tmp3227;
  assign tmp3190 = ~(s11 ? tmp3191 : tmp3221);
  assign tmp3189 = ~(s12 ? tmp2913 : tmp3190);
  assign tmp3169 = s13 ? tmp3170 : tmp3189;
  assign tmp3242 = s2 ? tmp2988 : 1;
  assign tmp3241 = s3 ? 1 : tmp3242;
  assign tmp3245 = s1 ? 1 : tmp2973;
  assign tmp3244 = s2 ? 1 : tmp3245;
  assign tmp3243 = s3 ? tmp3244 : 1;
  assign tmp3240 = s4 ? tmp3241 : tmp3243;
  assign tmp3239 = s5 ? 1 : tmp3240;
  assign tmp3238 = s6 ? tmp3239 : 1;
  assign tmp3237 = s7 ? 1 : tmp3238;
  assign tmp3249 = s4 ? tmp3241 : 1;
  assign tmp3248 = s5 ? 1 : tmp3249;
  assign tmp3247 = s6 ? 1 : tmp3248;
  assign tmp3246 = s7 ? 1 : tmp3247;
  assign tmp3236 = s8 ? tmp3237 : tmp3246;
  assign tmp3235 = s9 ? 1 : tmp3236;
  assign tmp3253 = s6 ? 1 : tmp3239;
  assign tmp3252 = s7 ? 1 : tmp3253;
  assign tmp3251 = s8 ? tmp3237 : tmp3252;
  assign tmp3250 = s9 ? 1 : tmp3251;
  assign tmp3234 = s10 ? tmp3235 : tmp3250;
  assign tmp3262 = s2 ? tmp3030 : tmp3025;
  assign tmp3261 = s3 ? tmp3262 : 1;
  assign tmp3260 = s4 ? tmp3261 : 1;
  assign tmp3259 = s5 ? 1 : tmp3260;
  assign tmp3258 = s6 ? tmp3259 : 1;
  assign tmp3257 = s7 ? 1 : tmp3258;
  assign tmp3268 = s2 ? tmp3030 : 1;
  assign tmp3267 = s3 ? tmp3268 : 1;
  assign tmp3266 = s4 ? tmp3267 : 1;
  assign tmp3265 = s5 ? 1 : tmp3266;
  assign tmp3264 = s6 ? 1 : tmp3265;
  assign tmp3263 = s7 ? 1 : tmp3264;
  assign tmp3256 = s8 ? tmp3257 : tmp3263;
  assign tmp3255 = s9 ? 1 : tmp3256;
  assign tmp3272 = s6 ? 1 : tmp3259;
  assign tmp3271 = s7 ? 1 : tmp3272;
  assign tmp3270 = s8 ? tmp3257 : tmp3271;
  assign tmp3269 = s9 ? 1 : tmp3270;
  assign tmp3254 = ~(s10 ? tmp3255 : tmp3269);
  assign tmp3233 = s11 ? tmp3234 : tmp3254;
  assign tmp3282 = s2 ? tmp2923 : tmp2918;
  assign tmp3281 = s3 ? tmp3282 : tmp2918;
  assign tmp3280 = s4 ? tmp2948 : tmp3281;
  assign tmp3279 = s5 ? tmp2918 : tmp3280;
  assign tmp3278 = s6 ? tmp3279 : tmp2937;
  assign tmp3277 = s7 ? tmp2936 : tmp3278;
  assign tmp3284 = s6 ? tmp2957 : tmp3279;
  assign tmp3283 = s7 ? tmp2956 : tmp3284;
  assign tmp3276 = s8 ? tmp3277 : tmp3283;
  assign tmp3275 = s9 ? tmp2917 : tmp3276;
  assign tmp3288 = s6 ? tmp2917 : tmp3279;
  assign tmp3287 = s7 ? tmp2936 : tmp3288;
  assign tmp3286 = s8 ? tmp3277 : tmp3287;
  assign tmp3285 = s9 ? tmp2917 : tmp3286;
  assign tmp3274 = s10 ? tmp3275 : tmp3285;
  assign tmp3273 = s11 ? tmp3274 : tmp2966;
  assign tmp3232 = s12 ? tmp3233 : tmp3273;
  assign tmp3300 = s1 ? 1 : tmp3026;
  assign tmp3299 = s2 ? tmp3300 : 1;
  assign tmp3301 = s2 ? 1 : tmp2932;
  assign tmp3298 = s3 ? tmp3299 : tmp3301;
  assign tmp3297 = s4 ? 1 : tmp3298;
  assign tmp3296 = s5 ? 1 : tmp3297;
  assign tmp3295 = s6 ? tmp3296 : 1;
  assign tmp3294 = s7 ? 1 : tmp3295;
  assign tmp3306 = s3 ? tmp3299 : 1;
  assign tmp3305 = s4 ? 1 : tmp3306;
  assign tmp3304 = s5 ? 1 : tmp3305;
  assign tmp3303 = s6 ? 1 : tmp3304;
  assign tmp3302 = s7 ? 1 : tmp3303;
  assign tmp3293 = s8 ? tmp3294 : tmp3302;
  assign tmp3292 = s9 ? 1 : tmp3293;
  assign tmp3310 = s6 ? 1 : tmp3296;
  assign tmp3309 = s7 ? 1 : tmp3310;
  assign tmp3308 = s8 ? tmp3294 : tmp3309;
  assign tmp3307 = s9 ? 1 : tmp3308;
  assign tmp3291 = s10 ? tmp3292 : tmp3307;
  assign tmp3319 = s2 ? tmp3245 : 1;
  assign tmp3318 = s3 ? 1 : tmp3319;
  assign tmp3320 = s3 ? 1 : tmp2988;
  assign tmp3317 = s4 ? tmp3318 : tmp3320;
  assign tmp3316 = s5 ? 1 : tmp3317;
  assign tmp3315 = s6 ? tmp3316 : 1;
  assign tmp3314 = s7 ? 1 : tmp3315;
  assign tmp3324 = s4 ? tmp3318 : 1;
  assign tmp3323 = s5 ? 1 : tmp3324;
  assign tmp3322 = s6 ? 1 : tmp3323;
  assign tmp3321 = s7 ? 1 : tmp3322;
  assign tmp3313 = s8 ? tmp3314 : tmp3321;
  assign tmp3312 = s9 ? 1 : tmp3313;
  assign tmp3328 = s6 ? 1 : tmp3316;
  assign tmp3327 = s7 ? 1 : tmp3328;
  assign tmp3326 = s8 ? tmp3314 : tmp3327;
  assign tmp3325 = s9 ? 1 : tmp3326;
  assign tmp3311 = ~(s10 ? tmp3312 : tmp3325);
  assign tmp3290 = s11 ? tmp3291 : tmp3311;
  assign tmp3339 = ~(s1 ? tmp3136 : tmp2918);
  assign tmp3338 = s2 ? tmp2954 : tmp3339;
  assign tmp3341 = s1 ? tmp3129 : tmp2918;
  assign tmp3340 = ~(s2 ? tmp3341 : tmp2918);
  assign tmp3337 = ~(s3 ? tmp3338 : tmp3340);
  assign tmp3336 = s4 ? tmp3133 : tmp3337;
  assign tmp3335 = s5 ? tmp3128 : tmp3336;
  assign tmp3334 = s6 ? tmp3335 : tmp3142;
  assign tmp3333 = s7 ? tmp3111 : tmp3334;
  assign tmp3346 = ~(s3 ? tmp3338 : tmp3141);
  assign tmp3345 = s4 ? tmp3133 : tmp3346;
  assign tmp3344 = s5 ? tmp3128 : tmp3345;
  assign tmp3343 = s6 ? tmp3161 : tmp3344;
  assign tmp3342 = s7 ? tmp3153 : tmp3343;
  assign tmp3332 = s8 ? tmp3333 : tmp3342;
  assign tmp3331 = s9 ? tmp3100 : tmp3332;
  assign tmp3350 = s6 ? tmp3122 : tmp3335;
  assign tmp3349 = s7 ? tmp3166 : tmp3350;
  assign tmp3348 = s8 ? tmp3333 : tmp3349;
  assign tmp3347 = s9 ? tmp3100 : tmp3348;
  assign tmp3330 = s10 ? tmp3331 : tmp3347;
  assign tmp3329 = ~(s11 ? tmp3017 : tmp3330);
  assign tmp3289 = ~(s12 ? tmp3290 : tmp3329);
  assign tmp3231 = s13 ? tmp3232 : tmp3289;
  assign tmp3168 = s15 ? tmp3169 : tmp3231;
  assign tmp2910 = s16 ? tmp2911 : tmp3168;
  assign s11n = tmp2910;

  assign tmp3357 = ~(l3 ? 1 : 0);
  assign tmp3356 = l2 ? 1 : tmp3357;
  assign tmp3355 = l1 ? tmp3356 : 1;
  assign tmp3358 = l1 ? 1 : tmp3356;
  assign tmp3354 = s11 ? tmp3355 : tmp3358;
  assign tmp3364 = l2 ? 1 : 0;
  assign tmp3363 = l1 ? tmp3356 : tmp3364;
  assign tmp3368 = s1 ? tmp3363 : tmp3358;
  assign tmp3370 = s0 ? tmp3363 : tmp3358;
  assign tmp3371 = s0 ? tmp3363 : tmp3356;
  assign tmp3369 = s1 ? tmp3370 : tmp3371;
  assign tmp3367 = s2 ? tmp3368 : tmp3369;
  assign tmp3375 = l1 ? 1 : tmp3364;
  assign tmp3374 = s0 ? tmp3355 : tmp3375;
  assign tmp3373 = s1 ? tmp3355 : tmp3374;
  assign tmp3372 = s2 ? tmp3373 : tmp3363;
  assign tmp3366 = s3 ? tmp3367 : tmp3372;
  assign tmp3382 = l3 ? 1 : 0;
  assign tmp3381 = l2 ? 1 : tmp3382;
  assign tmp3380 = l1 ? 1 : tmp3381;
  assign tmp3379 = s0 ? tmp3363 : tmp3380;
  assign tmp3384 = l1 ? tmp3356 : tmp3381;
  assign tmp3383 = s0 ? tmp3380 : tmp3384;
  assign tmp3378 = s1 ? tmp3379 : tmp3383;
  assign tmp3385 = s1 ? tmp3363 : tmp3384;
  assign tmp3377 = s2 ? tmp3378 : tmp3385;
  assign tmp3388 = s0 ? tmp3356 : tmp3363;
  assign tmp3387 = s1 ? tmp3388 : tmp3363;
  assign tmp3386 = s2 ? tmp3387 : tmp3379;
  assign tmp3376 = s3 ? tmp3377 : tmp3386;
  assign tmp3365 = s4 ? tmp3366 : tmp3376;
  assign tmp3362 = s5 ? tmp3363 : tmp3365;
  assign tmp3397 = s0 ? tmp3375 : tmp3356;
  assign tmp3396 = s1 ? tmp3397 : tmp3363;
  assign tmp3395 = s2 ? tmp3373 : tmp3396;
  assign tmp3394 = s3 ? tmp3367 : tmp3395;
  assign tmp3401 = s0 ? tmp3384 : tmp3363;
  assign tmp3400 = s1 ? tmp3401 : tmp3384;
  assign tmp3399 = s2 ? tmp3378 : tmp3400;
  assign tmp3404 = s0 ? tmp3375 : tmp3384;
  assign tmp3403 = s1 ? tmp3379 : tmp3404;
  assign tmp3402 = s2 ? tmp3387 : tmp3403;
  assign tmp3398 = s3 ? tmp3399 : tmp3402;
  assign tmp3393 = s4 ? tmp3394 : tmp3398;
  assign tmp3392 = s5 ? tmp3363 : tmp3393;
  assign tmp3391 = s6 ? tmp3392 : tmp3362;
  assign tmp3410 = s1 ? tmp3363 : tmp3371;
  assign tmp3409 = s2 ? tmp3368 : tmp3410;
  assign tmp3412 = s1 ? tmp3355 : tmp3375;
  assign tmp3413 = s1 ? tmp3356 : tmp3363;
  assign tmp3411 = s2 ? tmp3412 : tmp3413;
  assign tmp3408 = s3 ? tmp3409 : tmp3411;
  assign tmp3416 = s1 ? tmp3380 : tmp3384;
  assign tmp3415 = s2 ? tmp3416 : tmp3385;
  assign tmp3414 = s3 ? tmp3415 : tmp3363;
  assign tmp3407 = s4 ? tmp3408 : tmp3414;
  assign tmp3406 = s5 ? tmp3363 : tmp3407;
  assign tmp3421 = s1 ? tmp3397 : tmp3388;
  assign tmp3420 = s2 ? tmp3373 : tmp3421;
  assign tmp3419 = s3 ? tmp3367 : tmp3420;
  assign tmp3425 = s0 ? tmp3356 : tmp3384;
  assign tmp3424 = s1 ? tmp3401 : tmp3425;
  assign tmp3423 = s2 ? tmp3378 : tmp3424;
  assign tmp3426 = s2 ? tmp3388 : tmp3403;
  assign tmp3422 = s3 ? tmp3423 : tmp3426;
  assign tmp3418 = s4 ? tmp3419 : tmp3422;
  assign tmp3417 = s5 ? tmp3363 : tmp3418;
  assign tmp3405 = s6 ? tmp3406 : tmp3417;
  assign tmp3390 = s7 ? tmp3391 : tmp3405;
  assign tmp3431 = s3 ? tmp3409 : tmp3372;
  assign tmp3432 = s3 ? tmp3377 : tmp3363;
  assign tmp3430 = s4 ? tmp3431 : tmp3432;
  assign tmp3429 = s5 ? tmp3363 : tmp3430;
  assign tmp3428 = s6 ? tmp3392 : tmp3429;
  assign tmp3433 = s6 ? tmp3429 : tmp3406;
  assign tmp3427 = s7 ? tmp3428 : tmp3433;
  assign tmp3389 = s8 ? tmp3390 : tmp3427;
  assign tmp3361 = s9 ? tmp3362 : tmp3389;
  assign tmp3437 = s6 ? tmp3362 : tmp3406;
  assign tmp3436 = s7 ? tmp3391 : tmp3437;
  assign tmp3435 = s8 ? tmp3390 : tmp3436;
  assign tmp3434 = s9 ? tmp3362 : tmp3435;
  assign tmp3360 = s10 ? tmp3361 : tmp3434;
  assign tmp3441 = l1 ? tmp3364 : tmp3356;
  assign tmp3445 = s1 ? tmp3441 : tmp3358;
  assign tmp3447 = s0 ? tmp3441 : tmp3358;
  assign tmp3448 = s0 ? tmp3441 : tmp3355;
  assign tmp3446 = s1 ? tmp3447 : tmp3448;
  assign tmp3444 = s2 ? tmp3445 : tmp3446;
  assign tmp3452 = l1 ? tmp3381 : tmp3356;
  assign tmp3451 = s0 ? tmp3355 : tmp3452;
  assign tmp3450 = s1 ? tmp3355 : tmp3451;
  assign tmp3449 = s2 ? tmp3450 : tmp3441;
  assign tmp3443 = s3 ? tmp3444 : tmp3449;
  assign tmp3455 = l1 ? tmp3364 : 1;
  assign tmp3456 = s1 ? tmp3441 : tmp3455;
  assign tmp3454 = s2 ? tmp3455 : tmp3456;
  assign tmp3458 = s0 ? tmp3355 : tmp3441;
  assign tmp3457 = s1 ? tmp3458 : tmp3441;
  assign tmp3453 = s3 ? tmp3454 : tmp3457;
  assign tmp3442 = s4 ? tmp3443 : tmp3453;
  assign tmp3440 = s5 ? tmp3441 : tmp3442;
  assign tmp3467 = s0 ? tmp3452 : tmp3441;
  assign tmp3466 = s1 ? tmp3467 : tmp3441;
  assign tmp3465 = s2 ? tmp3450 : tmp3466;
  assign tmp3464 = s3 ? tmp3444 : tmp3465;
  assign tmp3471 = s0 ? tmp3356 : tmp3355;
  assign tmp3472 = s0 ? tmp3355 : tmp3455;
  assign tmp3470 = s1 ? tmp3471 : tmp3472;
  assign tmp3469 = s2 ? tmp3470 : tmp3456;
  assign tmp3475 = s0 ? tmp3452 : tmp3455;
  assign tmp3474 = s1 ? tmp3471 : tmp3475;
  assign tmp3473 = s2 ? tmp3457 : tmp3474;
  assign tmp3468 = s3 ? tmp3469 : tmp3473;
  assign tmp3463 = s4 ? tmp3464 : tmp3468;
  assign tmp3462 = s5 ? tmp3441 : tmp3463;
  assign tmp3480 = s1 ? tmp3355 : tmp3455;
  assign tmp3479 = s2 ? tmp3480 : tmp3456;
  assign tmp3478 = s3 ? tmp3479 : tmp3457;
  assign tmp3477 = s4 ? tmp3443 : tmp3478;
  assign tmp3476 = s5 ? tmp3441 : tmp3477;
  assign tmp3461 = s6 ? tmp3462 : tmp3476;
  assign tmp3486 = s1 ? tmp3441 : tmp3448;
  assign tmp3485 = s2 ? tmp3445 : tmp3486;
  assign tmp3488 = s1 ? tmp3355 : tmp3452;
  assign tmp3489 = s1 ? tmp3441 : tmp3356;
  assign tmp3487 = s2 ? tmp3488 : tmp3489;
  assign tmp3484 = s3 ? tmp3485 : tmp3487;
  assign tmp3491 = s2 ? tmp3480 : tmp3441;
  assign tmp3490 = s3 ? tmp3491 : tmp3441;
  assign tmp3483 = s4 ? tmp3484 : tmp3490;
  assign tmp3482 = s5 ? tmp3441 : tmp3483;
  assign tmp3497 = s0 ? tmp3441 : tmp3356;
  assign tmp3496 = s1 ? tmp3467 : tmp3497;
  assign tmp3495 = s2 ? tmp3450 : tmp3496;
  assign tmp3494 = s3 ? tmp3444 : tmp3495;
  assign tmp3500 = s1 ? tmp3441 : tmp3472;
  assign tmp3499 = s2 ? tmp3470 : tmp3500;
  assign tmp3498 = s3 ? tmp3499 : tmp3473;
  assign tmp3493 = s4 ? tmp3494 : tmp3498;
  assign tmp3492 = s5 ? tmp3441 : tmp3493;
  assign tmp3481 = s6 ? tmp3482 : tmp3492;
  assign tmp3460 = s7 ? tmp3461 : tmp3481;
  assign tmp3507 = s1 ? tmp3356 : tmp3455;
  assign tmp3506 = s2 ? tmp3507 : tmp3456;
  assign tmp3509 = s1 ? tmp3356 : tmp3475;
  assign tmp3508 = s2 ? tmp3457 : tmp3509;
  assign tmp3505 = s3 ? tmp3506 : tmp3508;
  assign tmp3504 = s4 ? tmp3464 : tmp3505;
  assign tmp3503 = s5 ? tmp3441 : tmp3504;
  assign tmp3512 = s3 ? tmp3485 : tmp3449;
  assign tmp3514 = s2 ? tmp3455 : tmp3441;
  assign tmp3513 = s3 ? tmp3514 : tmp3441;
  assign tmp3511 = s4 ? tmp3512 : tmp3513;
  assign tmp3510 = s5 ? tmp3441 : tmp3511;
  assign tmp3502 = s6 ? tmp3503 : tmp3510;
  assign tmp3517 = s4 ? tmp3512 : tmp3490;
  assign tmp3516 = s5 ? tmp3441 : tmp3517;
  assign tmp3515 = s6 ? tmp3516 : tmp3482;
  assign tmp3501 = s7 ? tmp3502 : tmp3515;
  assign tmp3459 = s8 ? tmp3460 : tmp3501;
  assign tmp3439 = s9 ? tmp3440 : tmp3459;
  assign tmp3521 = s6 ? tmp3503 : tmp3440;
  assign tmp3522 = s6 ? tmp3476 : tmp3482;
  assign tmp3520 = s7 ? tmp3521 : tmp3522;
  assign tmp3519 = s8 ? tmp3460 : tmp3520;
  assign tmp3518 = s9 ? tmp3440 : tmp3519;
  assign tmp3438 = s10 ? tmp3439 : tmp3518;
  assign tmp3359 = s11 ? tmp3360 : tmp3438;
  assign tmp3353 = s12 ? tmp3354 : tmp3359;
  assign tmp3524 = s11 ? tmp3380 : tmp3355;
  assign tmp3530 = l1 ? tmp3381 : tmp3364;
  assign tmp3532 = s0 ? tmp3375 : tmp3530;
  assign tmp3531 = s1 ? tmp3530 : tmp3532;
  assign tmp3529 = s2 ? tmp3530 : tmp3531;
  assign tmp3536 = s1 ? tmp3532 : tmp3375;
  assign tmp3537 = s0 ? tmp3530 : tmp3375;
  assign tmp3535 = s2 ? tmp3536 : tmp3537;
  assign tmp3539 = s1 ? tmp3381 : tmp3530;
  assign tmp3540 = s1 ? tmp3530 : tmp3375;
  assign tmp3538 = s2 ? tmp3539 : tmp3540;
  assign tmp3534 = s3 ? tmp3535 : tmp3538;
  assign tmp3544 = s0 ? tmp3380 : tmp3381;
  assign tmp3543 = s1 ? tmp3380 : tmp3544;
  assign tmp3545 = s1 ? tmp3530 : tmp3381;
  assign tmp3542 = s2 ? tmp3543 : tmp3545;
  assign tmp3547 = s1 ? tmp3380 : tmp3530;
  assign tmp3546 = s2 ? tmp3530 : tmp3547;
  assign tmp3541 = s3 ? tmp3542 : tmp3546;
  assign tmp3533 = s4 ? tmp3534 : tmp3541;
  assign tmp3528 = s5 ? tmp3529 : tmp3533;
  assign tmp3556 = s0 ? tmp3530 : tmp3358;
  assign tmp3555 = s1 ? tmp3537 : tmp3556;
  assign tmp3554 = s2 ? tmp3536 : tmp3555;
  assign tmp3559 = s0 ? tmp3358 : tmp3380;
  assign tmp3560 = s0 ? tmp3380 : tmp3530;
  assign tmp3558 = s1 ? tmp3559 : tmp3560;
  assign tmp3561 = s1 ? tmp3530 : tmp3537;
  assign tmp3557 = s2 ? tmp3558 : tmp3561;
  assign tmp3553 = s3 ? tmp3554 : tmp3557;
  assign tmp3565 = s0 ? tmp3375 : tmp3380;
  assign tmp3564 = s1 ? tmp3565 : tmp3544;
  assign tmp3567 = s0 ? tmp3381 : tmp3530;
  assign tmp3568 = s0 ? tmp3358 : tmp3381;
  assign tmp3566 = s1 ? tmp3567 : tmp3568;
  assign tmp3563 = s2 ? tmp3564 : tmp3566;
  assign tmp3570 = s1 ? tmp3560 : tmp3530;
  assign tmp3572 = s0 ? tmp3530 : tmp3381;
  assign tmp3571 = s1 ? tmp3565 : tmp3572;
  assign tmp3569 = s2 ? tmp3570 : tmp3571;
  assign tmp3562 = s3 ? tmp3563 : tmp3569;
  assign tmp3552 = s4 ? tmp3553 : tmp3562;
  assign tmp3551 = s5 ? tmp3529 : tmp3552;
  assign tmp3576 = s2 ? tmp3547 : tmp3540;
  assign tmp3575 = s3 ? tmp3554 : tmp3576;
  assign tmp3574 = s4 ? tmp3575 : tmp3541;
  assign tmp3573 = s5 ? tmp3529 : tmp3574;
  assign tmp3550 = s6 ? tmp3551 : tmp3573;
  assign tmp3582 = s1 ? tmp3532 : tmp3358;
  assign tmp3583 = s1 ? tmp3530 : tmp3556;
  assign tmp3581 = s2 ? tmp3582 : tmp3583;
  assign tmp3586 = s0 ? tmp3530 : tmp3452;
  assign tmp3585 = s1 ? tmp3586 : tmp3375;
  assign tmp3584 = s2 ? tmp3547 : tmp3585;
  assign tmp3580 = s3 ? tmp3581 : tmp3584;
  assign tmp3589 = s1 ? tmp3380 : tmp3381;
  assign tmp3588 = s2 ? tmp3589 : tmp3545;
  assign tmp3587 = s3 ? tmp3588 : tmp3530;
  assign tmp3579 = s4 ? tmp3580 : tmp3587;
  assign tmp3578 = s5 ? tmp3529 : tmp3579;
  assign tmp3593 = s2 ? tmp3582 : tmp3555;
  assign tmp3596 = s0 ? tmp3452 : tmp3375;
  assign tmp3595 = s1 ? tmp3586 : tmp3596;
  assign tmp3594 = s2 ? tmp3558 : tmp3595;
  assign tmp3592 = s3 ? tmp3593 : tmp3594;
  assign tmp3600 = s0 ? tmp3452 : tmp3530;
  assign tmp3599 = s1 ? tmp3560 : tmp3600;
  assign tmp3598 = s2 ? tmp3599 : tmp3571;
  assign tmp3597 = s3 ? tmp3563 : tmp3598;
  assign tmp3591 = s4 ? tmp3592 : tmp3597;
  assign tmp3590 = s5 ? tmp3529 : tmp3591;
  assign tmp3577 = s6 ? tmp3578 : tmp3590;
  assign tmp3549 = s7 ? tmp3550 : tmp3577;
  assign tmp3607 = s1 ? tmp3381 : tmp3567;
  assign tmp3606 = s2 ? tmp3607 : tmp3561;
  assign tmp3605 = s3 ? tmp3535 : tmp3606;
  assign tmp3610 = s1 ? tmp3567 : tmp3381;
  assign tmp3609 = s2 ? tmp3564 : tmp3610;
  assign tmp3612 = s1 ? tmp3567 : tmp3530;
  assign tmp3611 = s2 ? tmp3612 : tmp3571;
  assign tmp3608 = s3 ? tmp3609 : tmp3611;
  assign tmp3604 = s4 ? tmp3605 : tmp3608;
  assign tmp3603 = s5 ? tmp3529 : tmp3604;
  assign tmp3617 = s1 ? tmp3530 : tmp3572;
  assign tmp3616 = s2 ? tmp3536 : tmp3617;
  assign tmp3615 = s3 ? tmp3616 : tmp3538;
  assign tmp3618 = s3 ? tmp3542 : tmp3530;
  assign tmp3614 = s4 ? tmp3615 : tmp3618;
  assign tmp3613 = s5 ? tmp3529 : tmp3614;
  assign tmp3602 = s6 ? tmp3603 : tmp3613;
  assign tmp3623 = s2 ? tmp3536 : tmp3583;
  assign tmp3622 = s3 ? tmp3623 : tmp3576;
  assign tmp3621 = s4 ? tmp3622 : tmp3618;
  assign tmp3620 = s5 ? tmp3529 : tmp3621;
  assign tmp3619 = s6 ? tmp3620 : tmp3578;
  assign tmp3601 = s7 ? tmp3602 : tmp3619;
  assign tmp3548 = s8 ? tmp3549 : tmp3601;
  assign tmp3527 = s9 ? tmp3528 : tmp3548;
  assign tmp3627 = s6 ? tmp3603 : tmp3528;
  assign tmp3628 = s6 ? tmp3573 : tmp3578;
  assign tmp3626 = s7 ? tmp3627 : tmp3628;
  assign tmp3625 = s8 ? tmp3549 : tmp3626;
  assign tmp3624 = s9 ? tmp3528 : tmp3625;
  assign tmp3526 = s10 ? tmp3527 : tmp3624;
  assign tmp3632 = l1 ? tmp3364 : tmp3381;
  assign tmp3636 = s1 ? tmp3632 : tmp3381;
  assign tmp3638 = s0 ? tmp3632 : tmp3455;
  assign tmp3637 = s1 ? tmp3632 : tmp3638;
  assign tmp3635 = s2 ? tmp3636 : tmp3637;
  assign tmp3641 = s0 ? tmp3355 : tmp3381;
  assign tmp3640 = s1 ? tmp3355 : tmp3641;
  assign tmp3642 = s1 ? tmp3455 : tmp3632;
  assign tmp3639 = s2 ? tmp3640 : tmp3642;
  assign tmp3634 = s3 ? tmp3635 : tmp3639;
  assign tmp3646 = s0 ? tmp3380 : tmp3632;
  assign tmp3645 = s1 ? tmp3380 : tmp3646;
  assign tmp3648 = s0 ? tmp3455 : tmp3632;
  assign tmp3647 = s1 ? tmp3632 : tmp3648;
  assign tmp3644 = s2 ? tmp3645 : tmp3647;
  assign tmp3650 = s1 ? tmp3648 : tmp3632;
  assign tmp3651 = s1 ? tmp3380 : tmp3632;
  assign tmp3649 = s2 ? tmp3650 : tmp3651;
  assign tmp3643 = s3 ? tmp3644 : tmp3649;
  assign tmp3633 = s4 ? tmp3634 : tmp3643;
  assign tmp3631 = s5 ? tmp3632 : tmp3633;
  assign tmp3659 = s1 ? tmp3632 : tmp3355;
  assign tmp3661 = s0 ? tmp3632 : tmp3355;
  assign tmp3660 = s1 ? tmp3661 : tmp3638;
  assign tmp3658 = s2 ? tmp3659 : tmp3660;
  assign tmp3664 = s0 ? tmp3381 : tmp3455;
  assign tmp3663 = s1 ? tmp3664 : tmp3648;
  assign tmp3662 = s2 ? tmp3640 : tmp3663;
  assign tmp3657 = s3 ? tmp3658 : tmp3662;
  assign tmp3668 = s0 ? tmp3384 : tmp3380;
  assign tmp3667 = s1 ? tmp3668 : tmp3646;
  assign tmp3666 = s2 ? tmp3667 : tmp3647;
  assign tmp3671 = s0 ? tmp3381 : tmp3632;
  assign tmp3670 = s1 ? tmp3668 : tmp3671;
  assign tmp3669 = s2 ? tmp3650 : tmp3670;
  assign tmp3665 = s3 ? tmp3666 : tmp3669;
  assign tmp3656 = s4 ? tmp3657 : tmp3665;
  assign tmp3655 = s5 ? tmp3632 : tmp3656;
  assign tmp3675 = s2 ? tmp3659 : tmp3637;
  assign tmp3674 = s3 ? tmp3675 : tmp3639;
  assign tmp3673 = s4 ? tmp3674 : tmp3643;
  assign tmp3672 = s5 ? tmp3632 : tmp3673;
  assign tmp3654 = s6 ? tmp3655 : tmp3672;
  assign tmp3682 = s0 ? tmp3384 : tmp3632;
  assign tmp3681 = s1 ? tmp3682 : tmp3355;
  assign tmp3683 = s1 ? tmp3632 : tmp3661;
  assign tmp3680 = s2 ? tmp3681 : tmp3683;
  assign tmp3685 = s1 ? tmp3355 : tmp3381;
  assign tmp3686 = s1 ? tmp3455 : tmp3384;
  assign tmp3684 = s2 ? tmp3685 : tmp3686;
  assign tmp3679 = s3 ? tmp3680 : tmp3684;
  assign tmp3688 = s2 ? tmp3651 : tmp3632;
  assign tmp3687 = s3 ? tmp3688 : tmp3632;
  assign tmp3678 = s4 ? tmp3679 : tmp3687;
  assign tmp3677 = s5 ? tmp3632 : tmp3678;
  assign tmp3692 = s2 ? tmp3681 : tmp3661;
  assign tmp3695 = s0 ? tmp3455 : tmp3384;
  assign tmp3694 = s1 ? tmp3664 : tmp3695;
  assign tmp3693 = s2 ? tmp3640 : tmp3694;
  assign tmp3691 = s3 ? tmp3692 : tmp3693;
  assign tmp3699 = s0 ? tmp3355 : tmp3632;
  assign tmp3698 = s1 ? tmp3632 : tmp3699;
  assign tmp3697 = s2 ? tmp3667 : tmp3698;
  assign tmp3701 = s1 ? tmp3699 : tmp3648;
  assign tmp3700 = s2 ? tmp3701 : tmp3670;
  assign tmp3696 = s3 ? tmp3697 : tmp3700;
  assign tmp3690 = s4 ? tmp3691 : tmp3696;
  assign tmp3689 = s5 ? tmp3632 : tmp3690;
  assign tmp3676 = s6 ? tmp3677 : tmp3689;
  assign tmp3653 = s7 ? tmp3654 : tmp3676;
  assign tmp3709 = s0 ? tmp3632 : tmp3381;
  assign tmp3708 = s1 ? tmp3709 : tmp3638;
  assign tmp3707 = s2 ? tmp3636 : tmp3708;
  assign tmp3706 = s3 ? tmp3707 : tmp3662;
  assign tmp3705 = s4 ? tmp3706 : tmp3665;
  assign tmp3704 = s5 ? tmp3632 : tmp3705;
  assign tmp3713 = s2 ? tmp3645 : tmp3632;
  assign tmp3712 = s3 ? tmp3713 : tmp3632;
  assign tmp3711 = s4 ? tmp3634 : tmp3712;
  assign tmp3710 = s5 ? tmp3632 : tmp3711;
  assign tmp3703 = s6 ? tmp3704 : tmp3710;
  assign tmp3716 = s4 ? tmp3674 : tmp3712;
  assign tmp3715 = s5 ? tmp3632 : tmp3716;
  assign tmp3714 = s6 ? tmp3715 : tmp3677;
  assign tmp3702 = s7 ? tmp3703 : tmp3714;
  assign tmp3652 = s8 ? tmp3653 : tmp3702;
  assign tmp3630 = s9 ? tmp3631 : tmp3652;
  assign tmp3720 = s6 ? tmp3704 : tmp3631;
  assign tmp3721 = s6 ? tmp3672 : tmp3677;
  assign tmp3719 = s7 ? tmp3720 : tmp3721;
  assign tmp3718 = s8 ? tmp3653 : tmp3719;
  assign tmp3717 = s9 ? tmp3631 : tmp3718;
  assign tmp3629 = s10 ? tmp3630 : tmp3717;
  assign tmp3525 = s11 ? tmp3526 : tmp3629;
  assign tmp3523 = s12 ? tmp3524 : tmp3525;
  assign tmp3352 = s13 ? tmp3353 : tmp3523;
  assign tmp3732 = s1 ? tmp3356 : tmp3358;
  assign tmp3731 = s2 ? tmp3732 : tmp3356;
  assign tmp3734 = s1 ? tmp3355 : tmp3358;
  assign tmp3733 = s2 ? tmp3734 : tmp3356;
  assign tmp3730 = s3 ? tmp3731 : tmp3733;
  assign tmp3737 = s1 ? tmp3358 : tmp3356;
  assign tmp3736 = s2 ? tmp3737 : tmp3356;
  assign tmp3735 = s3 ? tmp3736 : tmp3356;
  assign tmp3729 = s4 ? tmp3730 : tmp3735;
  assign tmp3728 = s5 ? tmp3356 : tmp3729;
  assign tmp3745 = s1 ? tmp3380 : tmp3356;
  assign tmp3744 = s2 ? tmp3745 : tmp3356;
  assign tmp3743 = s3 ? tmp3744 : tmp3356;
  assign tmp3742 = s4 ? tmp3730 : tmp3743;
  assign tmp3741 = s5 ? tmp3356 : tmp3742;
  assign tmp3751 = s0 ? tmp3356 : tmp3358;
  assign tmp3750 = s1 ? tmp3751 : tmp3356;
  assign tmp3749 = s2 ? tmp3732 : tmp3750;
  assign tmp3754 = s0 ? tmp3355 : tmp3358;
  assign tmp3753 = s1 ? tmp3355 : tmp3754;
  assign tmp3752 = s2 ? tmp3753 : tmp3356;
  assign tmp3748 = s3 ? tmp3749 : tmp3752;
  assign tmp3758 = s0 ? tmp3356 : tmp3380;
  assign tmp3759 = s0 ? tmp3380 : tmp3356;
  assign tmp3757 = s1 ? tmp3758 : tmp3759;
  assign tmp3756 = s2 ? tmp3757 : tmp3356;
  assign tmp3760 = s2 ? tmp3356 : tmp3758;
  assign tmp3755 = s3 ? tmp3756 : tmp3760;
  assign tmp3747 = s4 ? tmp3748 : tmp3755;
  assign tmp3746 = s5 ? tmp3356 : tmp3747;
  assign tmp3740 = s6 ? tmp3741 : tmp3746;
  assign tmp3739 = s7 ? tmp3391 : tmp3740;
  assign tmp3765 = s3 ? tmp3731 : tmp3752;
  assign tmp3769 = s0 ? tmp3358 : tmp3356;
  assign tmp3768 = s1 ? tmp3751 : tmp3769;
  assign tmp3767 = s2 ? tmp3768 : tmp3356;
  assign tmp3766 = s3 ? tmp3767 : tmp3356;
  assign tmp3764 = s4 ? tmp3765 : tmp3766;
  assign tmp3763 = s5 ? tmp3356 : tmp3764;
  assign tmp3762 = s6 ? tmp3763 : tmp3728;
  assign tmp3770 = s6 ? tmp3429 : tmp3741;
  assign tmp3761 = s7 ? tmp3762 : tmp3770;
  assign tmp3738 = s8 ? tmp3739 : tmp3761;
  assign tmp3727 = s9 ? tmp3728 : tmp3738;
  assign tmp3778 = s2 ? tmp3356 : tmp3751;
  assign tmp3777 = s3 ? tmp3767 : tmp3778;
  assign tmp3776 = s4 ? tmp3748 : tmp3777;
  assign tmp3775 = s5 ? tmp3356 : tmp3776;
  assign tmp3774 = s6 ? tmp3775 : tmp3728;
  assign tmp3779 = s6 ? tmp3362 : tmp3741;
  assign tmp3773 = s7 ? tmp3774 : tmp3779;
  assign tmp3772 = s8 ? tmp3739 : tmp3773;
  assign tmp3771 = s9 ? tmp3728 : tmp3772;
  assign tmp3726 = s10 ? tmp3727 : tmp3771;
  assign tmp3782 = l1 ? tmp3381 : 1;
  assign tmp3790 = s1 ? tmp3782 : tmp3355;
  assign tmp3792 = s0 ? tmp3782 : tmp3355;
  assign tmp3791 = s1 ? tmp3782 : tmp3792;
  assign tmp3789 = s2 ? tmp3790 : tmp3791;
  assign tmp3794 = s1 ? tmp3355 : tmp3782;
  assign tmp3793 = s2 ? tmp3794 : tmp3790;
  assign tmp3788 = s3 ? tmp3789 : tmp3793;
  assign tmp3796 = s2 ? tmp3794 : tmp3782;
  assign tmp3795 = s3 ? tmp3796 : tmp3782;
  assign tmp3787 = s4 ? tmp3788 : tmp3795;
  assign tmp3786 = s5 ? tmp3782 : tmp3787;
  assign tmp3800 = s2 ? tmp3790 : tmp3792;
  assign tmp3803 = s0 ? tmp3355 : tmp3782;
  assign tmp3802 = s1 ? tmp3355 : tmp3803;
  assign tmp3801 = s2 ? tmp3802 : tmp3791;
  assign tmp3799 = s3 ? tmp3800 : tmp3801;
  assign tmp3806 = s1 ? tmp3782 : tmp3803;
  assign tmp3805 = s2 ? tmp3802 : tmp3806;
  assign tmp3808 = s1 ? tmp3803 : tmp3782;
  assign tmp3807 = s2 ? tmp3808 : tmp3794;
  assign tmp3804 = s3 ? tmp3805 : tmp3807;
  assign tmp3798 = s4 ? tmp3799 : tmp3804;
  assign tmp3797 = s5 ? tmp3782 : tmp3798;
  assign tmp3785 = s6 ? tmp3786 : tmp3797;
  assign tmp3784 = s7 ? tmp3461 : tmp3785;
  assign tmp3810 = s6 ? tmp3516 : tmp3786;
  assign tmp3809 = s7 ? tmp3782 : tmp3810;
  assign tmp3783 = s8 ? tmp3784 : tmp3809;
  assign tmp3781 = s9 ? tmp3782 : tmp3783;
  assign tmp3814 = s6 ? tmp3476 : tmp3786;
  assign tmp3813 = s7 ? tmp3782 : tmp3814;
  assign tmp3812 = s8 ? tmp3784 : tmp3813;
  assign tmp3811 = s9 ? tmp3782 : tmp3812;
  assign tmp3780 = s10 ? tmp3781 : tmp3811;
  assign tmp3725 = s11 ? tmp3726 : tmp3780;
  assign tmp3724 = s12 ? tmp3354 : tmp3725;
  assign tmp3824 = s1 ? tmp3452 : tmp3568;
  assign tmp3823 = s2 ? tmp3452 : tmp3824;
  assign tmp3829 = s0 ? tmp3380 : tmp3452;
  assign tmp3828 = s1 ? tmp3829 : tmp3358;
  assign tmp3831 = s0 ? tmp3452 : tmp3358;
  assign tmp3830 = s1 ? tmp3452 : tmp3831;
  assign tmp3827 = s2 ? tmp3828 : tmp3830;
  assign tmp3833 = s1 ? tmp3380 : tmp3782;
  assign tmp3834 = s1 ? tmp3782 : tmp3380;
  assign tmp3832 = s2 ? tmp3833 : tmp3834;
  assign tmp3826 = s3 ? tmp3827 : tmp3832;
  assign tmp3837 = s1 ? tmp3452 : tmp3381;
  assign tmp3836 = s2 ? tmp3833 : tmp3837;
  assign tmp3835 = s3 ? tmp3836 : tmp3837;
  assign tmp3825 = s4 ? tmp3826 : tmp3835;
  assign tmp3822 = s5 ? tmp3823 : tmp3825;
  assign tmp3841 = s2 ? tmp3828 : tmp3831;
  assign tmp3844 = s0 ? tmp3380 : tmp3782;
  assign tmp3843 = s1 ? tmp3559 : tmp3844;
  assign tmp3846 = s0 ? tmp3782 : tmp3380;
  assign tmp3845 = s1 ? tmp3782 : tmp3846;
  assign tmp3842 = s2 ? tmp3843 : tmp3845;
  assign tmp3840 = s3 ? tmp3841 : tmp3842;
  assign tmp3849 = s1 ? tmp3380 : tmp3844;
  assign tmp3851 = s0 ? tmp3381 : tmp3452;
  assign tmp3850 = s1 ? tmp3851 : tmp3568;
  assign tmp3848 = s2 ? tmp3849 : tmp3850;
  assign tmp3854 = s0 ? tmp3452 : tmp3381;
  assign tmp3853 = s1 ? tmp3844 : tmp3854;
  assign tmp3852 = s2 ? tmp3853 : tmp3833;
  assign tmp3847 = s3 ? tmp3848 : tmp3852;
  assign tmp3839 = s4 ? tmp3840 : tmp3847;
  assign tmp3838 = s5 ? tmp3823 : tmp3839;
  assign tmp3821 = s6 ? tmp3822 : tmp3838;
  assign tmp3820 = s7 ? tmp3550 : tmp3821;
  assign tmp3856 = s6 ? tmp3620 : tmp3822;
  assign tmp3855 = s7 ? tmp3782 : tmp3856;
  assign tmp3819 = s8 ? tmp3820 : tmp3855;
  assign tmp3818 = s9 ? tmp3782 : tmp3819;
  assign tmp3860 = s6 ? tmp3573 : tmp3822;
  assign tmp3859 = s7 ? tmp3782 : tmp3860;
  assign tmp3858 = s8 ? tmp3820 : tmp3859;
  assign tmp3857 = s9 ? tmp3782 : tmp3858;
  assign tmp3817 = s10 ? tmp3818 : tmp3857;
  assign tmp3864 = s7 ? tmp3654 : tmp3785;
  assign tmp3866 = s6 ? tmp3715 : tmp3786;
  assign tmp3865 = s7 ? tmp3782 : tmp3866;
  assign tmp3863 = s8 ? tmp3864 : tmp3865;
  assign tmp3862 = s9 ? tmp3782 : tmp3863;
  assign tmp3870 = s6 ? tmp3672 : tmp3786;
  assign tmp3869 = s7 ? tmp3782 : tmp3870;
  assign tmp3868 = s8 ? tmp3864 : tmp3869;
  assign tmp3867 = s9 ? tmp3782 : tmp3868;
  assign tmp3861 = s10 ? tmp3862 : tmp3867;
  assign tmp3816 = s11 ? tmp3817 : tmp3861;
  assign tmp3815 = s12 ? tmp3524 : tmp3816;
  assign tmp3723 = s13 ? tmp3724 : tmp3815;
  assign tmp3886 = l2 ? tmp3382 : 0;
  assign tmp3885 = l1 ? tmp3382 : tmp3886;
  assign tmp3887 = ~(l1 ? tmp3356 : 1);
  assign tmp3884 = s0 ? tmp3885 : tmp3887;
  assign tmp3883 = s1 ? tmp3884 : tmp3887;
  assign tmp3882 = ~(s2 ? tmp3883 : tmp3887);
  assign tmp3881 = s3 ? tmp3355 : tmp3882;
  assign tmp3891 = ~(s0 ? tmp3885 : tmp3887);
  assign tmp3890 = s1 ? tmp3355 : tmp3891;
  assign tmp3889 = s2 ? tmp3355 : tmp3890;
  assign tmp3888 = s3 ? tmp3889 : tmp3355;
  assign tmp3880 = s4 ? tmp3881 : tmp3888;
  assign tmp3879 = s5 ? tmp3355 : tmp3880;
  assign tmp3878 = s6 ? tmp3879 : tmp3355;
  assign tmp3877 = s7 ? tmp3355 : tmp3878;
  assign tmp3895 = s4 ? tmp3881 : tmp3355;
  assign tmp3894 = s5 ? tmp3355 : tmp3895;
  assign tmp3893 = s6 ? tmp3355 : tmp3894;
  assign tmp3892 = s7 ? tmp3355 : tmp3893;
  assign tmp3876 = s8 ? tmp3877 : tmp3892;
  assign tmp3875 = s9 ? tmp3355 : tmp3876;
  assign tmp3899 = s6 ? tmp3355 : tmp3879;
  assign tmp3898 = s7 ? tmp3355 : tmp3899;
  assign tmp3897 = s8 ? tmp3877 : tmp3898;
  assign tmp3896 = s9 ? tmp3355 : tmp3897;
  assign tmp3874 = s10 ? tmp3875 : tmp3896;
  assign tmp3911 = ~(l1 ? tmp3886 : tmp3382);
  assign tmp3910 = s0 ? tmp3358 : tmp3911;
  assign tmp3909 = s1 ? tmp3358 : tmp3910;
  assign tmp3912 = s1 ? tmp3910 : tmp3358;
  assign tmp3908 = s2 ? tmp3909 : tmp3912;
  assign tmp3907 = s3 ? tmp3908 : tmp3358;
  assign tmp3906 = s4 ? tmp3907 : tmp3358;
  assign tmp3905 = s5 ? tmp3358 : tmp3906;
  assign tmp3904 = s6 ? tmp3905 : tmp3358;
  assign tmp3903 = s7 ? tmp3358 : tmp3904;
  assign tmp3918 = s2 ? tmp3909 : tmp3358;
  assign tmp3917 = s3 ? tmp3918 : tmp3358;
  assign tmp3916 = s4 ? tmp3917 : tmp3358;
  assign tmp3915 = s5 ? tmp3358 : tmp3916;
  assign tmp3914 = s6 ? tmp3358 : tmp3915;
  assign tmp3913 = s7 ? tmp3358 : tmp3914;
  assign tmp3902 = s8 ? tmp3903 : tmp3913;
  assign tmp3901 = s9 ? tmp3358 : tmp3902;
  assign tmp3922 = s6 ? tmp3358 : tmp3905;
  assign tmp3921 = s7 ? tmp3358 : tmp3922;
  assign tmp3920 = s8 ? tmp3903 : tmp3921;
  assign tmp3919 = s9 ? tmp3358 : tmp3920;
  assign tmp3900 = s10 ? tmp3901 : tmp3919;
  assign tmp3873 = s11 ? tmp3874 : tmp3900;
  assign tmp3936 = ~(l2 ? tmp3382 : 0);
  assign tmp3935 = l1 ? tmp3382 : tmp3936;
  assign tmp3937 = ~(l1 ? 1 : tmp3381);
  assign tmp3934 = s0 ? tmp3935 : tmp3937;
  assign tmp3938 = ~(l1 ? tmp3356 : tmp3381);
  assign tmp3933 = s1 ? tmp3934 : tmp3938;
  assign tmp3939 = ~(s1 ? tmp3363 : tmp3384);
  assign tmp3932 = s2 ? tmp3933 : tmp3939;
  assign tmp3941 = ~(l1 ? tmp3382 : tmp3936);
  assign tmp3940 = ~(s2 ? tmp3363 : tmp3941);
  assign tmp3931 = ~(s3 ? tmp3932 : tmp3940);
  assign tmp3930 = s4 ? tmp3408 : tmp3931;
  assign tmp3929 = s5 ? tmp3363 : tmp3930;
  assign tmp3928 = s6 ? tmp3929 : tmp3417;
  assign tmp3927 = s7 ? tmp3391 : tmp3928;
  assign tmp3947 = ~(l1 ? tmp3356 : tmp3364);
  assign tmp3946 = ~(s3 ? tmp3932 : tmp3947);
  assign tmp3945 = s4 ? tmp3408 : tmp3946;
  assign tmp3944 = s5 ? tmp3363 : tmp3945;
  assign tmp3943 = s6 ? tmp3429 : tmp3944;
  assign tmp3942 = s7 ? tmp3428 : tmp3943;
  assign tmp3926 = s8 ? tmp3927 : tmp3942;
  assign tmp3925 = s9 ? tmp3362 : tmp3926;
  assign tmp3951 = s6 ? tmp3362 : tmp3929;
  assign tmp3950 = s7 ? tmp3391 : tmp3951;
  assign tmp3949 = s8 ? tmp3927 : tmp3950;
  assign tmp3948 = s9 ? tmp3362 : tmp3949;
  assign tmp3924 = s10 ? tmp3925 : tmp3948;
  assign tmp3963 = l1 ? tmp3364 : tmp3357;
  assign tmp3962 = s0 ? tmp3963 : tmp3356;
  assign tmp3961 = s1 ? tmp3441 : tmp3962;
  assign tmp3960 = s2 ? tmp3488 : tmp3961;
  assign tmp3959 = s3 ? tmp3485 : tmp3960;
  assign tmp3966 = s0 ? tmp3963 : tmp3441;
  assign tmp3965 = s1 ? tmp3441 : tmp3966;
  assign tmp3964 = s3 ? tmp3491 : tmp3965;
  assign tmp3958 = s4 ? tmp3959 : tmp3964;
  assign tmp3957 = s5 ? tmp3441 : tmp3958;
  assign tmp3956 = s6 ? tmp3957 : tmp3492;
  assign tmp3955 = s7 ? tmp3461 : tmp3956;
  assign tmp3970 = s4 ? tmp3959 : tmp3490;
  assign tmp3969 = s5 ? tmp3441 : tmp3970;
  assign tmp3968 = s6 ? tmp3516 : tmp3969;
  assign tmp3967 = s7 ? tmp3502 : tmp3968;
  assign tmp3954 = s8 ? tmp3955 : tmp3967;
  assign tmp3953 = s9 ? tmp3440 : tmp3954;
  assign tmp3974 = s6 ? tmp3476 : tmp3957;
  assign tmp3973 = s7 ? tmp3521 : tmp3974;
  assign tmp3972 = s8 ? tmp3955 : tmp3973;
  assign tmp3971 = s9 ? tmp3440 : tmp3972;
  assign tmp3952 = s10 ? tmp3953 : tmp3971;
  assign tmp3923 = s11 ? tmp3924 : tmp3952;
  assign tmp3872 = s12 ? tmp3873 : tmp3923;
  assign tmp3989 = l2 ? tmp3382 : 1;
  assign tmp3988 = l1 ? tmp3989 : tmp3382;
  assign tmp3987 = s0 ? tmp3988 : tmp3380;
  assign tmp3986 = s1 ? tmp3380 : tmp3987;
  assign tmp3985 = s2 ? tmp3986 : tmp3380;
  assign tmp3990 = s2 ? tmp3380 : tmp3988;
  assign tmp3984 = s3 ? tmp3985 : tmp3990;
  assign tmp3983 = s4 ? tmp3380 : tmp3984;
  assign tmp3982 = s5 ? tmp3380 : tmp3983;
  assign tmp3981 = s6 ? tmp3982 : tmp3380;
  assign tmp3980 = s7 ? tmp3380 : tmp3981;
  assign tmp3995 = s3 ? tmp3985 : tmp3380;
  assign tmp3994 = s4 ? tmp3380 : tmp3995;
  assign tmp3993 = s5 ? tmp3380 : tmp3994;
  assign tmp3992 = s6 ? tmp3380 : tmp3993;
  assign tmp3991 = s7 ? tmp3380 : tmp3992;
  assign tmp3979 = s8 ? tmp3980 : tmp3991;
  assign tmp3978 = s9 ? tmp3380 : tmp3979;
  assign tmp3999 = s6 ? tmp3380 : tmp3982;
  assign tmp3998 = s7 ? tmp3380 : tmp3999;
  assign tmp3997 = s8 ? tmp3980 : tmp3998;
  assign tmp3996 = s9 ? tmp3380 : tmp3997;
  assign tmp3977 = s10 ? tmp3978 : tmp3996;
  assign tmp4012 = l2 ? tmp3382 : tmp3357;
  assign tmp4011 = l1 ? tmp4012 : tmp3989;
  assign tmp4010 = s0 ? tmp4011 : tmp3355;
  assign tmp4009 = s1 ? tmp3355 : tmp4010;
  assign tmp4008 = s2 ? tmp4009 : tmp3355;
  assign tmp4007 = s3 ? tmp3355 : tmp4008;
  assign tmp4014 = s1 ? tmp4010 : tmp3355;
  assign tmp4013 = s3 ? tmp3355 : tmp4014;
  assign tmp4006 = s4 ? tmp4007 : tmp4013;
  assign tmp4005 = s5 ? tmp3355 : tmp4006;
  assign tmp4004 = s6 ? tmp4005 : tmp3355;
  assign tmp4003 = s7 ? tmp3355 : tmp4004;
  assign tmp4018 = s4 ? tmp4007 : tmp3355;
  assign tmp4017 = s5 ? tmp3355 : tmp4018;
  assign tmp4016 = s6 ? tmp3355 : tmp4017;
  assign tmp4015 = s7 ? tmp3355 : tmp4016;
  assign tmp4002 = s8 ? tmp4003 : tmp4015;
  assign tmp4001 = s9 ? tmp3355 : tmp4002;
  assign tmp4022 = s6 ? tmp3355 : tmp4005;
  assign tmp4021 = s7 ? tmp3355 : tmp4022;
  assign tmp4020 = s8 ? tmp4003 : tmp4021;
  assign tmp4019 = s9 ? tmp3355 : tmp4020;
  assign tmp4000 = s10 ? tmp4001 : tmp4019;
  assign tmp3976 = s11 ? tmp3977 : tmp4000;
  assign tmp4035 = l1 ? tmp3886 : tmp3381;
  assign tmp4034 = s0 ? tmp4035 : tmp3632;
  assign tmp4033 = s1 ? tmp4034 : tmp3632;
  assign tmp4032 = s2 ? tmp3651 : tmp4033;
  assign tmp4036 = s2 ? tmp3632 : tmp4035;
  assign tmp4031 = s3 ? tmp4032 : tmp4036;
  assign tmp4030 = s4 ? tmp3679 : tmp4031;
  assign tmp4029 = s5 ? tmp3632 : tmp4030;
  assign tmp4028 = s6 ? tmp4029 : tmp3689;
  assign tmp4027 = s7 ? tmp3654 : tmp4028;
  assign tmp4041 = s3 ? tmp4032 : tmp3632;
  assign tmp4040 = s4 ? tmp3679 : tmp4041;
  assign tmp4039 = s5 ? tmp3632 : tmp4040;
  assign tmp4038 = s6 ? tmp3715 : tmp4039;
  assign tmp4037 = s7 ? tmp3703 : tmp4038;
  assign tmp4026 = s8 ? tmp4027 : tmp4037;
  assign tmp4025 = s9 ? tmp3631 : tmp4026;
  assign tmp4045 = s6 ? tmp3672 : tmp4029;
  assign tmp4044 = s7 ? tmp3720 : tmp4045;
  assign tmp4043 = s8 ? tmp4027 : tmp4044;
  assign tmp4042 = s9 ? tmp3631 : tmp4043;
  assign tmp4024 = s10 ? tmp4025 : tmp4042;
  assign tmp4023 = s11 ? tmp3526 : tmp4024;
  assign tmp3975 = s12 ? tmp3976 : tmp4023;
  assign tmp3871 = s13 ? tmp3872 : tmp3975;
  assign tmp3722 = s15 ? tmp3723 : tmp3871;
  assign tmp3351 = s16 ? tmp3352 : tmp3722;
  assign s10n = tmp3351;

  assign tmp4057 = ~(l3 ? 1 : 0);
  assign tmp4056 = l2 ? 1 : tmp4057;
  assign tmp4055 = l1 ? tmp4056 : 1;
  assign tmp4061 = l2 ? 1 : 0;
  assign tmp4060 = l1 ? tmp4061 : 1;
  assign tmp4059 = s0 ? tmp4060 : tmp4055;
  assign tmp4058 = s1 ? tmp4055 : tmp4059;
  assign tmp4054 = s2 ? tmp4055 : tmp4058;
  assign tmp4065 = s1 ? tmp4059 : 1;
  assign tmp4067 = s0 ? tmp4055 : 1;
  assign tmp4068 = s0 ? tmp4055 : tmp4061;
  assign tmp4066 = s1 ? tmp4067 : tmp4068;
  assign tmp4064 = s2 ? tmp4065 : tmp4066;
  assign tmp4071 = s0 ? tmp4061 : 1;
  assign tmp4070 = s1 ? tmp4061 : tmp4071;
  assign tmp4073 = s0 ? 1 : tmp4055;
  assign tmp4074 = s0 ? tmp4055 : tmp4060;
  assign tmp4072 = s1 ? tmp4073 : tmp4074;
  assign tmp4069 = s2 ? tmp4070 : tmp4072;
  assign tmp4063 = s3 ? tmp4064 : tmp4069;
  assign tmp4078 = s0 ? tmp4060 : 1;
  assign tmp4079 = s0 ? 1 : tmp4056;
  assign tmp4077 = s1 ? tmp4078 : tmp4079;
  assign tmp4081 = s0 ? tmp4056 : tmp4055;
  assign tmp4082 = s0 ? tmp4061 : tmp4056;
  assign tmp4080 = s1 ? tmp4081 : tmp4082;
  assign tmp4076 = s2 ? tmp4077 : tmp4080;
  assign tmp4085 = s0 ? tmp4061 : tmp4055;
  assign tmp4084 = s1 ? tmp4085 : tmp4055;
  assign tmp4083 = s2 ? tmp4084 : tmp4077;
  assign tmp4075 = s3 ? tmp4076 : tmp4083;
  assign tmp4062 = s4 ? tmp4063 : tmp4075;
  assign tmp4053 = s5 ? tmp4054 : tmp4062;
  assign tmp4052 = s6 ? tmp4053 : 1;
  assign tmp4051 = s7 ? tmp4052 : 1;
  assign tmp4050 = s8 ? tmp4051 : 1;
  assign tmp4049 = s9 ? 1 : tmp4050;
  assign tmp4092 = l1 ? 1 : tmp4056;
  assign tmp4095 = l1 ? 1 : tmp4061;
  assign tmp4094 = s0 ? tmp4092 : tmp4095;
  assign tmp4093 = s1 ? tmp4094 : tmp4092;
  assign tmp4091 = s2 ? tmp4092 : tmp4093;
  assign tmp4099 = s1 ? tmp4092 : tmp4061;
  assign tmp4101 = s0 ? tmp4092 : tmp4061;
  assign tmp4102 = s0 ? tmp4092 : 1;
  assign tmp4100 = s1 ? tmp4101 : tmp4102;
  assign tmp4098 = s2 ? tmp4099 : tmp4100;
  assign tmp4104 = s1 ? 1 : tmp4079;
  assign tmp4106 = s0 ? tmp4056 : tmp4095;
  assign tmp4107 = s0 ? tmp4095 : tmp4092;
  assign tmp4105 = s1 ? tmp4106 : tmp4107;
  assign tmp4103 = s2 ? tmp4104 : tmp4105;
  assign tmp4097 = s3 ? tmp4098 : tmp4103;
  assign tmp4110 = s1 ? tmp4102 : 1;
  assign tmp4111 = s1 ? tmp4092 : 1;
  assign tmp4109 = s2 ? tmp4110 : tmp4111;
  assign tmp4114 = s0 ? 1 : tmp4092;
  assign tmp4113 = s1 ? tmp4114 : tmp4107;
  assign tmp4116 = s0 ? tmp4056 : 1;
  assign tmp4115 = s1 ? tmp4102 : tmp4116;
  assign tmp4112 = s2 ? tmp4113 : tmp4115;
  assign tmp4108 = s3 ? tmp4109 : tmp4112;
  assign tmp4096 = s4 ? tmp4097 : tmp4108;
  assign tmp4090 = s5 ? tmp4091 : tmp4096;
  assign tmp4089 = s6 ? tmp4090 : 1;
  assign tmp4088 = s7 ? tmp4089 : 1;
  assign tmp4087 = s8 ? tmp4088 : 1;
  assign tmp4086 = s9 ? 1 : tmp4087;
  assign tmp4048 = s11 ? tmp4049 : tmp4086;
  assign tmp4124 = l1 ? tmp4056 : tmp4061;
  assign tmp4126 = s0 ? tmp4061 : tmp4124;
  assign tmp4125 = s1 ? tmp4124 : tmp4126;
  assign tmp4123 = s2 ? tmp4124 : tmp4125;
  assign tmp4130 = s1 ? tmp4126 : tmp4061;
  assign tmp4131 = s0 ? tmp4124 : tmp4061;
  assign tmp4129 = s2 ? tmp4130 : tmp4131;
  assign tmp4134 = s0 ? tmp4061 : tmp4095;
  assign tmp4133 = s1 ? tmp4061 : tmp4134;
  assign tmp4135 = s1 ? tmp4124 : tmp4131;
  assign tmp4132 = s2 ? tmp4133 : tmp4135;
  assign tmp4128 = s3 ? tmp4129 : tmp4132;
  assign tmp4138 = s1 ? tmp4061 : tmp4126;
  assign tmp4137 = s2 ? tmp4138 : tmp4125;
  assign tmp4140 = s1 ? tmp4126 : tmp4124;
  assign tmp4141 = s1 ? tmp4061 : tmp4124;
  assign tmp4139 = s2 ? tmp4140 : tmp4141;
  assign tmp4136 = s3 ? tmp4137 : tmp4139;
  assign tmp4127 = s4 ? tmp4128 : tmp4136;
  assign tmp4122 = s5 ? tmp4123 : tmp4127;
  assign tmp4121 = s6 ? tmp4122 : 1;
  assign tmp4120 = s7 ? tmp4121 : 1;
  assign tmp4119 = s8 ? tmp4120 : 1;
  assign tmp4118 = s9 ? 1 : tmp4119;
  assign tmp4148 = l1 ? tmp4061 : tmp4056;
  assign tmp4150 = s0 ? tmp4148 : tmp4061;
  assign tmp4149 = s1 ? tmp4150 : tmp4148;
  assign tmp4147 = s2 ? tmp4148 : tmp4149;
  assign tmp4154 = s1 ? tmp4148 : tmp4061;
  assign tmp4153 = s2 ? tmp4154 : tmp4150;
  assign tmp4157 = s0 ? tmp4061 : tmp4148;
  assign tmp4156 = s1 ? tmp4061 : tmp4157;
  assign tmp4158 = s1 ? tmp4150 : tmp4157;
  assign tmp4155 = s2 ? tmp4156 : tmp4158;
  assign tmp4152 = s3 ? tmp4153 : tmp4155;
  assign tmp4162 = s0 ? tmp4061 : tmp4060;
  assign tmp4161 = s1 ? tmp4148 : tmp4162;
  assign tmp4160 = s2 ? tmp4148 : tmp4161;
  assign tmp4163 = s2 ? tmp4157 : tmp4148;
  assign tmp4159 = s3 ? tmp4160 : tmp4163;
  assign tmp4151 = s4 ? tmp4152 : tmp4159;
  assign tmp4146 = s5 ? tmp4147 : tmp4151;
  assign tmp4145 = s6 ? tmp4146 : 1;
  assign tmp4144 = s7 ? tmp4145 : 1;
  assign tmp4143 = s8 ? tmp4144 : 1;
  assign tmp4142 = s9 ? 1 : tmp4143;
  assign tmp4117 = s11 ? tmp4118 : tmp4142;
  assign tmp4047 = s12 ? tmp4048 : tmp4117;
  assign tmp4174 = l3 ? 1 : 0;
  assign tmp4173 = l2 ? 1 : tmp4174;
  assign tmp4172 = l1 ? 1 : tmp4173;
  assign tmp4176 = s0 ? tmp4173 : tmp4172;
  assign tmp4175 = s1 ? tmp4172 : tmp4176;
  assign tmp4171 = s2 ? tmp4172 : tmp4175;
  assign tmp4180 = s1 ? tmp4176 : 1;
  assign tmp4181 = s0 ? tmp4172 : 1;
  assign tmp4179 = s2 ? tmp4180 : tmp4181;
  assign tmp4184 = s0 ? 1 : tmp4172;
  assign tmp4183 = s1 ? 1 : tmp4184;
  assign tmp4186 = s0 ? 1 : tmp4173;
  assign tmp4185 = s1 ? tmp4181 : tmp4186;
  assign tmp4182 = s2 ? tmp4183 : tmp4185;
  assign tmp4178 = s3 ? tmp4179 : tmp4182;
  assign tmp4190 = s0 ? tmp4173 : tmp4061;
  assign tmp4189 = s1 ? tmp4190 : tmp4134;
  assign tmp4192 = s0 ? tmp4095 : tmp4172;
  assign tmp4193 = s0 ? 1 : tmp4095;
  assign tmp4191 = s1 ? tmp4192 : tmp4193;
  assign tmp4188 = s2 ? tmp4189 : tmp4191;
  assign tmp4195 = s1 ? tmp4184 : tmp4172;
  assign tmp4197 = s0 ? tmp4172 : tmp4095;
  assign tmp4196 = s1 ? tmp4190 : tmp4197;
  assign tmp4194 = s2 ? tmp4195 : tmp4196;
  assign tmp4187 = s3 ? tmp4188 : tmp4194;
  assign tmp4177 = s4 ? tmp4178 : tmp4187;
  assign tmp4170 = s5 ? tmp4171 : tmp4177;
  assign tmp4169 = s6 ? tmp4170 : 1;
  assign tmp4168 = s7 ? tmp4169 : 1;
  assign tmp4167 = s8 ? tmp4168 : 1;
  assign tmp4166 = s9 ? 1 : tmp4167;
  assign tmp4165 = s11 ? tmp4166 : tmp4049;
  assign tmp4204 = l1 ? tmp4173 : tmp4061;
  assign tmp4208 = s1 ? tmp4204 : tmp4061;
  assign tmp4210 = s0 ? tmp4204 : tmp4061;
  assign tmp4209 = s1 ? tmp4210 : tmp4204;
  assign tmp4207 = s2 ? tmp4208 : tmp4209;
  assign tmp4213 = s0 ? 1 : tmp4061;
  assign tmp4212 = s1 ? 1 : tmp4213;
  assign tmp4215 = s0 ? tmp4061 : tmp4204;
  assign tmp4214 = s1 ? tmp4215 : tmp4204;
  assign tmp4211 = s2 ? tmp4212 : tmp4214;
  assign tmp4206 = s3 ? tmp4207 : tmp4211;
  assign tmp4219 = s0 ? tmp4095 : tmp4061;
  assign tmp4218 = s1 ? tmp4219 : tmp4215;
  assign tmp4217 = s2 ? tmp4218 : tmp4204;
  assign tmp4220 = s2 ? tmp4204 : tmp4218;
  assign tmp4216 = s3 ? tmp4217 : tmp4220;
  assign tmp4205 = s4 ? tmp4206 : tmp4216;
  assign tmp4203 = s5 ? tmp4204 : tmp4205;
  assign tmp4202 = s6 ? tmp4203 : 1;
  assign tmp4201 = s7 ? tmp4202 : 1;
  assign tmp4200 = s8 ? tmp4201 : 1;
  assign tmp4199 = s9 ? 1 : tmp4200;
  assign tmp4226 = l1 ? tmp4061 : tmp4173;
  assign tmp4231 = s0 ? tmp4226 : tmp4061;
  assign tmp4230 = s1 ? tmp4226 : tmp4231;
  assign tmp4229 = s2 ? tmp4226 : tmp4230;
  assign tmp4234 = s0 ? tmp4061 : tmp4226;
  assign tmp4233 = s1 ? tmp4061 : tmp4234;
  assign tmp4232 = s2 ? tmp4233 : tmp4226;
  assign tmp4228 = s3 ? tmp4229 : tmp4232;
  assign tmp4237 = s1 ? tmp4231 : tmp4061;
  assign tmp4238 = s1 ? tmp4234 : tmp4061;
  assign tmp4236 = s2 ? tmp4237 : tmp4238;
  assign tmp4240 = s1 ? tmp4234 : tmp4226;
  assign tmp4239 = s2 ? tmp4240 : tmp4231;
  assign tmp4235 = s3 ? tmp4236 : tmp4239;
  assign tmp4227 = s4 ? tmp4228 : tmp4235;
  assign tmp4225 = s5 ? tmp4226 : tmp4227;
  assign tmp4224 = s6 ? tmp4225 : 1;
  assign tmp4223 = s7 ? tmp4224 : 1;
  assign tmp4222 = s8 ? tmp4223 : 1;
  assign tmp4221 = s9 ? 1 : tmp4222;
  assign tmp4198 = s11 ? tmp4199 : tmp4221;
  assign tmp4164 = s12 ? tmp4165 : tmp4198;
  assign tmp4046 = ~(s13 ? tmp4047 : tmp4164);
  assign s9n = tmp4046;

  assign tmp4242 = l2 ? 1 : 0;
  assign tmp4245 = s6 ? 1 : 0;
  assign tmp4244 = s7 ? 1 : tmp4245;
  assign tmp4247 = s6 ? 1 : tmp4242;
  assign tmp4246 = ~(s7 ? tmp4247 : 0);
  assign tmp4243 = ~(s8 ? tmp4244 : tmp4246);
  assign tmp4241 = s9 ? tmp4242 : tmp4243;
  assign s8n = tmp4241;

  assign tmp4259 = ~(l3 ? 1 : 0);
  assign tmp4258 = l2 ? 1 : tmp4259;
  assign tmp4257 = l1 ? tmp4258 : 1;
  assign tmp4263 = l2 ? 1 : 0;
  assign tmp4262 = l1 ? tmp4263 : 1;
  assign tmp4261 = s0 ? tmp4262 : tmp4257;
  assign tmp4260 = s1 ? tmp4257 : tmp4261;
  assign tmp4256 = s2 ? tmp4257 : tmp4260;
  assign tmp4267 = s1 ? tmp4261 : 1;
  assign tmp4269 = s0 ? tmp4257 : 1;
  assign tmp4270 = s0 ? tmp4257 : tmp4263;
  assign tmp4268 = s1 ? tmp4269 : tmp4270;
  assign tmp4266 = s2 ? tmp4267 : tmp4268;
  assign tmp4273 = s0 ? tmp4263 : 1;
  assign tmp4272 = s1 ? tmp4263 : tmp4273;
  assign tmp4275 = s0 ? 1 : tmp4257;
  assign tmp4276 = s0 ? tmp4257 : tmp4262;
  assign tmp4274 = s1 ? tmp4275 : tmp4276;
  assign tmp4271 = s2 ? tmp4272 : tmp4274;
  assign tmp4265 = s3 ? tmp4266 : tmp4271;
  assign tmp4280 = s0 ? tmp4262 : 1;
  assign tmp4281 = s0 ? 1 : tmp4258;
  assign tmp4279 = s1 ? tmp4280 : tmp4281;
  assign tmp4283 = s0 ? tmp4258 : tmp4257;
  assign tmp4284 = s0 ? tmp4263 : tmp4258;
  assign tmp4282 = s1 ? tmp4283 : tmp4284;
  assign tmp4278 = s2 ? tmp4279 : tmp4282;
  assign tmp4287 = s0 ? tmp4263 : tmp4257;
  assign tmp4286 = s1 ? tmp4287 : tmp4257;
  assign tmp4285 = s2 ? tmp4286 : tmp4279;
  assign tmp4277 = s3 ? tmp4278 : tmp4285;
  assign tmp4264 = s4 ? tmp4265 : tmp4277;
  assign tmp4255 = s5 ? tmp4256 : tmp4264;
  assign tmp4254 = s6 ? tmp4255 : 1;
  assign tmp4289 = ~(l2 ? 1 : 0);
  assign tmp4288 = ~(s6 ? 1 : tmp4289);
  assign tmp4253 = s7 ? tmp4254 : tmp4288;
  assign tmp4291 = ~(s6 ? 1 : 0);
  assign tmp4290 = ~(s7 ? 1 : tmp4291);
  assign tmp4252 = ~(s8 ? tmp4253 : tmp4290);
  assign tmp4251 = s9 ? 1 : tmp4252;
  assign tmp4298 = l1 ? 1 : tmp4258;
  assign tmp4301 = l1 ? 1 : tmp4263;
  assign tmp4300 = s0 ? tmp4298 : tmp4301;
  assign tmp4299 = s1 ? tmp4300 : tmp4298;
  assign tmp4297 = s2 ? tmp4298 : tmp4299;
  assign tmp4305 = s1 ? tmp4298 : tmp4263;
  assign tmp4307 = s0 ? tmp4298 : tmp4263;
  assign tmp4308 = s0 ? tmp4298 : 1;
  assign tmp4306 = s1 ? tmp4307 : tmp4308;
  assign tmp4304 = s2 ? tmp4305 : tmp4306;
  assign tmp4310 = s1 ? 1 : tmp4281;
  assign tmp4312 = s0 ? tmp4258 : tmp4301;
  assign tmp4313 = s0 ? tmp4301 : tmp4298;
  assign tmp4311 = s1 ? tmp4312 : tmp4313;
  assign tmp4309 = s2 ? tmp4310 : tmp4311;
  assign tmp4303 = s3 ? tmp4304 : tmp4309;
  assign tmp4316 = s1 ? tmp4308 : 1;
  assign tmp4317 = s1 ? tmp4298 : 1;
  assign tmp4315 = s2 ? tmp4316 : tmp4317;
  assign tmp4320 = s0 ? 1 : tmp4298;
  assign tmp4319 = s1 ? tmp4320 : tmp4313;
  assign tmp4322 = s0 ? tmp4258 : 1;
  assign tmp4321 = s1 ? tmp4308 : tmp4322;
  assign tmp4318 = s2 ? tmp4319 : tmp4321;
  assign tmp4314 = s3 ? tmp4315 : tmp4318;
  assign tmp4302 = s4 ? tmp4303 : tmp4314;
  assign tmp4296 = s5 ? tmp4297 : tmp4302;
  assign tmp4295 = s6 ? tmp4296 : 1;
  assign tmp4294 = s7 ? tmp4295 : tmp4288;
  assign tmp4293 = ~(s8 ? tmp4294 : tmp4290);
  assign tmp4292 = s9 ? 1 : tmp4293;
  assign tmp4250 = s11 ? tmp4251 : tmp4292;
  assign tmp4330 = l1 ? tmp4258 : tmp4263;
  assign tmp4332 = s0 ? tmp4263 : tmp4330;
  assign tmp4331 = s1 ? tmp4330 : tmp4332;
  assign tmp4329 = s2 ? tmp4330 : tmp4331;
  assign tmp4336 = s1 ? tmp4332 : tmp4263;
  assign tmp4337 = s0 ? tmp4330 : tmp4263;
  assign tmp4335 = s2 ? tmp4336 : tmp4337;
  assign tmp4340 = s0 ? tmp4263 : tmp4301;
  assign tmp4339 = s1 ? tmp4263 : tmp4340;
  assign tmp4341 = s1 ? tmp4330 : tmp4337;
  assign tmp4338 = s2 ? tmp4339 : tmp4341;
  assign tmp4334 = s3 ? tmp4335 : tmp4338;
  assign tmp4344 = s1 ? tmp4263 : tmp4332;
  assign tmp4343 = s2 ? tmp4344 : tmp4331;
  assign tmp4346 = s1 ? tmp4332 : tmp4330;
  assign tmp4347 = s1 ? tmp4263 : tmp4330;
  assign tmp4345 = s2 ? tmp4346 : tmp4347;
  assign tmp4342 = s3 ? tmp4343 : tmp4345;
  assign tmp4333 = s4 ? tmp4334 : tmp4342;
  assign tmp4328 = s5 ? tmp4329 : tmp4333;
  assign tmp4327 = s6 ? tmp4328 : 1;
  assign tmp4326 = s7 ? tmp4327 : tmp4288;
  assign tmp4325 = ~(s8 ? tmp4326 : tmp4290);
  assign tmp4324 = s9 ? 1 : tmp4325;
  assign tmp4354 = l1 ? tmp4263 : tmp4258;
  assign tmp4356 = s0 ? tmp4354 : tmp4263;
  assign tmp4355 = s1 ? tmp4356 : tmp4354;
  assign tmp4353 = s2 ? tmp4354 : tmp4355;
  assign tmp4360 = s1 ? tmp4354 : tmp4263;
  assign tmp4359 = s2 ? tmp4360 : tmp4356;
  assign tmp4363 = s0 ? tmp4263 : tmp4354;
  assign tmp4362 = s1 ? tmp4263 : tmp4363;
  assign tmp4364 = s1 ? tmp4356 : tmp4363;
  assign tmp4361 = s2 ? tmp4362 : tmp4364;
  assign tmp4358 = s3 ? tmp4359 : tmp4361;
  assign tmp4368 = s0 ? tmp4263 : tmp4262;
  assign tmp4367 = s1 ? tmp4354 : tmp4368;
  assign tmp4366 = s2 ? tmp4354 : tmp4367;
  assign tmp4369 = s2 ? tmp4363 : tmp4354;
  assign tmp4365 = s3 ? tmp4366 : tmp4369;
  assign tmp4357 = s4 ? tmp4358 : tmp4365;
  assign tmp4352 = s5 ? tmp4353 : tmp4357;
  assign tmp4351 = s6 ? tmp4352 : 1;
  assign tmp4350 = s7 ? tmp4351 : tmp4288;
  assign tmp4349 = ~(s8 ? tmp4350 : tmp4290);
  assign tmp4348 = s9 ? 1 : tmp4349;
  assign tmp4323 = s11 ? tmp4324 : tmp4348;
  assign tmp4249 = s12 ? tmp4250 : tmp4323;
  assign tmp4380 = l3 ? 1 : 0;
  assign tmp4379 = l2 ? 1 : tmp4380;
  assign tmp4378 = l1 ? 1 : tmp4379;
  assign tmp4382 = s0 ? tmp4379 : tmp4378;
  assign tmp4381 = s1 ? tmp4378 : tmp4382;
  assign tmp4377 = s2 ? tmp4378 : tmp4381;
  assign tmp4386 = s1 ? tmp4382 : 1;
  assign tmp4387 = s0 ? tmp4378 : 1;
  assign tmp4385 = s2 ? tmp4386 : tmp4387;
  assign tmp4390 = s0 ? 1 : tmp4378;
  assign tmp4389 = s1 ? 1 : tmp4390;
  assign tmp4392 = s0 ? 1 : tmp4379;
  assign tmp4391 = s1 ? tmp4387 : tmp4392;
  assign tmp4388 = s2 ? tmp4389 : tmp4391;
  assign tmp4384 = s3 ? tmp4385 : tmp4388;
  assign tmp4396 = s0 ? tmp4379 : tmp4263;
  assign tmp4395 = s1 ? tmp4396 : tmp4340;
  assign tmp4398 = s0 ? tmp4301 : tmp4378;
  assign tmp4399 = s0 ? 1 : tmp4301;
  assign tmp4397 = s1 ? tmp4398 : tmp4399;
  assign tmp4394 = s2 ? tmp4395 : tmp4397;
  assign tmp4401 = s1 ? tmp4390 : tmp4378;
  assign tmp4403 = s0 ? tmp4378 : tmp4301;
  assign tmp4402 = s1 ? tmp4396 : tmp4403;
  assign tmp4400 = s2 ? tmp4401 : tmp4402;
  assign tmp4393 = s3 ? tmp4394 : tmp4400;
  assign tmp4383 = s4 ? tmp4384 : tmp4393;
  assign tmp4376 = s5 ? tmp4377 : tmp4383;
  assign tmp4375 = s6 ? tmp4376 : 1;
  assign tmp4374 = s7 ? tmp4375 : tmp4288;
  assign tmp4373 = ~(s8 ? tmp4374 : tmp4290);
  assign tmp4372 = s9 ? 1 : tmp4373;
  assign tmp4371 = s11 ? tmp4372 : tmp4251;
  assign tmp4410 = l1 ? tmp4379 : tmp4263;
  assign tmp4414 = s1 ? tmp4410 : tmp4263;
  assign tmp4416 = s0 ? tmp4410 : tmp4263;
  assign tmp4415 = s1 ? tmp4416 : tmp4410;
  assign tmp4413 = s2 ? tmp4414 : tmp4415;
  assign tmp4419 = s0 ? 1 : tmp4263;
  assign tmp4418 = s1 ? 1 : tmp4419;
  assign tmp4421 = s0 ? tmp4263 : tmp4410;
  assign tmp4420 = s1 ? tmp4421 : tmp4410;
  assign tmp4417 = s2 ? tmp4418 : tmp4420;
  assign tmp4412 = s3 ? tmp4413 : tmp4417;
  assign tmp4425 = s0 ? tmp4301 : tmp4263;
  assign tmp4424 = s1 ? tmp4425 : tmp4421;
  assign tmp4423 = s2 ? tmp4424 : tmp4410;
  assign tmp4426 = s2 ? tmp4410 : tmp4424;
  assign tmp4422 = s3 ? tmp4423 : tmp4426;
  assign tmp4411 = s4 ? tmp4412 : tmp4422;
  assign tmp4409 = s5 ? tmp4410 : tmp4411;
  assign tmp4408 = s6 ? tmp4409 : 1;
  assign tmp4407 = s7 ? tmp4408 : tmp4288;
  assign tmp4406 = ~(s8 ? tmp4407 : tmp4290);
  assign tmp4405 = s9 ? 1 : tmp4406;
  assign tmp4432 = l1 ? tmp4263 : tmp4379;
  assign tmp4437 = s0 ? tmp4432 : tmp4263;
  assign tmp4436 = s1 ? tmp4432 : tmp4437;
  assign tmp4435 = s2 ? tmp4432 : tmp4436;
  assign tmp4440 = s0 ? tmp4263 : tmp4432;
  assign tmp4439 = s1 ? tmp4263 : tmp4440;
  assign tmp4438 = s2 ? tmp4439 : tmp4432;
  assign tmp4434 = s3 ? tmp4435 : tmp4438;
  assign tmp4443 = s1 ? tmp4437 : tmp4263;
  assign tmp4444 = s1 ? tmp4440 : tmp4263;
  assign tmp4442 = s2 ? tmp4443 : tmp4444;
  assign tmp4446 = s1 ? tmp4440 : tmp4432;
  assign tmp4445 = s2 ? tmp4446 : tmp4437;
  assign tmp4441 = s3 ? tmp4442 : tmp4445;
  assign tmp4433 = s4 ? tmp4434 : tmp4441;
  assign tmp4431 = s5 ? tmp4432 : tmp4433;
  assign tmp4430 = s6 ? tmp4431 : 1;
  assign tmp4429 = s7 ? tmp4430 : tmp4288;
  assign tmp4428 = ~(s8 ? tmp4429 : tmp4290);
  assign tmp4427 = s9 ? 1 : tmp4428;
  assign tmp4404 = s11 ? tmp4405 : tmp4427;
  assign tmp4370 = s12 ? tmp4371 : tmp4404;
  assign tmp4248 = ~(s13 ? tmp4249 : tmp4370);
  assign s7n = tmp4248;

  assign tmp4459 = ~(l3 ? 1 : 0);
  assign tmp4458 = l2 ? 1 : tmp4459;
  assign tmp4457 = l1 ? tmp4458 : 1;
  assign tmp4463 = l2 ? 1 : 0;
  assign tmp4462 = l1 ? tmp4463 : 1;
  assign tmp4461 = s0 ? tmp4462 : tmp4457;
  assign tmp4460 = s1 ? tmp4457 : tmp4461;
  assign tmp4456 = s2 ? tmp4457 : tmp4460;
  assign tmp4467 = s1 ? tmp4461 : 1;
  assign tmp4469 = s0 ? tmp4457 : 1;
  assign tmp4470 = s0 ? tmp4457 : tmp4463;
  assign tmp4468 = s1 ? tmp4469 : tmp4470;
  assign tmp4466 = s2 ? tmp4467 : tmp4468;
  assign tmp4473 = s0 ? tmp4463 : 1;
  assign tmp4472 = s1 ? tmp4463 : tmp4473;
  assign tmp4475 = s0 ? 1 : tmp4457;
  assign tmp4476 = s0 ? tmp4457 : tmp4462;
  assign tmp4474 = s1 ? tmp4475 : tmp4476;
  assign tmp4471 = s2 ? tmp4472 : tmp4474;
  assign tmp4465 = s3 ? tmp4466 : tmp4471;
  assign tmp4480 = s0 ? tmp4462 : 1;
  assign tmp4481 = s0 ? 1 : tmp4458;
  assign tmp4479 = s1 ? tmp4480 : tmp4481;
  assign tmp4483 = s0 ? tmp4458 : tmp4457;
  assign tmp4484 = s0 ? tmp4463 : tmp4458;
  assign tmp4482 = s1 ? tmp4483 : tmp4484;
  assign tmp4478 = s2 ? tmp4479 : tmp4482;
  assign tmp4487 = s0 ? tmp4463 : tmp4457;
  assign tmp4486 = s1 ? tmp4487 : tmp4457;
  assign tmp4485 = s2 ? tmp4486 : tmp4479;
  assign tmp4477 = s3 ? tmp4478 : tmp4485;
  assign tmp4464 = s4 ? tmp4465 : tmp4477;
  assign tmp4455 = s5 ? tmp4456 : tmp4464;
  assign tmp4454 = s6 ? tmp4455 : tmp4463;
  assign tmp4493 = s1 ? tmp4461 : tmp4462;
  assign tmp4494 = s1 ? tmp4476 : tmp4470;
  assign tmp4492 = s2 ? tmp4493 : tmp4494;
  assign tmp4498 = ~(l2 ? 1 : 0);
  assign tmp4497 = s0 ? tmp4463 : tmp4498;
  assign tmp4496 = s1 ? tmp4463 : tmp4497;
  assign tmp4503 = l3 ? 1 : 0;
  assign tmp4502 = l2 ? tmp4503 : tmp4459;
  assign tmp4501 = ~(l1 ? tmp4502 : 1);
  assign tmp4500 = s0 ? tmp4463 : tmp4501;
  assign tmp4505 = l1 ? tmp4502 : 1;
  assign tmp4504 = ~(s0 ? tmp4505 : tmp4462);
  assign tmp4499 = ~(s1 ? tmp4500 : tmp4504);
  assign tmp4495 = s2 ? tmp4496 : tmp4499;
  assign tmp4491 = s3 ? tmp4492 : tmp4495;
  assign tmp4509 = s0 ? tmp4462 : tmp4458;
  assign tmp4508 = s1 ? tmp4462 : tmp4509;
  assign tmp4507 = s2 ? tmp4508 : tmp4482;
  assign tmp4512 = s0 ? tmp4505 : tmp4457;
  assign tmp4511 = s1 ? tmp4487 : tmp4512;
  assign tmp4515 = ~(l2 ? 1 : tmp4459);
  assign tmp4514 = ~(s0 ? tmp4463 : tmp4515);
  assign tmp4513 = s1 ? tmp4462 : tmp4514;
  assign tmp4510 = s2 ? tmp4511 : tmp4513;
  assign tmp4506 = s3 ? tmp4507 : tmp4510;
  assign tmp4490 = s4 ? tmp4491 : tmp4506;
  assign tmp4489 = ~(s5 ? tmp4456 : tmp4490);
  assign tmp4488 = s6 ? tmp4463 : tmp4489;
  assign tmp4453 = s7 ? tmp4454 : tmp4488;
  assign tmp4517 = s6 ? tmp4455 : 1;
  assign tmp4516 = ~(s7 ? tmp4517 : tmp4498);
  assign tmp4452 = ~(s8 ? tmp4453 : tmp4516);
  assign tmp4451 = s9 ? 1 : tmp4452;
  assign tmp4524 = l1 ? 1 : tmp4458;
  assign tmp4527 = l1 ? 1 : tmp4463;
  assign tmp4526 = s0 ? tmp4524 : tmp4527;
  assign tmp4525 = s1 ? tmp4526 : tmp4524;
  assign tmp4523 = s2 ? tmp4524 : tmp4525;
  assign tmp4531 = s1 ? tmp4524 : tmp4463;
  assign tmp4533 = s0 ? tmp4524 : tmp4463;
  assign tmp4534 = s0 ? tmp4524 : 1;
  assign tmp4532 = s1 ? tmp4533 : tmp4534;
  assign tmp4530 = s2 ? tmp4531 : tmp4532;
  assign tmp4536 = s1 ? 1 : tmp4481;
  assign tmp4538 = s0 ? tmp4458 : tmp4527;
  assign tmp4539 = s0 ? tmp4527 : tmp4524;
  assign tmp4537 = s1 ? tmp4538 : tmp4539;
  assign tmp4535 = s2 ? tmp4536 : tmp4537;
  assign tmp4529 = s3 ? tmp4530 : tmp4535;
  assign tmp4542 = s1 ? tmp4534 : 1;
  assign tmp4543 = s1 ? tmp4524 : 1;
  assign tmp4541 = s2 ? tmp4542 : tmp4543;
  assign tmp4546 = s0 ? 1 : tmp4524;
  assign tmp4545 = s1 ? tmp4546 : tmp4539;
  assign tmp4548 = s0 ? tmp4458 : 1;
  assign tmp4547 = s1 ? tmp4534 : tmp4548;
  assign tmp4544 = s2 ? tmp4545 : tmp4547;
  assign tmp4540 = s3 ? tmp4541 : tmp4544;
  assign tmp4528 = s4 ? tmp4529 : tmp4540;
  assign tmp4522 = s5 ? tmp4523 : tmp4528;
  assign tmp4521 = s6 ? tmp4522 : tmp4463;
  assign tmp4554 = l2 ? tmp4503 : 1;
  assign tmp4553 = l1 ? tmp4554 : tmp4458;
  assign tmp4552 = s1 ? tmp4524 : tmp4553;
  assign tmp4556 = s0 ? tmp4553 : tmp4527;
  assign tmp4557 = s0 ? tmp4524 : tmp4553;
  assign tmp4555 = s1 ? tmp4556 : tmp4557;
  assign tmp4551 = s2 ? tmp4552 : tmp4555;
  assign tmp4561 = s1 ? tmp4553 : tmp4463;
  assign tmp4562 = s1 ? tmp4533 : tmp4556;
  assign tmp4560 = s2 ? tmp4561 : tmp4562;
  assign tmp4566 = ~(l1 ? tmp4463 : tmp4498);
  assign tmp4565 = s0 ? tmp4527 : tmp4566;
  assign tmp4568 = l1 ? tmp4463 : tmp4498;
  assign tmp4569 = ~(l2 ? tmp4503 : tmp4459);
  assign tmp4567 = ~(s0 ? tmp4568 : tmp4569);
  assign tmp4564 = s1 ? tmp4565 : tmp4567;
  assign tmp4571 = s0 ? tmp4502 : tmp4566;
  assign tmp4573 = ~(l1 ? 1 : tmp4458);
  assign tmp4572 = ~(s0 ? tmp4568 : tmp4573);
  assign tmp4570 = s1 ? tmp4571 : tmp4572;
  assign tmp4563 = s2 ? tmp4564 : tmp4570;
  assign tmp4559 = s3 ? tmp4560 : tmp4563;
  assign tmp4578 = ~(l1 ? tmp4463 : 0);
  assign tmp4577 = s0 ? tmp4524 : tmp4578;
  assign tmp4580 = l1 ? tmp4463 : 0;
  assign tmp4579 = ~(s0 ? tmp4580 : tmp4463);
  assign tmp4576 = s1 ? tmp4577 : tmp4579;
  assign tmp4582 = s0 ? tmp4527 : tmp4578;
  assign tmp4581 = s1 ? tmp4553 : tmp4582;
  assign tmp4575 = s2 ? tmp4576 : tmp4581;
  assign tmp4586 = l1 ? tmp4463 : tmp4515;
  assign tmp4585 = s0 ? tmp4568 : tmp4586;
  assign tmp4588 = ~(l1 ? tmp4554 : tmp4458);
  assign tmp4587 = s0 ? tmp4568 : tmp4588;
  assign tmp4584 = s1 ? tmp4585 : tmp4587;
  assign tmp4590 = s0 ? tmp4502 : tmp4498;
  assign tmp4589 = ~(s1 ? tmp4577 : tmp4590);
  assign tmp4583 = ~(s2 ? tmp4584 : tmp4589);
  assign tmp4574 = s3 ? tmp4575 : tmp4583;
  assign tmp4558 = s4 ? tmp4559 : tmp4574;
  assign tmp4550 = ~(s5 ? tmp4551 : tmp4558);
  assign tmp4549 = s6 ? tmp4463 : tmp4550;
  assign tmp4520 = s7 ? tmp4521 : tmp4549;
  assign tmp4592 = s6 ? tmp4522 : 1;
  assign tmp4591 = ~(s7 ? tmp4592 : tmp4498);
  assign tmp4519 = ~(s8 ? tmp4520 : tmp4591);
  assign tmp4518 = s9 ? 1 : tmp4519;
  assign tmp4450 = s11 ? tmp4451 : tmp4518;
  assign tmp4600 = l1 ? tmp4458 : tmp4463;
  assign tmp4602 = s0 ? tmp4463 : tmp4600;
  assign tmp4601 = s1 ? tmp4600 : tmp4602;
  assign tmp4599 = s2 ? tmp4600 : tmp4601;
  assign tmp4606 = s1 ? tmp4602 : tmp4463;
  assign tmp4607 = s0 ? tmp4600 : tmp4463;
  assign tmp4605 = s2 ? tmp4606 : tmp4607;
  assign tmp4610 = s0 ? tmp4463 : tmp4527;
  assign tmp4609 = s1 ? tmp4463 : tmp4610;
  assign tmp4611 = s1 ? tmp4600 : tmp4607;
  assign tmp4608 = s2 ? tmp4609 : tmp4611;
  assign tmp4604 = s3 ? tmp4605 : tmp4608;
  assign tmp4614 = s1 ? tmp4463 : tmp4602;
  assign tmp4613 = s2 ? tmp4614 : tmp4601;
  assign tmp4616 = s1 ? tmp4602 : tmp4600;
  assign tmp4617 = s1 ? tmp4463 : tmp4600;
  assign tmp4615 = s2 ? tmp4616 : tmp4617;
  assign tmp4612 = s3 ? tmp4613 : tmp4615;
  assign tmp4603 = s4 ? tmp4604 : tmp4612;
  assign tmp4598 = s5 ? tmp4599 : tmp4603;
  assign tmp4597 = s6 ? tmp4598 : tmp4463;
  assign tmp4624 = s0 ? tmp4463 : tmp4566;
  assign tmp4623 = s1 ? tmp4463 : tmp4624;
  assign tmp4626 = l1 ? tmp4502 : tmp4463;
  assign tmp4627 = s0 ? tmp4626 : tmp4463;
  assign tmp4625 = s1 ? tmp4626 : tmp4627;
  assign tmp4622 = s2 ? tmp4623 : tmp4625;
  assign tmp4621 = s3 ? tmp4605 : tmp4622;
  assign tmp4620 = s4 ? tmp4621 : tmp4612;
  assign tmp4619 = ~(s5 ? tmp4599 : tmp4620);
  assign tmp4618 = s6 ? tmp4463 : tmp4619;
  assign tmp4596 = s7 ? tmp4597 : tmp4618;
  assign tmp4629 = s6 ? tmp4598 : 1;
  assign tmp4628 = ~(s7 ? tmp4629 : tmp4498);
  assign tmp4595 = ~(s8 ? tmp4596 : tmp4628);
  assign tmp4594 = s9 ? 1 : tmp4595;
  assign tmp4636 = l1 ? tmp4463 : tmp4458;
  assign tmp4638 = s0 ? tmp4636 : tmp4463;
  assign tmp4637 = s1 ? tmp4638 : tmp4636;
  assign tmp4635 = s2 ? tmp4636 : tmp4637;
  assign tmp4642 = s1 ? tmp4636 : tmp4463;
  assign tmp4641 = s2 ? tmp4642 : tmp4638;
  assign tmp4645 = s0 ? tmp4463 : tmp4636;
  assign tmp4644 = s1 ? tmp4463 : tmp4645;
  assign tmp4646 = s1 ? tmp4638 : tmp4645;
  assign tmp4643 = s2 ? tmp4644 : tmp4646;
  assign tmp4640 = s3 ? tmp4641 : tmp4643;
  assign tmp4650 = s0 ? tmp4463 : tmp4462;
  assign tmp4649 = s1 ? tmp4636 : tmp4650;
  assign tmp4648 = s2 ? tmp4636 : tmp4649;
  assign tmp4651 = s2 ? tmp4645 : tmp4636;
  assign tmp4647 = s3 ? tmp4648 : tmp4651;
  assign tmp4639 = s4 ? tmp4640 : tmp4647;
  assign tmp4634 = s5 ? tmp4635 : tmp4639;
  assign tmp4633 = s6 ? tmp4634 : tmp4463;
  assign tmp4659 = l1 ? tmp4463 : tmp4502;
  assign tmp4658 = s0 ? tmp4463 : tmp4659;
  assign tmp4657 = s1 ? tmp4463 : tmp4658;
  assign tmp4661 = s0 ? tmp4659 : tmp4463;
  assign tmp4660 = s1 ? tmp4661 : tmp4645;
  assign tmp4656 = s2 ? tmp4657 : tmp4660;
  assign tmp4655 = s3 ? tmp4641 : tmp4656;
  assign tmp4654 = s4 ? tmp4655 : tmp4647;
  assign tmp4653 = ~(s5 ? tmp4635 : tmp4654);
  assign tmp4652 = s6 ? tmp4463 : tmp4653;
  assign tmp4632 = s7 ? tmp4633 : tmp4652;
  assign tmp4663 = s6 ? tmp4634 : 1;
  assign tmp4662 = ~(s7 ? tmp4663 : tmp4498);
  assign tmp4631 = ~(s8 ? tmp4632 : tmp4662);
  assign tmp4630 = s9 ? 1 : tmp4631;
  assign tmp4593 = s11 ? tmp4594 : tmp4630;
  assign tmp4449 = s12 ? tmp4450 : tmp4593;
  assign tmp4673 = l2 ? 1 : tmp4503;
  assign tmp4672 = l1 ? 1 : tmp4673;
  assign tmp4675 = s0 ? tmp4673 : tmp4672;
  assign tmp4674 = s1 ? tmp4672 : tmp4675;
  assign tmp4671 = s2 ? tmp4672 : tmp4674;
  assign tmp4679 = s1 ? tmp4675 : 1;
  assign tmp4680 = s0 ? tmp4672 : 1;
  assign tmp4678 = s2 ? tmp4679 : tmp4680;
  assign tmp4683 = s0 ? 1 : tmp4672;
  assign tmp4682 = s1 ? 1 : tmp4683;
  assign tmp4685 = s0 ? 1 : tmp4673;
  assign tmp4684 = s1 ? tmp4680 : tmp4685;
  assign tmp4681 = s2 ? tmp4682 : tmp4684;
  assign tmp4677 = s3 ? tmp4678 : tmp4681;
  assign tmp4689 = s0 ? tmp4673 : tmp4463;
  assign tmp4688 = s1 ? tmp4689 : tmp4610;
  assign tmp4691 = s0 ? tmp4527 : tmp4672;
  assign tmp4692 = s0 ? 1 : tmp4527;
  assign tmp4690 = s1 ? tmp4691 : tmp4692;
  assign tmp4687 = s2 ? tmp4688 : tmp4690;
  assign tmp4694 = s1 ? tmp4683 : tmp4672;
  assign tmp4696 = s0 ? tmp4672 : tmp4527;
  assign tmp4695 = s1 ? tmp4689 : tmp4696;
  assign tmp4693 = s2 ? tmp4694 : tmp4695;
  assign tmp4686 = s3 ? tmp4687 : tmp4693;
  assign tmp4676 = s4 ? tmp4677 : tmp4686;
  assign tmp4670 = s5 ? tmp4671 : tmp4676;
  assign tmp4669 = s6 ? tmp4670 : tmp4463;
  assign tmp4700 = l1 ? 1 : tmp4569;
  assign tmp4702 = s0 ? tmp4700 : tmp4672;
  assign tmp4701 = s1 ? tmp4700 : tmp4702;
  assign tmp4699 = s2 ? tmp4700 : tmp4701;
  assign tmp4707 = s0 ? tmp4673 : tmp4700;
  assign tmp4706 = s1 ? tmp4707 : tmp4568;
  assign tmp4709 = s0 ? tmp4700 : tmp4568;
  assign tmp4711 = l1 ? 1 : tmp4498;
  assign tmp4710 = s0 ? tmp4700 : tmp4711;
  assign tmp4708 = s1 ? tmp4709 : tmp4710;
  assign tmp4705 = s2 ? tmp4706 : tmp4708;
  assign tmp4714 = s0 ? tmp4711 : tmp4527;
  assign tmp4716 = ~(l1 ? tmp4463 : tmp4502);
  assign tmp4715 = s0 ? tmp4527 : tmp4716;
  assign tmp4713 = s1 ? tmp4714 : tmp4715;
  assign tmp4719 = ~(l2 ? 1 : tmp4503);
  assign tmp4718 = s0 ? tmp4463 : tmp4719;
  assign tmp4717 = ~(s1 ? tmp4661 : tmp4718);
  assign tmp4712 = s2 ? tmp4713 : tmp4717;
  assign tmp4704 = s3 ? tmp4705 : tmp4712;
  assign tmp4723 = s0 ? tmp4527 : tmp4700;
  assign tmp4722 = s1 ? tmp4723 : tmp4714;
  assign tmp4721 = s2 ? tmp4688 : tmp4722;
  assign tmp4727 = ~(l1 ? 1 : tmp4673);
  assign tmp4726 = ~(s0 ? tmp4463 : tmp4727);
  assign tmp4725 = s1 ? tmp4723 : tmp4726;
  assign tmp4730 = ~(l1 ? 1 : tmp4463);
  assign tmp4729 = ~(s0 ? tmp4659 : tmp4730);
  assign tmp4728 = s1 ? tmp4689 : tmp4729;
  assign tmp4724 = s2 ? tmp4725 : tmp4728;
  assign tmp4720 = s3 ? tmp4721 : tmp4724;
  assign tmp4703 = s4 ? tmp4704 : tmp4720;
  assign tmp4698 = ~(s5 ? tmp4699 : tmp4703);
  assign tmp4697 = s6 ? tmp4463 : tmp4698;
  assign tmp4668 = s7 ? tmp4669 : tmp4697;
  assign tmp4732 = s6 ? tmp4670 : 1;
  assign tmp4731 = ~(s7 ? tmp4732 : tmp4498);
  assign tmp4667 = ~(s8 ? tmp4668 : tmp4731);
  assign tmp4666 = s9 ? 1 : tmp4667;
  assign tmp4665 = s11 ? tmp4666 : tmp4451;
  assign tmp4739 = l1 ? tmp4673 : tmp4463;
  assign tmp4743 = s1 ? tmp4739 : tmp4463;
  assign tmp4745 = s0 ? tmp4739 : tmp4463;
  assign tmp4744 = s1 ? tmp4745 : tmp4739;
  assign tmp4742 = s2 ? tmp4743 : tmp4744;
  assign tmp4748 = s0 ? 1 : tmp4463;
  assign tmp4747 = s1 ? 1 : tmp4748;
  assign tmp4750 = s0 ? tmp4463 : tmp4739;
  assign tmp4749 = s1 ? tmp4750 : tmp4739;
  assign tmp4746 = s2 ? tmp4747 : tmp4749;
  assign tmp4741 = s3 ? tmp4742 : tmp4746;
  assign tmp4754 = s0 ? tmp4527 : tmp4463;
  assign tmp4753 = s1 ? tmp4754 : tmp4750;
  assign tmp4752 = s2 ? tmp4753 : tmp4739;
  assign tmp4755 = s2 ? tmp4739 : tmp4753;
  assign tmp4751 = s3 ? tmp4752 : tmp4755;
  assign tmp4740 = s4 ? tmp4741 : tmp4751;
  assign tmp4738 = s5 ? tmp4739 : tmp4740;
  assign tmp4737 = s6 ? tmp4738 : tmp4463;
  assign tmp4761 = s1 ? tmp4527 : tmp4754;
  assign tmp4764 = ~(l1 ? tmp4502 : tmp4498);
  assign tmp4763 = s0 ? tmp4463 : tmp4764;
  assign tmp4762 = s1 ? tmp4763 : tmp4739;
  assign tmp4760 = s2 ? tmp4761 : tmp4762;
  assign tmp4759 = s3 ? tmp4742 : tmp4760;
  assign tmp4758 = s4 ? tmp4759 : tmp4751;
  assign tmp4757 = ~(s5 ? tmp4739 : tmp4758);
  assign tmp4756 = s6 ? tmp4463 : tmp4757;
  assign tmp4736 = s7 ? tmp4737 : tmp4756;
  assign tmp4766 = s6 ? tmp4738 : 1;
  assign tmp4765 = ~(s7 ? tmp4766 : tmp4498);
  assign tmp4735 = ~(s8 ? tmp4736 : tmp4765);
  assign tmp4734 = s9 ? 1 : tmp4735;
  assign tmp4772 = l1 ? tmp4463 : tmp4673;
  assign tmp4777 = s0 ? tmp4772 : tmp4463;
  assign tmp4776 = s1 ? tmp4772 : tmp4777;
  assign tmp4775 = s2 ? tmp4772 : tmp4776;
  assign tmp4780 = s0 ? tmp4463 : tmp4772;
  assign tmp4779 = s1 ? tmp4463 : tmp4780;
  assign tmp4778 = s2 ? tmp4779 : tmp4772;
  assign tmp4774 = s3 ? tmp4775 : tmp4778;
  assign tmp4783 = s1 ? tmp4777 : tmp4463;
  assign tmp4784 = s1 ? tmp4780 : tmp4463;
  assign tmp4782 = s2 ? tmp4783 : tmp4784;
  assign tmp4786 = s1 ? tmp4780 : tmp4772;
  assign tmp4785 = s2 ? tmp4786 : tmp4777;
  assign tmp4781 = s3 ? tmp4782 : tmp4785;
  assign tmp4773 = s4 ? tmp4774 : tmp4781;
  assign tmp4771 = s5 ? tmp4772 : tmp4773;
  assign tmp4770 = s6 ? tmp4771 : tmp4463;
  assign tmp4794 = l1 ? tmp4463 : tmp4569;
  assign tmp4793 = s0 ? tmp4463 : tmp4794;
  assign tmp4792 = s1 ? tmp4463 : tmp4793;
  assign tmp4791 = s2 ? tmp4792 : tmp4772;
  assign tmp4790 = s3 ? tmp4775 : tmp4791;
  assign tmp4789 = s4 ? tmp4790 : tmp4781;
  assign tmp4788 = ~(s5 ? tmp4772 : tmp4789);
  assign tmp4787 = s6 ? tmp4463 : tmp4788;
  assign tmp4769 = s7 ? tmp4770 : tmp4787;
  assign tmp4796 = s6 ? tmp4771 : 1;
  assign tmp4795 = ~(s7 ? tmp4796 : tmp4498);
  assign tmp4768 = ~(s8 ? tmp4769 : tmp4795);
  assign tmp4767 = s9 ? 1 : tmp4768;
  assign tmp4733 = s11 ? tmp4734 : tmp4767;
  assign tmp4664 = s12 ? tmp4665 : tmp4733;
  assign tmp4448 = s13 ? tmp4449 : tmp4664;
  assign tmp4809 = s1 ? 1 : tmp4462;
  assign tmp4811 = s0 ? 1 : tmp4462;
  assign tmp4810 = s1 ? tmp4811 : tmp4692;
  assign tmp4808 = s2 ? tmp4809 : tmp4810;
  assign tmp4814 = s0 ? tmp4527 : tmp4498;
  assign tmp4813 = s1 ? tmp4527 : tmp4814;
  assign tmp4816 = s0 ? tmp4463 : tmp4580;
  assign tmp4817 = s0 ? tmp4580 : 0;
  assign tmp4815 = ~(s1 ? tmp4816 : tmp4817);
  assign tmp4812 = s2 ? tmp4813 : tmp4815;
  assign tmp4807 = s3 ? tmp4808 : tmp4812;
  assign tmp4821 = s0 ? tmp4462 : tmp4711;
  assign tmp4820 = s1 ? tmp4811 : tmp4821;
  assign tmp4823 = s0 ? tmp4711 : 1;
  assign tmp4824 = s0 ? tmp4527 : 1;
  assign tmp4822 = s1 ? tmp4823 : tmp4824;
  assign tmp4819 = s2 ? tmp4820 : tmp4822;
  assign tmp4827 = ~(s0 ? tmp4580 : 0);
  assign tmp4826 = s1 ? tmp4824 : tmp4827;
  assign tmp4830 = ~(l1 ? 1 : tmp4498);
  assign tmp4829 = ~(s0 ? tmp4463 : tmp4830);
  assign tmp4828 = s1 ? tmp4811 : tmp4829;
  assign tmp4825 = s2 ? tmp4826 : tmp4828;
  assign tmp4818 = s3 ? tmp4819 : tmp4825;
  assign tmp4806 = s4 ? tmp4807 : tmp4818;
  assign tmp4805 = ~(s5 ? 1 : tmp4806);
  assign tmp4804 = s6 ? tmp4463 : tmp4805;
  assign tmp4803 = s7 ? tmp4454 : tmp4804;
  assign tmp4831 = ~(s7 ? 1 : tmp4498);
  assign tmp4802 = ~(s8 ? tmp4803 : tmp4831);
  assign tmp4801 = s9 ? 1 : tmp4802;
  assign tmp4839 = l1 ? tmp4554 : 1;
  assign tmp4838 = s1 ? 1 : tmp4839;
  assign tmp4841 = s0 ? tmp4839 : 1;
  assign tmp4842 = s0 ? 1 : tmp4839;
  assign tmp4840 = s1 ? tmp4841 : tmp4842;
  assign tmp4837 = s2 ? tmp4838 : tmp4840;
  assign tmp4846 = s1 ? tmp4839 : tmp4462;
  assign tmp4848 = s0 ? tmp4839 : tmp4527;
  assign tmp4847 = s1 ? tmp4811 : tmp4848;
  assign tmp4845 = s2 ? tmp4846 : tmp4847;
  assign tmp4851 = ~(s0 ? tmp4568 : tmp4463);
  assign tmp4850 = s1 ? tmp4565 : tmp4851;
  assign tmp4849 = s2 ? tmp4850 : tmp4815;
  assign tmp4844 = s3 ? tmp4845 : tmp4849;
  assign tmp4855 = s0 ? 1 : tmp4578;
  assign tmp4854 = s1 ? tmp4855 : tmp4579;
  assign tmp4858 = ~(l1 ? tmp4554 : 1);
  assign tmp4857 = s0 ? tmp4463 : tmp4858;
  assign tmp4859 = ~(s0 ? tmp4527 : tmp4578);
  assign tmp4856 = ~(s1 ? tmp4857 : tmp4859);
  assign tmp4853 = s2 ? tmp4854 : tmp4856;
  assign tmp4862 = s0 ? tmp4568 : tmp4580;
  assign tmp4863 = s0 ? tmp4580 : tmp4858;
  assign tmp4861 = s1 ? tmp4862 : tmp4863;
  assign tmp4864 = ~(s1 ? tmp4855 : tmp4498);
  assign tmp4860 = ~(s2 ? tmp4861 : tmp4864);
  assign tmp4852 = s3 ? tmp4853 : tmp4860;
  assign tmp4843 = s4 ? tmp4844 : tmp4852;
  assign tmp4836 = ~(s5 ? tmp4837 : tmp4843);
  assign tmp4835 = s6 ? tmp4463 : tmp4836;
  assign tmp4834 = s7 ? tmp4521 : tmp4835;
  assign tmp4833 = ~(s8 ? tmp4834 : tmp4831);
  assign tmp4832 = s9 ? 1 : tmp4833;
  assign tmp4800 = s11 ? tmp4801 : tmp4832;
  assign tmp4868 = s7 ? tmp4597 : tmp4804;
  assign tmp4867 = ~(s8 ? tmp4868 : tmp4831);
  assign tmp4866 = s9 ? 1 : tmp4867;
  assign tmp4875 = l1 ? tmp4673 : 1;
  assign tmp4877 = s0 ? tmp4875 : tmp4673;
  assign tmp4876 = s1 ? tmp4877 : tmp4875;
  assign tmp4874 = s2 ? tmp4875 : tmp4876;
  assign tmp4881 = s1 ? tmp4875 : tmp4462;
  assign tmp4883 = s0 ? tmp4875 : tmp4462;
  assign tmp4884 = s0 ? tmp4875 : tmp4527;
  assign tmp4882 = s1 ? tmp4883 : tmp4884;
  assign tmp4880 = s2 ? tmp4881 : tmp4882;
  assign tmp4887 = s0 ? tmp4527 : tmp4568;
  assign tmp4886 = s1 ? tmp4527 : tmp4887;
  assign tmp4889 = s0 ? tmp4568 : tmp4673;
  assign tmp4890 = s0 ? tmp4673 : 1;
  assign tmp4888 = s1 ? tmp4889 : tmp4890;
  assign tmp4885 = s2 ? tmp4886 : tmp4888;
  assign tmp4879 = s3 ? tmp4880 : tmp4885;
  assign tmp4895 = l1 ? tmp4673 : tmp4498;
  assign tmp4894 = s0 ? tmp4462 : tmp4895;
  assign tmp4893 = s1 ? tmp4811 : tmp4894;
  assign tmp4897 = s0 ? tmp4895 : tmp4875;
  assign tmp4898 = s0 ? tmp4527 : tmp4875;
  assign tmp4896 = s1 ? tmp4897 : tmp4898;
  assign tmp4892 = s2 ? tmp4893 : tmp4896;
  assign tmp4901 = s0 ? tmp4673 : tmp4875;
  assign tmp4900 = s1 ? tmp4898 : tmp4901;
  assign tmp4903 = s0 ? tmp4568 : tmp4895;
  assign tmp4902 = s1 ? tmp4811 : tmp4903;
  assign tmp4899 = s2 ? tmp4900 : tmp4902;
  assign tmp4891 = s3 ? tmp4892 : tmp4899;
  assign tmp4878 = s4 ? tmp4879 : tmp4891;
  assign tmp4873 = ~(s5 ? tmp4874 : tmp4878);
  assign tmp4872 = s6 ? tmp4463 : tmp4873;
  assign tmp4871 = s7 ? tmp4633 : tmp4872;
  assign tmp4910 = s1 ? tmp4875 : 1;
  assign tmp4911 = s0 ? tmp4875 : 1;
  assign tmp4909 = s2 ? tmp4910 : tmp4911;
  assign tmp4913 = s1 ? 1 : tmp4811;
  assign tmp4915 = s0 ? tmp4462 : tmp4673;
  assign tmp4914 = s1 ? tmp4915 : tmp4890;
  assign tmp4912 = s2 ? tmp4913 : tmp4914;
  assign tmp4908 = s3 ? tmp4909 : tmp4912;
  assign tmp4919 = s0 ? 1 : tmp4875;
  assign tmp4918 = s1 ? 1 : tmp4919;
  assign tmp4920 = s1 ? tmp4875 : tmp4919;
  assign tmp4917 = s2 ? tmp4918 : tmp4920;
  assign tmp4922 = s1 ? tmp4919 : tmp4901;
  assign tmp4924 = s0 ? tmp4462 : tmp4875;
  assign tmp4923 = s1 ? 1 : tmp4924;
  assign tmp4921 = s2 ? tmp4922 : tmp4923;
  assign tmp4916 = s3 ? tmp4917 : tmp4921;
  assign tmp4907 = s4 ? tmp4908 : tmp4916;
  assign tmp4906 = s5 ? tmp4874 : tmp4907;
  assign tmp4905 = s6 ? tmp4906 : 1;
  assign tmp4904 = ~(s7 ? tmp4905 : tmp4498);
  assign tmp4870 = ~(s8 ? tmp4871 : tmp4904);
  assign tmp4869 = s9 ? 1 : tmp4870;
  assign tmp4865 = s11 ? tmp4866 : tmp4869;
  assign tmp4799 = s12 ? tmp4800 : tmp4865;
  assign tmp4934 = ~(l2 ? tmp4503 : 0);
  assign tmp4933 = l1 ? 1 : tmp4934;
  assign tmp4936 = s0 ? tmp4933 : tmp4711;
  assign tmp4937 = s0 ? tmp4933 : 1;
  assign tmp4935 = s1 ? tmp4936 : tmp4937;
  assign tmp4932 = s2 ? tmp4933 : tmp4935;
  assign tmp4942 = s0 ? 1 : tmp4933;
  assign tmp4941 = s1 ? tmp4942 : tmp4568;
  assign tmp4944 = s0 ? tmp4933 : tmp4568;
  assign tmp4943 = s1 ? tmp4944 : tmp4936;
  assign tmp4940 = s2 ? tmp4941 : tmp4943;
  assign tmp4946 = s1 ? tmp4714 : tmp4814;
  assign tmp4948 = s0 ? tmp4463 : 0;
  assign tmp4947 = ~(s1 ? tmp4463 : tmp4948);
  assign tmp4945 = s2 ? tmp4946 : tmp4947;
  assign tmp4939 = s3 ? tmp4940 : tmp4945;
  assign tmp4952 = s0 ? tmp4711 : tmp4933;
  assign tmp4951 = s1 ? tmp4952 : tmp4823;
  assign tmp4950 = s2 ? tmp4820 : tmp4951;
  assign tmp4955 = s0 ? tmp4527 : tmp4711;
  assign tmp4956 = ~(s0 ? tmp4463 : 0);
  assign tmp4954 = s1 ? tmp4955 : tmp4956;
  assign tmp4953 = s2 ? tmp4954 : tmp4828;
  assign tmp4949 = s3 ? tmp4950 : tmp4953;
  assign tmp4938 = s4 ? tmp4939 : tmp4949;
  assign tmp4931 = ~(s5 ? tmp4932 : tmp4938);
  assign tmp4930 = s6 ? tmp4463 : tmp4931;
  assign tmp4929 = s7 ? tmp4669 : tmp4930;
  assign tmp4928 = ~(s8 ? tmp4929 : tmp4831);
  assign tmp4927 = s9 ? 1 : tmp4928;
  assign tmp4926 = s11 ? tmp4927 : tmp4801;
  assign tmp4960 = s7 ? tmp4737 : tmp4872;
  assign tmp4959 = ~(s8 ? tmp4960 : tmp4904);
  assign tmp4958 = s9 ? 1 : tmp4959;
  assign tmp4963 = s7 ? tmp4770 : tmp4872;
  assign tmp4962 = ~(s8 ? tmp4963 : tmp4904);
  assign tmp4961 = s9 ? 1 : tmp4962;
  assign tmp4957 = s11 ? tmp4958 : tmp4961;
  assign tmp4925 = s12 ? tmp4926 : tmp4957;
  assign tmp4798 = s13 ? tmp4799 : tmp4925;
  assign tmp4797 = s15 ? tmp4798 : tmp4448;
  assign tmp4447 = ~(s16 ? tmp4448 : tmp4797);
  assign s6n = tmp4447;

  assign tmp4975 = l3 ? 1 : 0;
  assign tmp4974 = l2 ? tmp4975 : 1;
  assign tmp4973 = l1 ? tmp4974 : 1;
  assign tmp4972 = s1 ? tmp4973 : 1;
  assign tmp4978 = l1 ? tmp4974 : tmp4975;
  assign tmp4977 = s0 ? 1 : tmp4978;
  assign tmp4980 = l1 ? tmp4975 : 1;
  assign tmp4979 = s0 ? tmp4980 : 1;
  assign tmp4976 = s1 ? tmp4977 : tmp4979;
  assign tmp4971 = s2 ? tmp4972 : tmp4976;
  assign tmp4987 = l2 ? 1 : tmp4975;
  assign tmp4988 = ~(l2 ? tmp4975 : 0);
  assign tmp4986 = l1 ? tmp4987 : tmp4988;
  assign tmp4985 = s0 ? tmp4986 : 1;
  assign tmp4990 = l2 ? tmp4975 : 0;
  assign tmp4989 = l1 ? tmp4990 : tmp4975;
  assign tmp4984 = s1 ? tmp4985 : tmp4989;
  assign tmp4993 = l1 ? tmp4975 : tmp4990;
  assign tmp4992 = s0 ? 1 : tmp4993;
  assign tmp4991 = s1 ? tmp4973 : tmp4992;
  assign tmp4983 = s2 ? tmp4984 : tmp4991;
  assign tmp4996 = s0 ? tmp4993 : 1;
  assign tmp4995 = s1 ? tmp4996 : 1;
  assign tmp4994 = s2 ? tmp4995 : 1;
  assign tmp4982 = s3 ? tmp4983 : tmp4994;
  assign tmp5001 = ~(l1 ? tmp4990 : tmp4975);
  assign tmp5000 = s0 ? tmp4993 : tmp5001;
  assign tmp4999 = s1 ? 1 : tmp5000;
  assign tmp4998 = s2 ? 1 : tmp4999;
  assign tmp4997 = s3 ? tmp4998 : 1;
  assign tmp4981 = s4 ? tmp4982 : tmp4997;
  assign tmp4970 = s5 ? tmp4971 : tmp4981;
  assign tmp5010 = s0 ? tmp4973 : tmp4989;
  assign tmp5009 = s1 ? tmp5010 : tmp4992;
  assign tmp5008 = s2 ? tmp4984 : tmp5009;
  assign tmp5007 = s3 ? tmp5008 : tmp4994;
  assign tmp5006 = s4 ? tmp5007 : tmp4997;
  assign tmp5005 = s5 ? tmp4971 : tmp5006;
  assign tmp5004 = s6 ? tmp5005 : tmp4970;
  assign tmp5014 = s3 ? tmp4983 : 1;
  assign tmp5017 = s1 ? 1 : tmp5001;
  assign tmp5016 = s2 ? 1 : tmp5017;
  assign tmp5015 = s3 ? tmp5016 : 1;
  assign tmp5013 = s4 ? tmp5014 : tmp5015;
  assign tmp5012 = s5 ? tmp4971 : tmp5013;
  assign tmp5011 = s6 ? tmp5012 : tmp5005;
  assign tmp5003 = s7 ? tmp5004 : tmp5011;
  assign tmp5021 = s4 ? tmp4982 : tmp5015;
  assign tmp5020 = s5 ? tmp4971 : tmp5021;
  assign tmp5019 = s6 ? tmp5005 : tmp5020;
  assign tmp5022 = s6 ? tmp5020 : tmp5012;
  assign tmp5018 = s7 ? tmp5019 : tmp5022;
  assign tmp5002 = s8 ? tmp5003 : tmp5018;
  assign tmp4969 = s9 ? tmp4970 : tmp5002;
  assign tmp5026 = s6 ? tmp4970 : tmp5012;
  assign tmp5025 = s7 ? tmp5004 : tmp5026;
  assign tmp5024 = s8 ? tmp5003 : tmp5025;
  assign tmp5023 = s9 ? tmp4970 : tmp5024;
  assign tmp4968 = s10 ? tmp4969 : tmp5023;
  assign tmp5031 = s3 ? tmp5008 : 1;
  assign tmp5030 = s4 ? tmp5031 : tmp5015;
  assign tmp5029 = s5 ? tmp4971 : tmp5030;
  assign tmp5034 = s6 ? tmp5005 : tmp5029;
  assign tmp5033 = s7 ? tmp5034 : tmp5011;
  assign tmp5036 = s6 ? tmp5005 : tmp5012;
  assign tmp5035 = s7 ? tmp5036 : tmp5012;
  assign tmp5032 = s8 ? tmp5033 : tmp5035;
  assign tmp5028 = s9 ? tmp5029 : tmp5032;
  assign tmp5040 = s6 ? tmp5029 : tmp5012;
  assign tmp5039 = s7 ? tmp5034 : tmp5040;
  assign tmp5038 = s8 ? tmp5033 : tmp5039;
  assign tmp5037 = s9 ? tmp5029 : tmp5038;
  assign tmp5027 = s10 ? tmp5028 : tmp5037;
  assign tmp4967 = s11 ? tmp4968 : tmp5027;
  assign tmp5044 = s7 ? tmp5005 : tmp5011;
  assign tmp5043 = s8 ? tmp5044 : tmp5018;
  assign tmp5042 = s9 ? tmp5005 : tmp5043;
  assign tmp5047 = s7 ? tmp5005 : tmp5036;
  assign tmp5046 = s8 ? tmp5044 : tmp5047;
  assign tmp5045 = s9 ? tmp5005 : tmp5046;
  assign tmp5041 = s10 ? tmp5042 : tmp5045;
  assign tmp4966 = s12 ? tmp4967 : tmp5041;
  assign tmp5052 = s7 ? tmp5036 : tmp5011;
  assign tmp5051 = s8 ? tmp5052 : tmp5035;
  assign tmp5050 = s9 ? tmp5012 : tmp5051;
  assign tmp5049 = s11 ? tmp5050 : tmp4968;
  assign tmp5053 = s11 ? tmp5027 : tmp4968;
  assign tmp5048 = s12 ? tmp5049 : tmp5053;
  assign tmp4965 = s13 ? tmp4966 : tmp5048;
  assign tmp5061 = s7 ? tmp5036 : tmp5022;
  assign tmp5060 = s8 ? tmp5003 : tmp5061;
  assign tmp5059 = s9 ? tmp5012 : tmp5060;
  assign tmp5064 = s7 ? tmp5036 : tmp5026;
  assign tmp5063 = s8 ? tmp5003 : tmp5064;
  assign tmp5062 = s9 ? tmp5012 : tmp5063;
  assign tmp5058 = s10 ? tmp5059 : tmp5062;
  assign tmp5066 = s9 ? tmp5012 : tmp5032;
  assign tmp5069 = s7 ? tmp5036 : tmp5040;
  assign tmp5068 = s8 ? tmp5033 : tmp5069;
  assign tmp5067 = s9 ? tmp5012 : tmp5068;
  assign tmp5065 = s10 ? tmp5066 : tmp5067;
  assign tmp5057 = s11 ? tmp5058 : tmp5065;
  assign tmp5072 = s8 ? tmp5044 : tmp5061;
  assign tmp5071 = s9 ? tmp5012 : tmp5072;
  assign tmp5074 = s8 ? tmp5044 : tmp5036;
  assign tmp5073 = s9 ? tmp5012 : tmp5074;
  assign tmp5070 = s10 ? tmp5071 : tmp5073;
  assign tmp5056 = s12 ? tmp5057 : tmp5070;
  assign tmp5076 = s11 ? tmp5050 : tmp5058;
  assign tmp5077 = s11 ? tmp5065 : tmp5058;
  assign tmp5075 = s12 ? tmp5076 : tmp5077;
  assign tmp5055 = s13 ? tmp5056 : tmp5075;
  assign tmp5085 = s6 ? tmp4970 : tmp5005;
  assign tmp5084 = s7 ? tmp5004 : tmp5085;
  assign tmp5086 = s7 ? tmp5019 : tmp5020;
  assign tmp5083 = s8 ? tmp5084 : tmp5086;
  assign tmp5082 = s9 ? tmp4970 : tmp5083;
  assign tmp5089 = s7 ? tmp5004 : tmp4970;
  assign tmp5088 = s8 ? tmp5084 : tmp5089;
  assign tmp5087 = s9 ? tmp4970 : tmp5088;
  assign tmp5081 = s10 ? tmp5082 : tmp5087;
  assign tmp5094 = s6 ? tmp5029 : tmp5005;
  assign tmp5093 = s7 ? tmp5034 : tmp5094;
  assign tmp5092 = s8 ? tmp5093 : tmp5035;
  assign tmp5091 = s9 ? tmp5029 : tmp5092;
  assign tmp5097 = s7 ? tmp5034 : tmp5029;
  assign tmp5096 = s8 ? tmp5093 : tmp5097;
  assign tmp5095 = s9 ? tmp5029 : tmp5096;
  assign tmp5090 = s10 ? tmp5091 : tmp5095;
  assign tmp5080 = s11 ? tmp5081 : tmp5090;
  assign tmp5079 = s12 ? tmp5080 : tmp5041;
  assign tmp5078 = s13 ? tmp5079 : tmp5048;
  assign tmp5054 = s15 ? tmp5055 : tmp5078;
  assign tmp4964 = ~(s16 ? tmp4965 : tmp5054);
  assign s5n = tmp4964;

  assign tmp5117 = l3 ? 1 : 0;
  assign tmp5118 = ~(l3 ? 1 : 0);
  assign tmp5116 = l2 ? tmp5117 : tmp5118;
  assign tmp5119 = l2 ? 1 : tmp5117;
  assign tmp5115 = ~(l1 ? tmp5116 : tmp5119);
  assign tmp5114 = s0 ? 1 : tmp5115;
  assign tmp5113 = s1 ? tmp5114 : tmp5115;
  assign tmp5122 = l1 ? tmp5116 : tmp5119;
  assign tmp5123 = l1 ? tmp5116 : tmp5117;
  assign tmp5121 = s0 ? tmp5122 : tmp5123;
  assign tmp5126 = l2 ? tmp5117 : 0;
  assign tmp5125 = l1 ? tmp5126 : tmp5119;
  assign tmp5124 = s0 ? tmp5125 : tmp5122;
  assign tmp5120 = ~(s1 ? tmp5121 : tmp5124);
  assign tmp5112 = s2 ? tmp5113 : tmp5120;
  assign tmp5111 = s3 ? 1 : tmp5112;
  assign tmp5110 = s4 ? 1 : tmp5111;
  assign tmp5133 = ~(l2 ? tmp5117 : tmp5118);
  assign tmp5132 = l1 ? tmp5126 : tmp5133;
  assign tmp5131 = s0 ? tmp5132 : tmp5122;
  assign tmp5135 = l1 ? tmp5126 : tmp5117;
  assign tmp5134 = s0 ? tmp5135 : 0;
  assign tmp5130 = s1 ? tmp5131 : tmp5134;
  assign tmp5137 = s0 ? tmp5122 : 0;
  assign tmp5138 = s0 ? tmp5122 : tmp5126;
  assign tmp5136 = s1 ? tmp5137 : tmp5138;
  assign tmp5129 = s2 ? tmp5130 : tmp5136;
  assign tmp5143 = ~(l2 ? tmp5117 : 0);
  assign tmp5142 = l1 ? 1 : tmp5143;
  assign tmp5144 = ~(l1 ? tmp5116 : 1);
  assign tmp5141 = s0 ? tmp5142 : tmp5144;
  assign tmp5147 = l2 ? tmp5117 : 1;
  assign tmp5146 = l1 ? tmp5116 : tmp5147;
  assign tmp5149 = l2 ? 1 : tmp5118;
  assign tmp5148 = ~(l1 ? tmp5119 : tmp5149);
  assign tmp5145 = ~(s0 ? tmp5146 : tmp5148);
  assign tmp5140 = s1 ? tmp5141 : tmp5145;
  assign tmp5152 = ~(l1 ? tmp5149 : 1);
  assign tmp5151 = s0 ? 1 : tmp5152;
  assign tmp5154 = ~(l1 ? tmp5126 : tmp5133);
  assign tmp5153 = s0 ? 1 : tmp5154;
  assign tmp5150 = s1 ? tmp5151 : tmp5153;
  assign tmp5139 = ~(s2 ? tmp5140 : tmp5150);
  assign tmp5128 = s3 ? tmp5129 : tmp5139;
  assign tmp5159 = l1 ? 1 : tmp5147;
  assign tmp5158 = s0 ? 1 : tmp5159;
  assign tmp5161 = l1 ? tmp5119 : 1;
  assign tmp5160 = s0 ? 1 : tmp5161;
  assign tmp5157 = s1 ? tmp5158 : tmp5160;
  assign tmp5164 = l1 ? tmp5119 : tmp5147;
  assign tmp5163 = s0 ? tmp5142 : tmp5164;
  assign tmp5162 = s1 ? tmp5114 : tmp5163;
  assign tmp5156 = s2 ? tmp5157 : tmp5162;
  assign tmp5167 = s0 ? tmp5146 : tmp5122;
  assign tmp5168 = ~(s0 ? 1 : tmp5115);
  assign tmp5166 = s1 ? tmp5167 : tmp5168;
  assign tmp5165 = ~(s2 ? tmp5166 : 0);
  assign tmp5155 = ~(s3 ? tmp5156 : tmp5165);
  assign tmp5127 = ~(s4 ? tmp5128 : tmp5155);
  assign tmp5109 = s5 ? tmp5110 : tmp5127;
  assign tmp5108 = s6 ? 1 : tmp5109;
  assign tmp5107 = s7 ? 1 : tmp5108;
  assign tmp5106 = s8 ? 1 : tmp5107;
  assign tmp5178 = ~(l1 ? 1 : tmp5143);
  assign tmp5177 = s0 ? tmp5135 : tmp5178;
  assign tmp5176 = s1 ? tmp5131 : tmp5177;
  assign tmp5180 = s0 ? tmp5122 : tmp5178;
  assign tmp5179 = s1 ? tmp5180 : tmp5138;
  assign tmp5175 = s2 ? tmp5176 : tmp5179;
  assign tmp5185 = l2 ? 1 : 0;
  assign tmp5184 = l1 ? tmp5185 : tmp5149;
  assign tmp5183 = ~(s0 ? tmp5184 : tmp5132);
  assign tmp5182 = s1 ? tmp5151 : tmp5183;
  assign tmp5181 = ~(s2 ? tmp5140 : tmp5182);
  assign tmp5174 = s3 ? tmp5175 : tmp5181;
  assign tmp5189 = s0 ? tmp5184 : tmp5122;
  assign tmp5188 = s1 ? tmp5167 : tmp5189;
  assign tmp5187 = ~(s2 ? tmp5188 : 0);
  assign tmp5186 = ~(s3 ? tmp5156 : tmp5187);
  assign tmp5173 = ~(s4 ? tmp5174 : tmp5186);
  assign tmp5172 = s5 ? tmp5110 : tmp5173;
  assign tmp5171 = s6 ? tmp5172 : tmp5109;
  assign tmp5196 = s0 ? 1 : tmp5144;
  assign tmp5198 = l1 ? tmp5119 : tmp5149;
  assign tmp5197 = s0 ? 1 : tmp5198;
  assign tmp5195 = s1 ? tmp5196 : tmp5197;
  assign tmp5194 = ~(s2 ? tmp5195 : tmp5150);
  assign tmp5193 = s3 ? tmp5129 : tmp5194;
  assign tmp5202 = s0 ? 1 : tmp5164;
  assign tmp5201 = s1 ? tmp5114 : tmp5202;
  assign tmp5200 = s2 ? tmp5157 : tmp5201;
  assign tmp5203 = s2 ? tmp5114 : 1;
  assign tmp5199 = ~(s3 ? tmp5200 : tmp5203);
  assign tmp5192 = ~(s4 ? tmp5193 : tmp5199);
  assign tmp5191 = s5 ? tmp5110 : tmp5192;
  assign tmp5190 = s6 ? tmp5191 : tmp5172;
  assign tmp5170 = s7 ? tmp5171 : tmp5190;
  assign tmp5207 = ~(s4 ? tmp5128 : tmp5199);
  assign tmp5206 = s5 ? tmp5110 : tmp5207;
  assign tmp5205 = s6 ? tmp5172 : tmp5206;
  assign tmp5208 = s6 ? tmp5206 : tmp5191;
  assign tmp5204 = s7 ? tmp5205 : tmp5208;
  assign tmp5169 = s8 ? tmp5170 : tmp5204;
  assign tmp5105 = s9 ? tmp5106 : tmp5169;
  assign tmp5212 = s6 ? tmp5109 : tmp5191;
  assign tmp5211 = s7 ? tmp5171 : tmp5212;
  assign tmp5210 = s8 ? tmp5170 : tmp5211;
  assign tmp5209 = s9 ? tmp5106 : tmp5210;
  assign tmp5104 = s10 ? tmp5105 : tmp5209;
  assign tmp5224 = ~(l1 ? tmp5147 : tmp5119);
  assign tmp5223 = s0 ? 1 : tmp5224;
  assign tmp5222 = s1 ? tmp5223 : tmp5224;
  assign tmp5227 = l1 ? tmp5147 : tmp5119;
  assign tmp5228 = l1 ? tmp5147 : tmp5117;
  assign tmp5226 = s0 ? tmp5227 : tmp5228;
  assign tmp5230 = l1 ? tmp5117 : tmp5119;
  assign tmp5229 = s0 ? tmp5230 : tmp5227;
  assign tmp5225 = ~(s1 ? tmp5226 : tmp5229);
  assign tmp5221 = s2 ? tmp5222 : tmp5225;
  assign tmp5220 = s3 ? 1 : tmp5221;
  assign tmp5219 = s4 ? 1 : tmp5220;
  assign tmp5236 = l1 ? tmp5117 : tmp5133;
  assign tmp5235 = s0 ? tmp5236 : tmp5227;
  assign tmp5234 = s1 ? tmp5235 : tmp5177;
  assign tmp5238 = s0 ? tmp5227 : tmp5178;
  assign tmp5240 = l1 ? tmp5117 : tmp5126;
  assign tmp5239 = s0 ? tmp5227 : tmp5240;
  assign tmp5237 = s1 ? tmp5238 : tmp5239;
  assign tmp5233 = s2 ? tmp5234 : tmp5237;
  assign tmp5244 = ~(l1 ? tmp5147 : 1);
  assign tmp5243 = s0 ? 1 : tmp5244;
  assign tmp5242 = s1 ? tmp5243 : tmp5197;
  assign tmp5246 = s0 ? 1 : 0;
  assign tmp5248 = ~(l1 ? tmp5117 : tmp5133);
  assign tmp5247 = s0 ? 1 : tmp5248;
  assign tmp5245 = s1 ? tmp5246 : tmp5247;
  assign tmp5241 = ~(s2 ? tmp5242 : tmp5245);
  assign tmp5232 = s3 ? tmp5233 : tmp5241;
  assign tmp5253 = l1 ? tmp5185 : 1;
  assign tmp5252 = s0 ? 1 : tmp5253;
  assign tmp5251 = s1 ? tmp5158 : tmp5252;
  assign tmp5256 = l1 ? tmp5185 : tmp5147;
  assign tmp5255 = s0 ? 1 : tmp5256;
  assign tmp5254 = s1 ? tmp5223 : tmp5255;
  assign tmp5250 = s2 ? tmp5251 : tmp5254;
  assign tmp5257 = s2 ? tmp5223 : 1;
  assign tmp5249 = ~(s3 ? tmp5250 : tmp5257);
  assign tmp5231 = ~(s4 ? tmp5232 : tmp5249);
  assign tmp5218 = s5 ? tmp5219 : tmp5231;
  assign tmp5217 = s6 ? 1 : tmp5218;
  assign tmp5216 = s7 ? 1 : tmp5217;
  assign tmp5215 = s8 ? 1 : tmp5216;
  assign tmp5260 = s6 ? tmp5172 : tmp5218;
  assign tmp5266 = s1 ? tmp5235 : tmp5134;
  assign tmp5268 = s0 ? tmp5227 : 0;
  assign tmp5267 = s1 ? tmp5268 : tmp5239;
  assign tmp5265 = s2 ? tmp5266 : tmp5267;
  assign tmp5264 = s3 ? tmp5265 : tmp5241;
  assign tmp5263 = ~(s4 ? tmp5264 : tmp5249);
  assign tmp5262 = s5 ? tmp5219 : tmp5263;
  assign tmp5261 = s6 ? tmp5262 : tmp5172;
  assign tmp5259 = s7 ? tmp5260 : tmp5261;
  assign tmp5274 = s2 ? tmp5234 : tmp5267;
  assign tmp5273 = s3 ? tmp5274 : tmp5241;
  assign tmp5272 = ~(s4 ? tmp5273 : tmp5249);
  assign tmp5271 = s5 ? tmp5219 : tmp5272;
  assign tmp5270 = s6 ? tmp5172 : tmp5271;
  assign tmp5275 = s6 ? tmp5271 : tmp5262;
  assign tmp5269 = s7 ? tmp5270 : tmp5275;
  assign tmp5258 = s8 ? tmp5259 : tmp5269;
  assign tmp5214 = s9 ? tmp5215 : tmp5258;
  assign tmp5279 = s6 ? tmp5218 : tmp5262;
  assign tmp5278 = s7 ? tmp5260 : tmp5279;
  assign tmp5277 = s8 ? tmp5259 : tmp5278;
  assign tmp5276 = s9 ? tmp5215 : tmp5277;
  assign tmp5213 = s10 ? tmp5214 : tmp5276;
  assign tmp5103 = s11 ? tmp5104 : tmp5213;
  assign tmp5288 = s3 ? tmp5175 : tmp5139;
  assign tmp5287 = ~(s4 ? tmp5288 : tmp5155);
  assign tmp5286 = s5 ? tmp5110 : tmp5287;
  assign tmp5285 = s6 ? 1 : tmp5286;
  assign tmp5284 = s7 ? 1 : tmp5285;
  assign tmp5283 = s8 ? 1 : tmp5284;
  assign tmp5291 = s6 ? tmp5172 : tmp5286;
  assign tmp5290 = s7 ? tmp5291 : tmp5190;
  assign tmp5297 = s2 ? tmp5176 : tmp5136;
  assign tmp5296 = s3 ? tmp5297 : tmp5139;
  assign tmp5295 = ~(s4 ? tmp5296 : tmp5199);
  assign tmp5294 = s5 ? tmp5110 : tmp5295;
  assign tmp5293 = s6 ? tmp5172 : tmp5294;
  assign tmp5298 = s6 ? tmp5294 : tmp5191;
  assign tmp5292 = s7 ? tmp5293 : tmp5298;
  assign tmp5289 = s8 ? tmp5290 : tmp5292;
  assign tmp5282 = s9 ? tmp5283 : tmp5289;
  assign tmp5302 = s6 ? tmp5286 : tmp5191;
  assign tmp5301 = s7 ? tmp5291 : tmp5302;
  assign tmp5300 = s8 ? tmp5290 : tmp5301;
  assign tmp5299 = s9 ? tmp5283 : tmp5300;
  assign tmp5281 = s10 ? tmp5282 : tmp5299;
  assign tmp5307 = s6 ? 1 : tmp5172;
  assign tmp5306 = s7 ? 1 : tmp5307;
  assign tmp5305 = s8 ? 1 : tmp5306;
  assign tmp5309 = s7 ? tmp5172 : tmp5190;
  assign tmp5314 = s3 ? tmp5297 : tmp5181;
  assign tmp5313 = ~(s4 ? tmp5314 : tmp5199);
  assign tmp5312 = s5 ? tmp5110 : tmp5313;
  assign tmp5311 = s6 ? tmp5172 : tmp5312;
  assign tmp5315 = s6 ? tmp5312 : tmp5191;
  assign tmp5310 = s7 ? tmp5311 : tmp5315;
  assign tmp5308 = s8 ? tmp5309 : tmp5310;
  assign tmp5304 = s9 ? tmp5305 : tmp5308;
  assign tmp5319 = s6 ? tmp5172 : tmp5191;
  assign tmp5318 = s7 ? tmp5172 : tmp5319;
  assign tmp5317 = s8 ? tmp5309 : tmp5318;
  assign tmp5316 = s9 ? tmp5305 : tmp5317;
  assign tmp5303 = s10 ? tmp5304 : tmp5316;
  assign tmp5280 = s11 ? tmp5281 : tmp5303;
  assign tmp5102 = s12 ? tmp5103 : tmp5280;
  assign tmp5325 = s6 ? 1 : tmp5262;
  assign tmp5324 = s7 ? 1 : tmp5325;
  assign tmp5323 = s8 ? 1 : tmp5324;
  assign tmp5328 = s6 ? tmp5172 : tmp5262;
  assign tmp5327 = s7 ? tmp5328 : tmp5261;
  assign tmp5329 = s7 ? tmp5328 : tmp5262;
  assign tmp5326 = s8 ? tmp5327 : tmp5329;
  assign tmp5322 = s9 ? tmp5323 : tmp5326;
  assign tmp5321 = s11 ? tmp5322 : tmp5104;
  assign tmp5330 = s11 ? tmp5213 : tmp5104;
  assign tmp5320 = s12 ? tmp5321 : tmp5330;
  assign tmp5101 = s13 ? tmp5102 : tmp5320;
  assign tmp5100 = s14 ? 1 : tmp5101;
  assign tmp5099 = s15 ? 1 : tmp5100;
  assign tmp5339 = s7 ? tmp5171 : tmp5261;
  assign tmp5347 = s0 ? tmp5142 : tmp5244;
  assign tmp5346 = s1 ? tmp5347 : tmp5145;
  assign tmp5349 = ~(s0 ? tmp5184 : tmp5236);
  assign tmp5348 = s1 ? tmp5246 : tmp5349;
  assign tmp5345 = ~(s2 ? tmp5346 : tmp5348);
  assign tmp5344 = s3 ? tmp5233 : tmp5345;
  assign tmp5353 = s0 ? tmp5142 : tmp5256;
  assign tmp5352 = s1 ? tmp5223 : tmp5353;
  assign tmp5351 = s2 ? tmp5251 : tmp5352;
  assign tmp5356 = s0 ? tmp5146 : tmp5227;
  assign tmp5357 = s0 ? tmp5184 : tmp5227;
  assign tmp5355 = s1 ? tmp5356 : tmp5357;
  assign tmp5354 = ~(s2 ? tmp5355 : 0);
  assign tmp5350 = ~(s3 ? tmp5351 : tmp5354);
  assign tmp5343 = ~(s4 ? tmp5344 : tmp5350);
  assign tmp5342 = s5 ? tmp5219 : tmp5343;
  assign tmp5341 = s6 ? tmp5342 : tmp5262;
  assign tmp5358 = s6 ? tmp5206 : tmp5262;
  assign tmp5340 = s7 ? tmp5341 : tmp5358;
  assign tmp5338 = s8 ? tmp5339 : tmp5340;
  assign tmp5337 = s9 ? tmp5323 : tmp5338;
  assign tmp5362 = s6 ? tmp5109 : tmp5262;
  assign tmp5361 = s7 ? tmp5341 : tmp5362;
  assign tmp5360 = s8 ? tmp5339 : tmp5361;
  assign tmp5359 = s9 ? tmp5323 : tmp5360;
  assign tmp5336 = s10 ? tmp5337 : tmp5359;
  assign tmp5366 = s7 ? tmp5341 : tmp5275;
  assign tmp5365 = s8 ? tmp5259 : tmp5366;
  assign tmp5364 = s9 ? tmp5323 : tmp5365;
  assign tmp5369 = s7 ? tmp5341 : tmp5279;
  assign tmp5368 = s8 ? tmp5259 : tmp5369;
  assign tmp5367 = s9 ? tmp5323 : tmp5368;
  assign tmp5363 = s10 ? tmp5364 : tmp5367;
  assign tmp5335 = s11 ? tmp5336 : tmp5363;
  assign tmp5374 = s7 ? tmp5291 : tmp5261;
  assign tmp5376 = s6 ? tmp5294 : tmp5262;
  assign tmp5375 = s7 ? tmp5341 : tmp5376;
  assign tmp5373 = s8 ? tmp5374 : tmp5375;
  assign tmp5372 = s9 ? tmp5323 : tmp5373;
  assign tmp5380 = s6 ? tmp5286 : tmp5262;
  assign tmp5379 = s7 ? tmp5341 : tmp5380;
  assign tmp5378 = s8 ? tmp5374 : tmp5379;
  assign tmp5377 = s9 ? tmp5323 : tmp5378;
  assign tmp5371 = s10 ? tmp5372 : tmp5377;
  assign tmp5384 = s7 ? tmp5172 : tmp5261;
  assign tmp5386 = s6 ? tmp5312 : tmp5262;
  assign tmp5385 = s7 ? tmp5328 : tmp5386;
  assign tmp5383 = s8 ? tmp5384 : tmp5385;
  assign tmp5382 = s9 ? tmp5323 : tmp5383;
  assign tmp5388 = s8 ? tmp5384 : tmp5328;
  assign tmp5387 = s9 ? tmp5323 : tmp5388;
  assign tmp5381 = s10 ? tmp5382 : tmp5387;
  assign tmp5370 = s11 ? tmp5371 : tmp5381;
  assign tmp5334 = s12 ? tmp5335 : tmp5370;
  assign tmp5393 = s7 ? tmp5341 : tmp5262;
  assign tmp5392 = s8 ? tmp5327 : tmp5393;
  assign tmp5391 = s9 ? tmp5323 : tmp5392;
  assign tmp5390 = s11 ? tmp5391 : tmp5336;
  assign tmp5398 = s7 ? tmp5328 : tmp5275;
  assign tmp5397 = s8 ? tmp5259 : tmp5398;
  assign tmp5396 = s9 ? tmp5323 : tmp5397;
  assign tmp5401 = s7 ? tmp5328 : tmp5279;
  assign tmp5400 = s8 ? tmp5259 : tmp5401;
  assign tmp5399 = s9 ? tmp5323 : tmp5400;
  assign tmp5395 = s10 ? tmp5396 : tmp5399;
  assign tmp5405 = s7 ? tmp5328 : tmp5358;
  assign tmp5404 = s8 ? tmp5339 : tmp5405;
  assign tmp5403 = s9 ? tmp5323 : tmp5404;
  assign tmp5408 = s7 ? tmp5328 : tmp5362;
  assign tmp5407 = s8 ? tmp5339 : tmp5408;
  assign tmp5406 = s9 ? tmp5323 : tmp5407;
  assign tmp5402 = s10 ? tmp5403 : tmp5406;
  assign tmp5394 = s11 ? tmp5395 : tmp5402;
  assign tmp5389 = s12 ? tmp5390 : tmp5394;
  assign tmp5333 = s13 ? tmp5334 : tmp5389;
  assign tmp5332 = s14 ? 1 : tmp5333;
  assign tmp5422 = s1 ? tmp5141 : tmp5197;
  assign tmp5421 = ~(s2 ? tmp5422 : tmp5150);
  assign tmp5420 = s3 ? tmp5129 : tmp5421;
  assign tmp5423 = ~(s3 ? tmp5156 : tmp5203);
  assign tmp5419 = ~(s4 ? tmp5420 : tmp5423);
  assign tmp5418 = s5 ? tmp5110 : tmp5419;
  assign tmp5417 = s6 ? tmp5418 : tmp5172;
  assign tmp5416 = s7 ? tmp5171 : tmp5417;
  assign tmp5427 = ~(s4 ? tmp5420 : tmp5199);
  assign tmp5426 = s5 ? tmp5110 : tmp5427;
  assign tmp5425 = s6 ? tmp5206 : tmp5426;
  assign tmp5424 = s7 ? tmp5205 : tmp5425;
  assign tmp5415 = s8 ? tmp5416 : tmp5424;
  assign tmp5414 = s9 ? tmp5106 : tmp5415;
  assign tmp5431 = s6 ? tmp5109 : tmp5418;
  assign tmp5430 = s7 ? tmp5171 : tmp5431;
  assign tmp5429 = s8 ? tmp5416 : tmp5430;
  assign tmp5428 = s9 ? tmp5106 : tmp5429;
  assign tmp5413 = s10 ? tmp5414 : tmp5428;
  assign tmp5436 = s6 ? tmp5218 : tmp5172;
  assign tmp5435 = s7 ? tmp5260 : tmp5436;
  assign tmp5437 = s7 ? tmp5270 : tmp5271;
  assign tmp5434 = s8 ? tmp5435 : tmp5437;
  assign tmp5433 = s9 ? tmp5215 : tmp5434;
  assign tmp5440 = s7 ? tmp5260 : tmp5218;
  assign tmp5439 = s8 ? tmp5435 : tmp5440;
  assign tmp5438 = s9 ? tmp5215 : tmp5439;
  assign tmp5432 = s10 ? tmp5433 : tmp5438;
  assign tmp5412 = s11 ? tmp5413 : tmp5432;
  assign tmp5450 = ~(s2 ? tmp5195 : tmp5182);
  assign tmp5449 = s3 ? tmp5129 : tmp5450;
  assign tmp5454 = ~(s0 ? tmp5184 : tmp5122);
  assign tmp5453 = s1 ? tmp5114 : tmp5454;
  assign tmp5452 = s2 ? tmp5453 : 1;
  assign tmp5451 = ~(s3 ? tmp5200 : tmp5452);
  assign tmp5448 = ~(s4 ? tmp5449 : tmp5451);
  assign tmp5447 = s5 ? tmp5110 : tmp5448;
  assign tmp5446 = s6 ? tmp5447 : tmp5172;
  assign tmp5445 = s7 ? tmp5172 : tmp5446;
  assign tmp5458 = ~(s4 ? tmp5449 : tmp5199);
  assign tmp5457 = s5 ? tmp5110 : tmp5458;
  assign tmp5456 = s6 ? tmp5312 : tmp5457;
  assign tmp5455 = s7 ? tmp5311 : tmp5456;
  assign tmp5444 = s8 ? tmp5445 : tmp5455;
  assign tmp5443 = s9 ? tmp5305 : tmp5444;
  assign tmp5462 = s6 ? tmp5172 : tmp5447;
  assign tmp5461 = s7 ? tmp5172 : tmp5462;
  assign tmp5460 = s8 ? tmp5445 : tmp5461;
  assign tmp5459 = s9 ? tmp5305 : tmp5460;
  assign tmp5442 = s10 ? tmp5443 : tmp5459;
  assign tmp5441 = s11 ? tmp5281 : tmp5442;
  assign tmp5411 = s12 ? tmp5412 : tmp5441;
  assign tmp5474 = s1 ? tmp5196 : tmp5145;
  assign tmp5473 = ~(s2 ? tmp5474 : tmp5150);
  assign tmp5472 = s3 ? tmp5129 : tmp5473;
  assign tmp5475 = ~(s3 ? tmp5200 : tmp5165);
  assign tmp5471 = ~(s4 ? tmp5472 : tmp5475);
  assign tmp5470 = s5 ? tmp5110 : tmp5471;
  assign tmp5469 = s6 ? tmp5470 : tmp5172;
  assign tmp5468 = s7 ? tmp5171 : tmp5469;
  assign tmp5479 = ~(s4 ? tmp5472 : tmp5199);
  assign tmp5478 = s5 ? tmp5110 : tmp5479;
  assign tmp5477 = s6 ? tmp5206 : tmp5478;
  assign tmp5476 = s7 ? tmp5205 : tmp5477;
  assign tmp5467 = s8 ? tmp5468 : tmp5476;
  assign tmp5466 = s9 ? tmp5106 : tmp5467;
  assign tmp5483 = s6 ? tmp5109 : tmp5470;
  assign tmp5482 = s7 ? tmp5171 : tmp5483;
  assign tmp5481 = s8 ? tmp5468 : tmp5482;
  assign tmp5480 = s9 ? tmp5106 : tmp5481;
  assign tmp5465 = s10 ? tmp5466 : tmp5480;
  assign tmp5464 = s11 ? tmp5322 : tmp5465;
  assign tmp5463 = s12 ? tmp5464 : tmp5330;
  assign tmp5410 = s13 ? tmp5411 : tmp5463;
  assign tmp5409 = s14 ? 1 : tmp5410;
  assign tmp5331 = s15 ? tmp5332 : tmp5409;
  assign tmp5098 = ~(s16 ? tmp5099 : tmp5331);
  assign s4n = tmp5098;

  assign tmp5495 = ~(l3 ? 1 : 0);
  assign tmp5494 = l2 ? 1 : tmp5495;
  assign tmp5497 = l3 ? 1 : 0;
  assign tmp5496 = ~(l2 ? tmp5497 : tmp5495);
  assign tmp5493 = l1 ? tmp5494 : tmp5496;
  assign tmp5499 = l2 ? tmp5497 : tmp5495;
  assign tmp5498 = l1 ? tmp5499 : tmp5496;
  assign tmp5492 = s1 ? tmp5493 : tmp5498;
  assign tmp5503 = ~(l2 ? tmp5497 : 0);
  assign tmp5502 = l1 ? tmp5494 : tmp5503;
  assign tmp5501 = s0 ? tmp5498 : tmp5502;
  assign tmp5504 = s0 ? tmp5493 : tmp5498;
  assign tmp5500 = s1 ? tmp5501 : tmp5504;
  assign tmp5491 = s2 ? tmp5492 : tmp5500;
  assign tmp5511 = l2 ? 1 : tmp5497;
  assign tmp5510 = l1 ? tmp5499 : tmp5511;
  assign tmp5509 = s0 ? tmp5510 : tmp5498;
  assign tmp5508 = s1 ? tmp5509 : tmp5503;
  assign tmp5512 = s1 ? tmp5493 : tmp5501;
  assign tmp5507 = s2 ? tmp5508 : tmp5512;
  assign tmp5516 = l2 ? tmp5497 : 0;
  assign tmp5518 = l2 ? tmp5497 : 1;
  assign tmp5517 = l1 ? 1 : tmp5518;
  assign tmp5515 = s0 ? tmp5516 : tmp5517;
  assign tmp5520 = l1 ? tmp5499 : tmp5518;
  assign tmp5521 = ~(l1 ? 1 : tmp5511);
  assign tmp5519 = s0 ? tmp5520 : tmp5521;
  assign tmp5514 = s1 ? tmp5515 : tmp5519;
  assign tmp5523 = l1 ? tmp5511 : tmp5494;
  assign tmp5524 = ~(l1 ? tmp5516 : tmp5496);
  assign tmp5522 = s1 ? tmp5523 : tmp5524;
  assign tmp5513 = ~(s2 ? tmp5514 : tmp5522);
  assign tmp5506 = s3 ? tmp5507 : tmp5513;
  assign tmp5528 = ~(l1 ? tmp5499 : tmp5511);
  assign tmp5527 = s1 ? tmp5517 : tmp5528;
  assign tmp5530 = ~(s0 ? tmp5516 : tmp5528);
  assign tmp5529 = ~(s1 ? tmp5498 : tmp5530);
  assign tmp5526 = s2 ? tmp5527 : tmp5529;
  assign tmp5532 = s0 ? tmp5520 : tmp5523;
  assign tmp5533 = ~(l1 ? tmp5499 : tmp5496);
  assign tmp5531 = s1 ? tmp5532 : tmp5533;
  assign tmp5525 = ~(s3 ? tmp5526 : tmp5531);
  assign tmp5505 = s4 ? tmp5506 : tmp5525;
  assign tmp5490 = s5 ? tmp5491 : tmp5505;
  assign tmp5543 = l1 ? 1 : tmp5503;
  assign tmp5542 = s0 ? tmp5543 : tmp5503;
  assign tmp5541 = s1 ? tmp5509 : tmp5542;
  assign tmp5545 = s0 ? tmp5493 : tmp5503;
  assign tmp5544 = s1 ? tmp5545 : tmp5501;
  assign tmp5540 = s2 ? tmp5541 : tmp5544;
  assign tmp5549 = ~(l1 ? tmp5511 : tmp5494);
  assign tmp5548 = s0 ? 1 : tmp5549;
  assign tmp5552 = l2 ? 1 : 0;
  assign tmp5551 = l1 ? tmp5552 : tmp5494;
  assign tmp5550 = ~(s0 ? tmp5551 : tmp5524);
  assign tmp5547 = ~(s1 ? tmp5548 : tmp5550);
  assign tmp5546 = ~(s2 ? tmp5514 : tmp5547);
  assign tmp5539 = s3 ? tmp5540 : tmp5546;
  assign tmp5557 = l1 ? tmp5494 : tmp5516;
  assign tmp5556 = s0 ? tmp5557 : tmp5517;
  assign tmp5559 = l1 ? tmp5518 : tmp5497;
  assign tmp5558 = s0 ? tmp5559 : tmp5528;
  assign tmp5555 = s1 ? tmp5556 : tmp5558;
  assign tmp5561 = s0 ? 1 : tmp5498;
  assign tmp5560 = ~(s1 ? tmp5561 : tmp5530);
  assign tmp5554 = s2 ? tmp5555 : tmp5560;
  assign tmp5564 = s0 ? tmp5551 : tmp5533;
  assign tmp5563 = s1 ? tmp5532 : tmp5564;
  assign tmp5566 = s0 ? tmp5557 : tmp5559;
  assign tmp5565 = s1 ? tmp5566 : 0;
  assign tmp5562 = s2 ? tmp5563 : tmp5565;
  assign tmp5553 = ~(s3 ? tmp5554 : tmp5562);
  assign tmp5538 = s4 ? tmp5539 : tmp5553;
  assign tmp5537 = s5 ? tmp5491 : tmp5538;
  assign tmp5536 = s6 ? tmp5537 : tmp5490;
  assign tmp5572 = s1 ? tmp5509 : tmp5543;
  assign tmp5571 = s2 ? tmp5572 : tmp5512;
  assign tmp5574 = s1 ? tmp5517 : tmp5521;
  assign tmp5573 = ~(s2 ? tmp5574 : tmp5522);
  assign tmp5570 = s3 ? tmp5571 : tmp5573;
  assign tmp5577 = ~(s1 ? tmp5498 : tmp5510);
  assign tmp5576 = s2 ? tmp5527 : tmp5577;
  assign tmp5578 = s1 ? tmp5523 : tmp5533;
  assign tmp5575 = ~(s3 ? tmp5576 : tmp5578);
  assign tmp5569 = s4 ? tmp5570 : tmp5575;
  assign tmp5568 = s5 ? tmp5491 : tmp5569;
  assign tmp5567 = s6 ? tmp5568 : tmp5537;
  assign tmp5535 = s7 ? tmp5536 : tmp5567;
  assign tmp5582 = s4 ? tmp5506 : tmp5575;
  assign tmp5581 = s5 ? tmp5491 : tmp5582;
  assign tmp5580 = s6 ? tmp5537 : tmp5581;
  assign tmp5586 = s3 ? tmp5571 : tmp5513;
  assign tmp5585 = s4 ? tmp5586 : tmp5575;
  assign tmp5584 = s5 ? tmp5491 : tmp5585;
  assign tmp5583 = s6 ? tmp5584 : tmp5568;
  assign tmp5579 = s7 ? tmp5580 : tmp5583;
  assign tmp5534 = s8 ? tmp5535 : tmp5579;
  assign tmp5489 = s9 ? tmp5490 : tmp5534;
  assign tmp5592 = s4 ? tmp5586 : tmp5525;
  assign tmp5591 = s5 ? tmp5491 : tmp5592;
  assign tmp5590 = s6 ? tmp5591 : tmp5568;
  assign tmp5589 = s7 ? tmp5536 : tmp5590;
  assign tmp5588 = s8 ? tmp5535 : tmp5589;
  assign tmp5587 = s9 ? tmp5490 : tmp5588;
  assign tmp5488 = s10 ? tmp5489 : tmp5587;
  assign tmp5598 = l1 ? tmp5516 : tmp5499;
  assign tmp5599 = l1 ? tmp5552 : tmp5499;
  assign tmp5597 = s1 ? tmp5598 : tmp5599;
  assign tmp5601 = s0 ? tmp5599 : tmp5516;
  assign tmp5602 = s0 ? tmp5598 : tmp5599;
  assign tmp5600 = s1 ? tmp5601 : tmp5602;
  assign tmp5596 = s2 ? tmp5597 : tmp5600;
  assign tmp5609 = ~(l2 ? 1 : tmp5497);
  assign tmp5608 = l1 ? tmp5552 : tmp5609;
  assign tmp5607 = s0 ? tmp5608 : tmp5599;
  assign tmp5610 = ~(s0 ? tmp5543 : tmp5503);
  assign tmp5606 = s1 ? tmp5607 : tmp5610;
  assign tmp5612 = s0 ? tmp5598 : tmp5516;
  assign tmp5611 = s1 ? tmp5612 : tmp5601;
  assign tmp5605 = s2 ? tmp5606 : tmp5611;
  assign tmp5615 = l1 ? tmp5494 : tmp5518;
  assign tmp5614 = s1 ? tmp5615 : tmp5521;
  assign tmp5617 = l1 ? tmp5494 : tmp5499;
  assign tmp5616 = s1 ? tmp5551 : tmp5617;
  assign tmp5613 = s2 ? tmp5614 : tmp5616;
  assign tmp5604 = s3 ? tmp5605 : tmp5613;
  assign tmp5621 = ~(l1 ? tmp5518 : tmp5511);
  assign tmp5620 = s1 ? tmp5517 : tmp5621;
  assign tmp5622 = s1 ? tmp5599 : tmp5621;
  assign tmp5619 = s2 ? tmp5620 : tmp5622;
  assign tmp5623 = s1 ? tmp5551 : tmp5599;
  assign tmp5618 = s3 ? tmp5619 : tmp5623;
  assign tmp5603 = s4 ? tmp5604 : tmp5618;
  assign tmp5595 = s5 ? tmp5596 : tmp5603;
  assign tmp5627 = ~(s5 ? tmp5596 : tmp5603);
  assign tmp5626 = s6 ? tmp5537 : tmp5627;
  assign tmp5632 = l1 ? 1 : tmp5496;
  assign tmp5633 = l1 ? tmp5518 : tmp5496;
  assign tmp5631 = s1 ? tmp5632 : tmp5633;
  assign tmp5635 = s0 ? tmp5633 : tmp5543;
  assign tmp5636 = s0 ? tmp5632 : tmp5633;
  assign tmp5634 = s1 ? tmp5635 : tmp5636;
  assign tmp5630 = s2 ? tmp5631 : tmp5634;
  assign tmp5642 = l1 ? tmp5518 : tmp5511;
  assign tmp5641 = s0 ? tmp5642 : tmp5633;
  assign tmp5640 = s1 ? tmp5641 : tmp5543;
  assign tmp5643 = s1 ? tmp5632 : tmp5635;
  assign tmp5639 = s2 ? tmp5640 : tmp5643;
  assign tmp5646 = ~(l1 ? tmp5497 : tmp5496);
  assign tmp5645 = s1 ? tmp5551 : tmp5646;
  assign tmp5644 = ~(s2 ? tmp5614 : tmp5645);
  assign tmp5638 = s3 ? tmp5639 : tmp5644;
  assign tmp5649 = ~(s1 ? tmp5633 : tmp5642);
  assign tmp5648 = s2 ? tmp5620 : tmp5649;
  assign tmp5651 = ~(l1 ? tmp5518 : tmp5496);
  assign tmp5650 = s1 ? tmp5551 : tmp5651;
  assign tmp5647 = ~(s3 ? tmp5648 : tmp5650);
  assign tmp5637 = s4 ? tmp5638 : tmp5647;
  assign tmp5629 = s5 ? tmp5630 : tmp5637;
  assign tmp5628 = s6 ? tmp5629 : tmp5537;
  assign tmp5625 = s7 ? tmp5626 : tmp5628;
  assign tmp5658 = s1 ? tmp5598 : tmp5601;
  assign tmp5657 = s2 ? tmp5606 : tmp5658;
  assign tmp5656 = s3 ? tmp5657 : tmp5613;
  assign tmp5655 = s4 ? tmp5656 : tmp5618;
  assign tmp5654 = ~(s5 ? tmp5596 : tmp5655);
  assign tmp5653 = s6 ? tmp5537 : tmp5654;
  assign tmp5660 = s5 ? tmp5596 : tmp5655;
  assign tmp5661 = ~(s5 ? tmp5630 : tmp5637);
  assign tmp5659 = ~(s6 ? tmp5660 : tmp5661);
  assign tmp5652 = s7 ? tmp5653 : tmp5659;
  assign tmp5624 = ~(s8 ? tmp5625 : tmp5652);
  assign tmp5594 = s9 ? tmp5595 : tmp5624;
  assign tmp5665 = ~(s6 ? tmp5595 : tmp5661);
  assign tmp5664 = s7 ? tmp5626 : tmp5665;
  assign tmp5663 = ~(s8 ? tmp5625 : tmp5664);
  assign tmp5662 = s9 ? tmp5595 : tmp5663;
  assign tmp5593 = ~(s10 ? tmp5594 : tmp5662);
  assign tmp5487 = s11 ? tmp5488 : tmp5593;
  assign tmp5671 = s3 ? tmp5540 : tmp5513;
  assign tmp5673 = s2 ? tmp5555 : tmp5529;
  assign tmp5674 = s2 ? tmp5531 : tmp5566;
  assign tmp5672 = ~(s3 ? tmp5673 : tmp5674);
  assign tmp5670 = s4 ? tmp5671 : tmp5672;
  assign tmp5669 = s5 ? tmp5491 : tmp5670;
  assign tmp5677 = s6 ? tmp5537 : tmp5669;
  assign tmp5676 = s7 ? tmp5677 : tmp5567;
  assign tmp5683 = s2 ? tmp5541 : tmp5512;
  assign tmp5682 = s3 ? tmp5683 : tmp5513;
  assign tmp5685 = s2 ? tmp5555 : tmp5577;
  assign tmp5684 = ~(s3 ? tmp5685 : tmp5578);
  assign tmp5681 = s4 ? tmp5682 : tmp5684;
  assign tmp5680 = s5 ? tmp5491 : tmp5681;
  assign tmp5679 = s6 ? tmp5537 : tmp5680;
  assign tmp5686 = s6 ? tmp5680 : tmp5568;
  assign tmp5678 = s7 ? tmp5679 : tmp5686;
  assign tmp5675 = s8 ? tmp5676 : tmp5678;
  assign tmp5668 = s9 ? tmp5669 : tmp5675;
  assign tmp5690 = s6 ? tmp5669 : tmp5568;
  assign tmp5689 = s7 ? tmp5677 : tmp5690;
  assign tmp5688 = s8 ? tmp5676 : tmp5689;
  assign tmp5687 = s9 ? tmp5669 : tmp5688;
  assign tmp5667 = s10 ? tmp5668 : tmp5687;
  assign tmp5698 = s0 ? tmp5551 : tmp5524;
  assign tmp5697 = s1 ? tmp5523 : tmp5698;
  assign tmp5696 = ~(s2 ? tmp5514 : tmp5697);
  assign tmp5695 = s3 ? tmp5540 : tmp5696;
  assign tmp5699 = ~(s3 ? tmp5526 : tmp5563);
  assign tmp5694 = s4 ? tmp5695 : tmp5699;
  assign tmp5693 = s5 ? tmp5491 : tmp5694;
  assign tmp5702 = s6 ? tmp5537 : tmp5693;
  assign tmp5701 = s7 ? tmp5702 : tmp5567;
  assign tmp5707 = s3 ? tmp5683 : tmp5696;
  assign tmp5706 = s4 ? tmp5707 : tmp5575;
  assign tmp5705 = s5 ? tmp5491 : tmp5706;
  assign tmp5704 = s6 ? tmp5537 : tmp5705;
  assign tmp5708 = s6 ? tmp5705 : tmp5568;
  assign tmp5703 = s7 ? tmp5704 : tmp5708;
  assign tmp5700 = s8 ? tmp5701 : tmp5703;
  assign tmp5692 = s9 ? tmp5693 : tmp5700;
  assign tmp5712 = s6 ? tmp5693 : tmp5568;
  assign tmp5711 = s7 ? tmp5702 : tmp5712;
  assign tmp5710 = s8 ? tmp5701 : tmp5711;
  assign tmp5709 = s9 ? tmp5693 : tmp5710;
  assign tmp5691 = s10 ? tmp5692 : tmp5709;
  assign tmp5666 = s11 ? tmp5667 : tmp5691;
  assign tmp5486 = s12 ? tmp5487 : tmp5666;
  assign tmp5721 = s1 ? tmp5607 : tmp5516;
  assign tmp5720 = s2 ? tmp5721 : tmp5658;
  assign tmp5719 = s3 ? tmp5720 : tmp5613;
  assign tmp5725 = s0 ? tmp5559 : tmp5621;
  assign tmp5724 = s1 ? tmp5517 : tmp5725;
  assign tmp5723 = s2 ? tmp5724 : tmp5622;
  assign tmp5726 = s2 ? tmp5623 : tmp5559;
  assign tmp5722 = s3 ? tmp5723 : tmp5726;
  assign tmp5718 = s4 ? tmp5719 : tmp5722;
  assign tmp5717 = s5 ? tmp5596 : tmp5718;
  assign tmp5730 = ~(s5 ? tmp5596 : tmp5718);
  assign tmp5729 = s6 ? tmp5537 : tmp5730;
  assign tmp5728 = s7 ? tmp5729 : tmp5628;
  assign tmp5735 = s3 ? tmp5723 : tmp5623;
  assign tmp5734 = s4 ? tmp5719 : tmp5735;
  assign tmp5733 = ~(s5 ? tmp5596 : tmp5734);
  assign tmp5732 = s6 ? tmp5537 : tmp5733;
  assign tmp5737 = s5 ? tmp5596 : tmp5734;
  assign tmp5736 = ~(s6 ? tmp5737 : tmp5661);
  assign tmp5731 = s7 ? tmp5732 : tmp5736;
  assign tmp5727 = ~(s8 ? tmp5728 : tmp5731);
  assign tmp5716 = s9 ? tmp5717 : tmp5727;
  assign tmp5741 = ~(s6 ? tmp5717 : tmp5661);
  assign tmp5740 = s7 ? tmp5729 : tmp5741;
  assign tmp5739 = ~(s8 ? tmp5728 : tmp5740);
  assign tmp5738 = s9 ? tmp5717 : tmp5739;
  assign tmp5715 = s10 ? tmp5716 : tmp5738;
  assign tmp5742 = ~(s10 ? tmp5489 : tmp5587);
  assign tmp5714 = s11 ? tmp5715 : tmp5742;
  assign tmp5752 = ~(l1 ? tmp5552 : tmp5494);
  assign tmp5751 = s0 ? 1 : tmp5752;
  assign tmp5753 = ~(l1 ? tmp5494 : tmp5499);
  assign tmp5750 = ~(s1 ? tmp5751 : tmp5753);
  assign tmp5749 = s2 ? tmp5614 : tmp5750;
  assign tmp5748 = s3 ? tmp5605 : tmp5749;
  assign tmp5756 = s1 ? tmp5559 : 0;
  assign tmp5755 = s2 ? tmp5623 : tmp5756;
  assign tmp5754 = s3 ? tmp5723 : tmp5755;
  assign tmp5747 = s4 ? tmp5748 : tmp5754;
  assign tmp5746 = s5 ? tmp5596 : tmp5747;
  assign tmp5760 = ~(s5 ? tmp5596 : tmp5747);
  assign tmp5759 = s6 ? tmp5537 : tmp5760;
  assign tmp5767 = l1 ? tmp5497 : tmp5496;
  assign tmp5766 = ~(s1 ? tmp5751 : tmp5767);
  assign tmp5765 = ~(s2 ? tmp5614 : tmp5766);
  assign tmp5764 = s3 ? tmp5639 : tmp5765;
  assign tmp5769 = s2 ? tmp5650 : 0;
  assign tmp5768 = ~(s3 ? tmp5648 : tmp5769);
  assign tmp5763 = s4 ? tmp5764 : tmp5768;
  assign tmp5762 = s5 ? tmp5630 : tmp5763;
  assign tmp5761 = s6 ? tmp5762 : tmp5537;
  assign tmp5758 = s7 ? tmp5759 : tmp5761;
  assign tmp5774 = s3 ? tmp5657 : tmp5749;
  assign tmp5773 = s4 ? tmp5774 : tmp5735;
  assign tmp5772 = ~(s5 ? tmp5596 : tmp5773);
  assign tmp5771 = s6 ? tmp5537 : tmp5772;
  assign tmp5780 = s1 ? tmp5641 : tmp5542;
  assign tmp5779 = s2 ? tmp5780 : tmp5643;
  assign tmp5778 = s3 ? tmp5779 : tmp5765;
  assign tmp5782 = s2 ? tmp5724 : tmp5649;
  assign tmp5781 = ~(s3 ? tmp5782 : tmp5650);
  assign tmp5777 = s4 ? tmp5778 : tmp5781;
  assign tmp5776 = s5 ? tmp5630 : tmp5777;
  assign tmp5784 = s4 ? tmp5764 : tmp5647;
  assign tmp5783 = s5 ? tmp5630 : tmp5784;
  assign tmp5775 = s6 ? tmp5776 : tmp5783;
  assign tmp5770 = s7 ? tmp5771 : tmp5775;
  assign tmp5757 = ~(s8 ? tmp5758 : tmp5770);
  assign tmp5745 = s9 ? tmp5746 : tmp5757;
  assign tmp5794 = s0 ? tmp5632 : tmp5503;
  assign tmp5793 = s1 ? tmp5794 : tmp5635;
  assign tmp5792 = s2 ? tmp5780 : tmp5793;
  assign tmp5791 = s3 ? tmp5792 : tmp5765;
  assign tmp5796 = s2 ? tmp5650 : tmp5756;
  assign tmp5795 = ~(s3 ? tmp5782 : tmp5796);
  assign tmp5790 = s4 ? tmp5791 : tmp5795;
  assign tmp5789 = s5 ? tmp5630 : tmp5790;
  assign tmp5788 = s6 ? tmp5789 : tmp5762;
  assign tmp5787 = s7 ? tmp5759 : tmp5788;
  assign tmp5786 = ~(s8 ? tmp5758 : tmp5787);
  assign tmp5785 = s9 ? tmp5746 : tmp5786;
  assign tmp5744 = s10 ? tmp5745 : tmp5785;
  assign tmp5803 = s1 ? tmp5517 : tmp5558;
  assign tmp5802 = s2 ? tmp5803 : tmp5560;
  assign tmp5804 = s2 ? tmp5531 : tmp5756;
  assign tmp5801 = ~(s3 ? tmp5802 : tmp5804);
  assign tmp5800 = s4 ? tmp5506 : tmp5801;
  assign tmp5799 = s5 ? tmp5491 : tmp5800;
  assign tmp5807 = s6 ? tmp5537 : tmp5799;
  assign tmp5806 = s7 ? tmp5807 : tmp5567;
  assign tmp5814 = ~(s1 ? tmp5561 : tmp5510);
  assign tmp5813 = s2 ? tmp5803 : tmp5814;
  assign tmp5812 = ~(s3 ? tmp5813 : tmp5578);
  assign tmp5811 = s4 ? tmp5506 : tmp5812;
  assign tmp5810 = s5 ? tmp5491 : tmp5811;
  assign tmp5809 = s6 ? tmp5537 : tmp5810;
  assign tmp5817 = s4 ? tmp5586 : tmp5812;
  assign tmp5816 = s5 ? tmp5491 : tmp5817;
  assign tmp5815 = s6 ? tmp5816 : tmp5568;
  assign tmp5808 = s7 ? tmp5809 : tmp5815;
  assign tmp5805 = s8 ? tmp5806 : tmp5808;
  assign tmp5798 = s9 ? tmp5799 : tmp5805;
  assign tmp5823 = s4 ? tmp5586 : tmp5801;
  assign tmp5822 = s5 ? tmp5491 : tmp5823;
  assign tmp5821 = s6 ? tmp5822 : tmp5568;
  assign tmp5820 = s7 ? tmp5807 : tmp5821;
  assign tmp5819 = s8 ? tmp5806 : tmp5820;
  assign tmp5818 = s9 ? tmp5799 : tmp5819;
  assign tmp5797 = ~(s10 ? tmp5798 : tmp5818);
  assign tmp5743 = s11 ? tmp5744 : tmp5797;
  assign tmp5713 = ~(s12 ? tmp5714 : tmp5743);
  assign tmp5485 = s13 ? tmp5486 : tmp5713;
  assign tmp5831 = s4 ? tmp5719 : tmp5618;
  assign tmp5830 = s5 ? tmp5596 : tmp5831;
  assign tmp5833 = s7 ? tmp5536 : tmp5628;
  assign tmp5839 = s2 ? tmp5721 : tmp5611;
  assign tmp5842 = s0 ? tmp5516 : tmp5615;
  assign tmp5841 = s1 ? tmp5842 : tmp5519;
  assign tmp5844 = ~(s0 ? tmp5551 : tmp5617);
  assign tmp5843 = ~(s1 ? tmp5751 : tmp5844);
  assign tmp5840 = s2 ? tmp5841 : tmp5843;
  assign tmp5838 = s3 ? tmp5839 : tmp5840;
  assign tmp5847 = s1 ? tmp5556 : tmp5725;
  assign tmp5850 = ~(l1 ? tmp5552 : tmp5499);
  assign tmp5849 = s0 ? 1 : tmp5850;
  assign tmp5851 = ~(s0 ? tmp5516 : tmp5621);
  assign tmp5848 = ~(s1 ? tmp5849 : tmp5851);
  assign tmp5846 = s2 ? tmp5847 : tmp5848;
  assign tmp5854 = s0 ? tmp5520 : tmp5551;
  assign tmp5855 = s0 ? tmp5551 : tmp5599;
  assign tmp5853 = s1 ? tmp5854 : tmp5855;
  assign tmp5852 = s2 ? tmp5853 : tmp5565;
  assign tmp5845 = s3 ? tmp5846 : tmp5852;
  assign tmp5837 = s4 ? tmp5838 : tmp5845;
  assign tmp5836 = s5 ? tmp5596 : tmp5837;
  assign tmp5835 = s6 ? tmp5836 : tmp5830;
  assign tmp5856 = ~(s6 ? tmp5581 : tmp5629);
  assign tmp5834 = ~(s7 ? tmp5835 : tmp5856);
  assign tmp5832 = ~(s8 ? tmp5833 : tmp5834);
  assign tmp5829 = s9 ? tmp5830 : tmp5832;
  assign tmp5860 = ~(s6 ? tmp5490 : tmp5629);
  assign tmp5859 = ~(s7 ? tmp5835 : tmp5860);
  assign tmp5858 = ~(s8 ? tmp5833 : tmp5859);
  assign tmp5857 = s9 ? tmp5830 : tmp5858;
  assign tmp5828 = s10 ? tmp5829 : tmp5857;
  assign tmp5865 = s6 ? tmp5660 : tmp5661;
  assign tmp5864 = ~(s7 ? tmp5835 : tmp5865);
  assign tmp5863 = ~(s8 ? tmp5625 : tmp5864);
  assign tmp5862 = s9 ? tmp5830 : tmp5863;
  assign tmp5869 = s6 ? tmp5595 : tmp5661;
  assign tmp5868 = ~(s7 ? tmp5835 : tmp5869);
  assign tmp5867 = ~(s8 ? tmp5625 : tmp5868);
  assign tmp5866 = s9 ? tmp5830 : tmp5867;
  assign tmp5861 = s10 ? tmp5862 : tmp5866;
  assign tmp5827 = s11 ? tmp5828 : tmp5861;
  assign tmp5874 = s7 ? tmp5677 : tmp5628;
  assign tmp5876 = ~(s6 ? tmp5680 : tmp5629);
  assign tmp5875 = ~(s7 ? tmp5835 : tmp5876);
  assign tmp5873 = ~(s8 ? tmp5874 : tmp5875);
  assign tmp5872 = s9 ? tmp5830 : tmp5873;
  assign tmp5880 = ~(s6 ? tmp5669 : tmp5629);
  assign tmp5879 = ~(s7 ? tmp5835 : tmp5880);
  assign tmp5878 = ~(s8 ? tmp5874 : tmp5879);
  assign tmp5877 = s9 ? tmp5830 : tmp5878;
  assign tmp5871 = s10 ? tmp5872 : tmp5877;
  assign tmp5884 = s7 ? tmp5702 : tmp5628;
  assign tmp5887 = ~(s5 ? tmp5596 : tmp5831);
  assign tmp5886 = s6 ? tmp5537 : tmp5887;
  assign tmp5888 = s6 ? tmp5705 : tmp5629;
  assign tmp5885 = s7 ? tmp5886 : tmp5888;
  assign tmp5883 = ~(s8 ? tmp5884 : tmp5885);
  assign tmp5882 = s9 ? tmp5830 : tmp5883;
  assign tmp5892 = s6 ? tmp5693 : tmp5629;
  assign tmp5891 = s7 ? tmp5886 : tmp5892;
  assign tmp5890 = ~(s8 ? tmp5884 : tmp5891);
  assign tmp5889 = s9 ? tmp5830 : tmp5890;
  assign tmp5881 = s10 ? tmp5882 : tmp5889;
  assign tmp5870 = s11 ? tmp5871 : tmp5881;
  assign tmp5826 = s12 ? tmp5827 : tmp5870;
  assign tmp5899 = s6 ? tmp5737 : tmp5661;
  assign tmp5898 = ~(s7 ? tmp5835 : tmp5899);
  assign tmp5897 = ~(s8 ? tmp5728 : tmp5898);
  assign tmp5896 = s9 ? tmp5830 : tmp5897;
  assign tmp5903 = s6 ? tmp5717 : tmp5661;
  assign tmp5902 = ~(s7 ? tmp5835 : tmp5903);
  assign tmp5901 = ~(s8 ? tmp5728 : tmp5902);
  assign tmp5900 = s9 ? tmp5830 : tmp5901;
  assign tmp5895 = s10 ? tmp5896 : tmp5900;
  assign tmp5894 = s11 ? tmp5895 : tmp5828;
  assign tmp5908 = s7 ? tmp5759 : tmp5628;
  assign tmp5911 = s5 ? tmp5596 : tmp5773;
  assign tmp5910 = ~(s6 ? tmp5911 : tmp5661);
  assign tmp5909 = s7 ? tmp5886 : tmp5910;
  assign tmp5907 = ~(s8 ? tmp5908 : tmp5909);
  assign tmp5906 = s9 ? tmp5830 : tmp5907;
  assign tmp5915 = ~(s6 ? tmp5746 : tmp5661);
  assign tmp5914 = s7 ? tmp5886 : tmp5915;
  assign tmp5913 = ~(s8 ? tmp5908 : tmp5914);
  assign tmp5912 = s9 ? tmp5830 : tmp5913;
  assign tmp5905 = s10 ? tmp5906 : tmp5912;
  assign tmp5919 = s7 ? tmp5807 : tmp5628;
  assign tmp5921 = s6 ? tmp5810 : tmp5629;
  assign tmp5920 = s7 ? tmp5886 : tmp5921;
  assign tmp5918 = ~(s8 ? tmp5919 : tmp5920);
  assign tmp5917 = s9 ? tmp5830 : tmp5918;
  assign tmp5925 = s6 ? tmp5799 : tmp5629;
  assign tmp5924 = s7 ? tmp5886 : tmp5925;
  assign tmp5923 = ~(s8 ? tmp5919 : tmp5924);
  assign tmp5922 = s9 ? tmp5830 : tmp5923;
  assign tmp5916 = s10 ? tmp5917 : tmp5922;
  assign tmp5904 = s11 ? tmp5905 : tmp5916;
  assign tmp5893 = s12 ? tmp5894 : tmp5904;
  assign tmp5825 = s13 ? tmp5826 : tmp5893;
  assign tmp5938 = s1 ? tmp5515 : tmp5521;
  assign tmp5937 = ~(s2 ? tmp5938 : tmp5522);
  assign tmp5936 = s3 ? tmp5571 : tmp5937;
  assign tmp5939 = ~(s3 ? tmp5526 : tmp5578);
  assign tmp5935 = s4 ? tmp5936 : tmp5939;
  assign tmp5934 = s5 ? tmp5491 : tmp5935;
  assign tmp5933 = s6 ? tmp5934 : tmp5537;
  assign tmp5932 = s7 ? tmp5536 : tmp5933;
  assign tmp5943 = s4 ? tmp5936 : tmp5575;
  assign tmp5942 = s5 ? tmp5491 : tmp5943;
  assign tmp5941 = s6 ? tmp5584 : tmp5942;
  assign tmp5940 = s7 ? tmp5580 : tmp5941;
  assign tmp5931 = s8 ? tmp5932 : tmp5940;
  assign tmp5930 = s9 ? tmp5490 : tmp5931;
  assign tmp5947 = s6 ? tmp5591 : tmp5934;
  assign tmp5946 = s7 ? tmp5536 : tmp5947;
  assign tmp5945 = s8 ? tmp5932 : tmp5946;
  assign tmp5944 = s9 ? tmp5490 : tmp5945;
  assign tmp5929 = s10 ? tmp5930 : tmp5944;
  assign tmp5955 = s3 ? tmp5792 : tmp5644;
  assign tmp5954 = s4 ? tmp5955 : tmp5647;
  assign tmp5953 = s5 ? tmp5630 : tmp5954;
  assign tmp5952 = s6 ? tmp5953 : tmp5537;
  assign tmp5951 = s7 ? tmp5626 : tmp5952;
  assign tmp5960 = s3 ? tmp5779 : tmp5644;
  assign tmp5959 = s4 ? tmp5960 : tmp5647;
  assign tmp5958 = ~(s5 ? tmp5630 : tmp5959);
  assign tmp5957 = ~(s6 ? tmp5660 : tmp5958);
  assign tmp5956 = s7 ? tmp5653 : tmp5957;
  assign tmp5950 = ~(s8 ? tmp5951 : tmp5956);
  assign tmp5949 = s9 ? tmp5595 : tmp5950;
  assign tmp5965 = ~(s5 ? tmp5630 : tmp5954);
  assign tmp5964 = ~(s6 ? tmp5595 : tmp5965);
  assign tmp5963 = s7 ? tmp5626 : tmp5964;
  assign tmp5962 = ~(s8 ? tmp5951 : tmp5963);
  assign tmp5961 = s9 ? tmp5595 : tmp5962;
  assign tmp5948 = ~(s10 ? tmp5949 : tmp5961);
  assign tmp5928 = s11 ? tmp5929 : tmp5948;
  assign tmp5976 = s1 ? tmp5556 : tmp5528;
  assign tmp5975 = s2 ? tmp5976 : tmp5577;
  assign tmp5977 = s2 ? tmp5578 : tmp5557;
  assign tmp5974 = ~(s3 ? tmp5975 : tmp5977);
  assign tmp5973 = s4 ? tmp5570 : tmp5974;
  assign tmp5972 = s5 ? tmp5491 : tmp5973;
  assign tmp5971 = s6 ? tmp5972 : tmp5537;
  assign tmp5970 = s7 ? tmp5677 : tmp5971;
  assign tmp5982 = ~(s3 ? tmp5975 : tmp5578);
  assign tmp5981 = s4 ? tmp5570 : tmp5982;
  assign tmp5980 = s5 ? tmp5491 : tmp5981;
  assign tmp5979 = s6 ? tmp5680 : tmp5980;
  assign tmp5978 = s7 ? tmp5679 : tmp5979;
  assign tmp5969 = s8 ? tmp5970 : tmp5978;
  assign tmp5968 = s9 ? tmp5669 : tmp5969;
  assign tmp5986 = s6 ? tmp5669 : tmp5972;
  assign tmp5985 = s7 ? tmp5677 : tmp5986;
  assign tmp5984 = s8 ? tmp5970 : tmp5985;
  assign tmp5983 = s9 ? tmp5669 : tmp5984;
  assign tmp5967 = s10 ? tmp5968 : tmp5983;
  assign tmp5995 = ~(s2 ? tmp5574 : tmp5697);
  assign tmp5994 = s3 ? tmp5571 : tmp5995;
  assign tmp5997 = s1 ? tmp5523 : tmp5564;
  assign tmp5996 = ~(s3 ? tmp5576 : tmp5997);
  assign tmp5993 = s4 ? tmp5994 : tmp5996;
  assign tmp5992 = s5 ? tmp5491 : tmp5993;
  assign tmp5991 = s6 ? tmp5992 : tmp5537;
  assign tmp5990 = s7 ? tmp5702 : tmp5991;
  assign tmp6001 = s4 ? tmp5994 : tmp5575;
  assign tmp6000 = s5 ? tmp5491 : tmp6001;
  assign tmp5999 = s6 ? tmp5705 : tmp6000;
  assign tmp5998 = s7 ? tmp5704 : tmp5999;
  assign tmp5989 = s8 ? tmp5990 : tmp5998;
  assign tmp5988 = s9 ? tmp5693 : tmp5989;
  assign tmp6005 = s6 ? tmp5693 : tmp5992;
  assign tmp6004 = s7 ? tmp5702 : tmp6005;
  assign tmp6003 = s8 ? tmp5990 : tmp6004;
  assign tmp6002 = s9 ? tmp5693 : tmp6003;
  assign tmp5987 = s10 ? tmp5988 : tmp6002;
  assign tmp5966 = s11 ? tmp5967 : tmp5987;
  assign tmp5927 = s12 ? tmp5928 : tmp5966;
  assign tmp6016 = s2 ? tmp5650 : tmp5559;
  assign tmp6015 = ~(s3 ? tmp5782 : tmp6016);
  assign tmp6014 = s4 ? tmp5638 : tmp6015;
  assign tmp6013 = s5 ? tmp5630 : tmp6014;
  assign tmp6012 = s6 ? tmp6013 : tmp5537;
  assign tmp6011 = s7 ? tmp5729 : tmp6012;
  assign tmp6020 = s4 ? tmp5638 : tmp5781;
  assign tmp6019 = ~(s5 ? tmp5630 : tmp6020);
  assign tmp6018 = ~(s6 ? tmp5737 : tmp6019);
  assign tmp6017 = s7 ? tmp5732 : tmp6018;
  assign tmp6010 = ~(s8 ? tmp6011 : tmp6017);
  assign tmp6009 = s9 ? tmp5717 : tmp6010;
  assign tmp6025 = ~(s5 ? tmp5630 : tmp6014);
  assign tmp6024 = ~(s6 ? tmp5717 : tmp6025);
  assign tmp6023 = s7 ? tmp5729 : tmp6024;
  assign tmp6022 = ~(s8 ? tmp6011 : tmp6023);
  assign tmp6021 = s9 ? tmp5717 : tmp6022;
  assign tmp6008 = s10 ? tmp6009 : tmp6021;
  assign tmp6035 = s1 ? tmp5517 : tmp5519;
  assign tmp6034 = ~(s2 ? tmp6035 : tmp5522);
  assign tmp6033 = s3 ? tmp5571 : tmp6034;
  assign tmp6036 = ~(s3 ? tmp5576 : tmp5531);
  assign tmp6032 = s4 ? tmp6033 : tmp6036;
  assign tmp6031 = s5 ? tmp5491 : tmp6032;
  assign tmp6030 = s6 ? tmp6031 : tmp5537;
  assign tmp6029 = s7 ? tmp5536 : tmp6030;
  assign tmp6040 = s4 ? tmp6033 : tmp5575;
  assign tmp6039 = s5 ? tmp5491 : tmp6040;
  assign tmp6038 = s6 ? tmp5584 : tmp6039;
  assign tmp6037 = s7 ? tmp5580 : tmp6038;
  assign tmp6028 = s8 ? tmp6029 : tmp6037;
  assign tmp6027 = s9 ? tmp5490 : tmp6028;
  assign tmp6044 = s6 ? tmp5591 : tmp6031;
  assign tmp6043 = s7 ? tmp5536 : tmp6044;
  assign tmp6042 = s8 ? tmp6029 : tmp6043;
  assign tmp6041 = s9 ? tmp5490 : tmp6042;
  assign tmp6026 = ~(s10 ? tmp6027 : tmp6041);
  assign tmp6007 = s11 ? tmp6008 : tmp6026;
  assign tmp6054 = s2 ? tmp5527 : tmp5814;
  assign tmp6055 = s2 ? tmp5578 : 0;
  assign tmp6053 = ~(s3 ? tmp6054 : tmp6055);
  assign tmp6052 = s4 ? tmp5570 : tmp6053;
  assign tmp6051 = s5 ? tmp5491 : tmp6052;
  assign tmp6050 = s6 ? tmp6051 : tmp5537;
  assign tmp6049 = s7 ? tmp5807 : tmp6050;
  assign tmp6060 = ~(s3 ? tmp6054 : tmp5578);
  assign tmp6059 = s4 ? tmp5570 : tmp6060;
  assign tmp6058 = s5 ? tmp5491 : tmp6059;
  assign tmp6057 = s6 ? tmp5816 : tmp6058;
  assign tmp6056 = s7 ? tmp5809 : tmp6057;
  assign tmp6048 = s8 ? tmp6049 : tmp6056;
  assign tmp6047 = s9 ? tmp5799 : tmp6048;
  assign tmp6064 = s6 ? tmp5822 : tmp6051;
  assign tmp6063 = s7 ? tmp5807 : tmp6064;
  assign tmp6062 = s8 ? tmp6049 : tmp6063;
  assign tmp6061 = s9 ? tmp5799 : tmp6062;
  assign tmp6046 = ~(s10 ? tmp6047 : tmp6061);
  assign tmp6045 = s11 ? tmp5744 : tmp6046;
  assign tmp6006 = ~(s12 ? tmp6007 : tmp6045);
  assign tmp5926 = ~(s13 ? tmp5927 : tmp6006);
  assign tmp5824 = ~(s15 ? tmp5825 : tmp5926);
  assign tmp5484 = ~(s16 ? tmp5485 : tmp5824);
  assign s3n = tmp5484;

  assign tmp6076 = l3 ? 1 : 0;
  assign tmp6075 = l2 ? tmp6076 : 1;
  assign tmp6078 = ~(l3 ? 1 : 0);
  assign tmp6077 = l2 ? 1 : tmp6078;
  assign tmp6074 = l1 ? tmp6075 : tmp6077;
  assign tmp6079 = l1 ? 1 : tmp6077;
  assign tmp6073 = s1 ? tmp6074 : tmp6079;
  assign tmp6082 = l1 ? 1 : tmp6078;
  assign tmp6081 = s0 ? tmp6079 : tmp6082;
  assign tmp6080 = s1 ? tmp6079 : tmp6081;
  assign tmp6072 = s2 ? tmp6073 : tmp6080;
  assign tmp6088 = ~(l2 ? tmp6076 : 0);
  assign tmp6087 = ~(l1 ? 1 : tmp6088);
  assign tmp6086 = s1 ? tmp6079 : tmp6087;
  assign tmp6092 = l2 ? tmp6076 : 0;
  assign tmp6091 = l1 ? tmp6076 : tmp6092;
  assign tmp6090 = s0 ? tmp6079 : tmp6091;
  assign tmp6089 = s1 ? tmp6074 : tmp6090;
  assign tmp6085 = s2 ? tmp6086 : tmp6089;
  assign tmp6095 = s0 ? 1 : 0;
  assign tmp6098 = l2 ? tmp6076 : tmp6078;
  assign tmp6097 = l1 ? tmp6098 : 1;
  assign tmp6096 = ~(s0 ? tmp6097 : tmp6079);
  assign tmp6094 = s1 ? tmp6095 : tmp6096;
  assign tmp6101 = l2 ? 1 : 0;
  assign tmp6100 = l1 ? tmp6101 : tmp6088;
  assign tmp6102 = ~(l1 ? tmp6076 : tmp6078);
  assign tmp6099 = s1 ? tmp6100 : tmp6102;
  assign tmp6093 = ~(s2 ? tmp6094 : tmp6099);
  assign tmp6084 = s3 ? tmp6085 : tmp6093;
  assign tmp6106 = l1 ? tmp6075 : tmp6076;
  assign tmp6105 = s1 ? tmp6106 : 0;
  assign tmp6109 = l1 ? tmp6092 : tmp6076;
  assign tmp6108 = ~(s0 ? 1 : tmp6109);
  assign tmp6107 = ~(s1 ? tmp6079 : tmp6108);
  assign tmp6104 = s2 ? tmp6105 : tmp6107;
  assign tmp6111 = s0 ? tmp6097 : tmp6079;
  assign tmp6110 = ~(s1 ? tmp6111 : tmp6082);
  assign tmp6103 = ~(s3 ? tmp6104 : tmp6110);
  assign tmp6083 = s4 ? tmp6084 : tmp6103;
  assign tmp6071 = s5 ? tmp6072 : tmp6083;
  assign tmp6118 = l1 ? tmp6076 : tmp6101;
  assign tmp6120 = l2 ? 1 : tmp6076;
  assign tmp6119 = l1 ? tmp6120 : tmp6101;
  assign tmp6117 = s1 ? tmp6118 : tmp6119;
  assign tmp6123 = l1 ? tmp6120 : tmp6077;
  assign tmp6122 = s0 ? tmp6119 : tmp6123;
  assign tmp6125 = l1 ? 1 : tmp6101;
  assign tmp6127 = ~(l2 ? tmp6076 : 1);
  assign tmp6126 = l1 ? tmp6120 : tmp6127;
  assign tmp6124 = s0 ? tmp6125 : tmp6126;
  assign tmp6121 = s1 ? tmp6122 : tmp6124;
  assign tmp6116 = s2 ? tmp6117 : tmp6121;
  assign tmp6132 = s0 ? tmp6125 : tmp6119;
  assign tmp6134 = ~(l1 ? 1 : tmp6077);
  assign tmp6133 = s0 ? tmp6092 : tmp6134;
  assign tmp6131 = s1 ? tmp6132 : tmp6133;
  assign tmp6136 = s0 ? tmp6118 : tmp6134;
  assign tmp6137 = s0 ? tmp6119 : tmp6091;
  assign tmp6135 = s1 ? tmp6136 : tmp6137;
  assign tmp6130 = s2 ? tmp6131 : tmp6135;
  assign tmp6140 = ~(s0 ? tmp6097 : tmp6119);
  assign tmp6139 = s1 ? tmp6095 : tmp6140;
  assign tmp6143 = ~(l1 ? tmp6077 : tmp6088);
  assign tmp6142 = s0 ? tmp6120 : tmp6143;
  assign tmp6145 = ~(l1 ? tmp6076 : tmp6127);
  assign tmp6144 = ~(s0 ? tmp6079 : tmp6145);
  assign tmp6141 = ~(s1 ? tmp6142 : tmp6144);
  assign tmp6138 = ~(s2 ? tmp6139 : tmp6141);
  assign tmp6129 = s3 ? tmp6130 : tmp6138;
  assign tmp6150 = l1 ? 1 : tmp6098;
  assign tmp6149 = s0 ? tmp6150 : tmp6075;
  assign tmp6152 = l1 ? 1 : tmp6075;
  assign tmp6153 = ~(l2 ? 1 : tmp6076);
  assign tmp6151 = s0 ? tmp6152 : tmp6153;
  assign tmp6148 = s1 ? tmp6149 : tmp6151;
  assign tmp6156 = l1 ? tmp6092 : tmp6120;
  assign tmp6155 = s0 ? tmp6156 : tmp6119;
  assign tmp6158 = l1 ? tmp6098 : tmp6075;
  assign tmp6157 = ~(s0 ? 1 : tmp6158);
  assign tmp6154 = ~(s1 ? tmp6155 : tmp6157);
  assign tmp6147 = s2 ? tmp6148 : tmp6154;
  assign tmp6161 = s0 ? tmp6097 : tmp6119;
  assign tmp6163 = ~(l1 ? tmp6120 : tmp6127);
  assign tmp6162 = ~(s0 ? tmp6079 : tmp6163);
  assign tmp6160 = s1 ? tmp6161 : tmp6162;
  assign tmp6165 = s0 ? tmp6150 : tmp6152;
  assign tmp6166 = ~(s0 ? tmp6120 : tmp6156);
  assign tmp6164 = ~(s1 ? tmp6165 : tmp6166);
  assign tmp6159 = ~(s2 ? tmp6160 : tmp6164);
  assign tmp6146 = ~(s3 ? tmp6147 : tmp6159);
  assign tmp6128 = s4 ? tmp6129 : tmp6146;
  assign tmp6115 = s5 ? tmp6116 : tmp6128;
  assign tmp6114 = s6 ? tmp6115 : tmp6071;
  assign tmp6172 = s1 ? tmp6079 : tmp6092;
  assign tmp6171 = s2 ? tmp6172 : tmp6089;
  assign tmp6174 = s1 ? 1 : tmp6079;
  assign tmp6175 = ~(s1 ? tmp6100 : tmp6102);
  assign tmp6173 = s2 ? tmp6174 : tmp6175;
  assign tmp6170 = s3 ? tmp6171 : tmp6173;
  assign tmp6179 = ~(l1 ? tmp6092 : tmp6076);
  assign tmp6178 = ~(s1 ? tmp6079 : tmp6179);
  assign tmp6177 = s2 ? tmp6105 : tmp6178;
  assign tmp6180 = ~(s1 ? tmp6079 : tmp6082);
  assign tmp6176 = ~(s3 ? tmp6177 : tmp6180);
  assign tmp6169 = s4 ? tmp6170 : tmp6176;
  assign tmp6168 = s5 ? tmp6072 : tmp6169;
  assign tmp6167 = s6 ? tmp6168 : tmp6115;
  assign tmp6113 = s7 ? tmp6114 : tmp6167;
  assign tmp6184 = s4 ? tmp6084 : tmp6176;
  assign tmp6183 = s5 ? tmp6072 : tmp6184;
  assign tmp6182 = s6 ? tmp6115 : tmp6183;
  assign tmp6188 = s3 ? tmp6171 : tmp6093;
  assign tmp6187 = s4 ? tmp6188 : tmp6176;
  assign tmp6186 = s5 ? tmp6072 : tmp6187;
  assign tmp6185 = s6 ? tmp6186 : tmp6168;
  assign tmp6181 = s7 ? tmp6182 : tmp6185;
  assign tmp6112 = s8 ? tmp6113 : tmp6181;
  assign tmp6070 = s9 ? tmp6071 : tmp6112;
  assign tmp6194 = s4 ? tmp6188 : tmp6103;
  assign tmp6193 = s5 ? tmp6072 : tmp6194;
  assign tmp6192 = s6 ? tmp6193 : tmp6168;
  assign tmp6191 = s7 ? tmp6114 : tmp6192;
  assign tmp6190 = s8 ? tmp6113 : tmp6191;
  assign tmp6189 = s9 ? tmp6071 : tmp6190;
  assign tmp6069 = s10 ? tmp6070 : tmp6189;
  assign tmp6201 = ~(l2 ? 1 : tmp6078);
  assign tmp6200 = l1 ? tmp6120 : tmp6201;
  assign tmp6202 = l1 ? tmp6076 : tmp6201;
  assign tmp6199 = s1 ? tmp6200 : tmp6202;
  assign tmp6204 = s0 ? tmp6202 : tmp6076;
  assign tmp6203 = s1 ? tmp6202 : tmp6204;
  assign tmp6198 = s2 ? tmp6199 : tmp6203;
  assign tmp6209 = ~(s0 ? tmp6092 : tmp6134);
  assign tmp6208 = s1 ? tmp6202 : tmp6209;
  assign tmp6211 = s0 ? tmp6200 : tmp6079;
  assign tmp6213 = l1 ? 1 : tmp6088;
  assign tmp6212 = s0 ? tmp6202 : tmp6213;
  assign tmp6210 = s1 ? tmp6211 : tmp6212;
  assign tmp6207 = s2 ? tmp6208 : tmp6210;
  assign tmp6216 = l1 ? tmp6077 : 1;
  assign tmp6215 = s1 ? tmp6216 : tmp6079;
  assign tmp6218 = l1 ? tmp6120 : tmp6088;
  assign tmp6219 = l1 ? 1 : tmp6076;
  assign tmp6217 = ~(s1 ? tmp6218 : tmp6219);
  assign tmp6214 = ~(s2 ? tmp6215 : tmp6217);
  assign tmp6206 = s3 ? tmp6207 : tmp6214;
  assign tmp6223 = ~(l1 ? tmp6077 : 1);
  assign tmp6222 = s1 ? tmp6106 : tmp6223;
  assign tmp6224 = s1 ? tmp6202 : tmp6076;
  assign tmp6221 = s2 ? tmp6222 : tmp6224;
  assign tmp6225 = ~(s1 ? tmp6077 : tmp6078);
  assign tmp6220 = s3 ? tmp6221 : tmp6225;
  assign tmp6205 = s4 ? tmp6206 : tmp6220;
  assign tmp6197 = s5 ? tmp6198 : tmp6205;
  assign tmp6229 = ~(s5 ? tmp6198 : tmp6205);
  assign tmp6228 = s6 ? tmp6115 : tmp6229;
  assign tmp6234 = l1 ? tmp6098 : tmp6077;
  assign tmp6233 = s1 ? tmp6234 : tmp6077;
  assign tmp6237 = l1 ? tmp6077 : tmp6078;
  assign tmp6236 = s0 ? tmp6077 : tmp6237;
  assign tmp6235 = s1 ? tmp6077 : tmp6236;
  assign tmp6232 = s2 ? tmp6233 : tmp6235;
  assign tmp6241 = s1 ? tmp6077 : tmp6092;
  assign tmp6243 = s0 ? tmp6077 : tmp6092;
  assign tmp6242 = s1 ? tmp6234 : tmp6243;
  assign tmp6240 = s2 ? tmp6241 : tmp6242;
  assign tmp6246 = ~(l1 ? tmp6092 : tmp6078);
  assign tmp6245 = ~(s1 ? tmp6218 : tmp6246);
  assign tmp6244 = s2 ? tmp6215 : tmp6245;
  assign tmp6239 = s3 ? tmp6240 : tmp6244;
  assign tmp6248 = s2 ? tmp6222 : tmp6225;
  assign tmp6249 = ~(s1 ? tmp6077 : tmp6237);
  assign tmp6247 = ~(s3 ? tmp6248 : tmp6249);
  assign tmp6238 = s4 ? tmp6239 : tmp6247;
  assign tmp6231 = s5 ? tmp6232 : tmp6238;
  assign tmp6230 = s6 ? tmp6231 : tmp6115;
  assign tmp6227 = s7 ? tmp6228 : tmp6230;
  assign tmp6256 = s1 ? tmp6200 : tmp6212;
  assign tmp6255 = s2 ? tmp6208 : tmp6256;
  assign tmp6254 = s3 ? tmp6255 : tmp6214;
  assign tmp6253 = s4 ? tmp6254 : tmp6220;
  assign tmp6252 = ~(s5 ? tmp6198 : tmp6253);
  assign tmp6251 = s6 ? tmp6115 : tmp6252;
  assign tmp6258 = s5 ? tmp6198 : tmp6253;
  assign tmp6259 = ~(s5 ? tmp6232 : tmp6238);
  assign tmp6257 = ~(s6 ? tmp6258 : tmp6259);
  assign tmp6250 = s7 ? tmp6251 : tmp6257;
  assign tmp6226 = ~(s8 ? tmp6227 : tmp6250);
  assign tmp6196 = s9 ? tmp6197 : tmp6226;
  assign tmp6263 = ~(s6 ? tmp6197 : tmp6259);
  assign tmp6262 = s7 ? tmp6228 : tmp6263;
  assign tmp6261 = ~(s8 ? tmp6227 : tmp6262);
  assign tmp6260 = s9 ? tmp6197 : tmp6261;
  assign tmp6195 = ~(s10 ? tmp6196 : tmp6260);
  assign tmp6068 = s11 ? tmp6069 : tmp6195;
  assign tmp6270 = l1 ? tmp6075 : tmp6101;
  assign tmp6269 = s1 ? tmp6270 : tmp6125;
  assign tmp6272 = s0 ? tmp6125 : tmp6079;
  assign tmp6274 = l1 ? 1 : tmp6127;
  assign tmp6273 = s0 ? tmp6125 : tmp6274;
  assign tmp6271 = s1 ? tmp6272 : tmp6273;
  assign tmp6268 = s2 ? tmp6269 : tmp6271;
  assign tmp6278 = s1 ? tmp6125 : tmp6133;
  assign tmp6280 = s0 ? tmp6270 : tmp6134;
  assign tmp6281 = s0 ? tmp6125 : tmp6091;
  assign tmp6279 = s1 ? tmp6280 : tmp6281;
  assign tmp6277 = s2 ? tmp6278 : tmp6279;
  assign tmp6284 = ~(s0 ? tmp6097 : tmp6125);
  assign tmp6283 = s1 ? tmp6095 : tmp6284;
  assign tmp6285 = s1 ? tmp6100 : tmp6145;
  assign tmp6282 = ~(s2 ? tmp6283 : tmp6285);
  assign tmp6276 = s3 ? tmp6277 : tmp6282;
  assign tmp6290 = ~(l1 ? 1 : tmp6120);
  assign tmp6289 = s0 ? tmp6152 : tmp6290;
  assign tmp6288 = s1 ? tmp6149 : tmp6289;
  assign tmp6293 = l1 ? tmp6092 : tmp6075;
  assign tmp6292 = ~(s0 ? 1 : tmp6293);
  assign tmp6291 = ~(s1 ? tmp6125 : tmp6292);
  assign tmp6287 = s2 ? tmp6288 : tmp6291;
  assign tmp6296 = s0 ? tmp6097 : tmp6125;
  assign tmp6295 = s1 ? tmp6296 : tmp6274;
  assign tmp6297 = ~(s0 ? tmp6150 : tmp6152);
  assign tmp6294 = ~(s2 ? tmp6295 : tmp6297);
  assign tmp6286 = ~(s3 ? tmp6287 : tmp6294);
  assign tmp6275 = s4 ? tmp6276 : tmp6286;
  assign tmp6267 = s5 ? tmp6268 : tmp6275;
  assign tmp6300 = s6 ? tmp6115 : tmp6267;
  assign tmp6306 = s1 ? tmp6125 : tmp6092;
  assign tmp6307 = s1 ? tmp6270 : tmp6281;
  assign tmp6305 = s2 ? tmp6306 : tmp6307;
  assign tmp6309 = s1 ? 1 : tmp6125;
  assign tmp6310 = ~(s1 ? tmp6100 : tmp6145);
  assign tmp6308 = s2 ? tmp6309 : tmp6310;
  assign tmp6304 = s3 ? tmp6305 : tmp6308;
  assign tmp6313 = s1 ? tmp6075 : tmp6290;
  assign tmp6315 = ~(l1 ? tmp6092 : tmp6075);
  assign tmp6314 = ~(s1 ? tmp6125 : tmp6315);
  assign tmp6312 = s2 ? tmp6313 : tmp6314;
  assign tmp6316 = ~(s1 ? tmp6125 : tmp6274);
  assign tmp6311 = ~(s3 ? tmp6312 : tmp6316);
  assign tmp6303 = s4 ? tmp6304 : tmp6311;
  assign tmp6302 = s5 ? tmp6268 : tmp6303;
  assign tmp6301 = s6 ? tmp6302 : tmp6115;
  assign tmp6299 = s7 ? tmp6300 : tmp6301;
  assign tmp6322 = s2 ? tmp6278 : tmp6307;
  assign tmp6321 = s3 ? tmp6322 : tmp6282;
  assign tmp6324 = s2 ? tmp6288 : tmp6314;
  assign tmp6323 = ~(s3 ? tmp6324 : tmp6316);
  assign tmp6320 = s4 ? tmp6321 : tmp6323;
  assign tmp6319 = s5 ? tmp6268 : tmp6320;
  assign tmp6318 = s6 ? tmp6115 : tmp6319;
  assign tmp6325 = s6 ? tmp6319 : tmp6302;
  assign tmp6317 = s7 ? tmp6318 : tmp6325;
  assign tmp6298 = s8 ? tmp6299 : tmp6317;
  assign tmp6266 = s9 ? tmp6267 : tmp6298;
  assign tmp6329 = s6 ? tmp6267 : tmp6302;
  assign tmp6328 = s7 ? tmp6300 : tmp6329;
  assign tmp6327 = s8 ? tmp6299 : tmp6328;
  assign tmp6326 = s9 ? tmp6267 : tmp6327;
  assign tmp6265 = s10 ? tmp6266 : tmp6326;
  assign tmp6335 = l1 ? tmp6076 : tmp6077;
  assign tmp6334 = s1 ? tmp6335 : tmp6123;
  assign tmp6338 = l1 ? tmp6120 : tmp6078;
  assign tmp6337 = s0 ? tmp6079 : tmp6338;
  assign tmp6336 = s1 ? tmp6123 : tmp6337;
  assign tmp6333 = s2 ? tmp6334 : tmp6336;
  assign tmp6343 = s0 ? tmp6079 : tmp6123;
  assign tmp6342 = s1 ? tmp6343 : tmp6133;
  assign tmp6345 = s0 ? tmp6335 : tmp6134;
  assign tmp6346 = s0 ? tmp6123 : tmp6091;
  assign tmp6344 = s1 ? tmp6345 : tmp6346;
  assign tmp6341 = s2 ? tmp6342 : tmp6344;
  assign tmp6349 = ~(s0 ? tmp6097 : tmp6123);
  assign tmp6348 = s1 ? tmp6095 : tmp6349;
  assign tmp6351 = l1 ? tmp6077 : tmp6088;
  assign tmp6352 = s0 ? tmp6079 : tmp6102;
  assign tmp6350 = s1 ? tmp6351 : tmp6352;
  assign tmp6347 = ~(s2 ? tmp6348 : tmp6350);
  assign tmp6340 = s3 ? tmp6341 : tmp6347;
  assign tmp6356 = ~(l1 ? tmp6120 : 1);
  assign tmp6355 = s1 ? tmp6106 : tmp6356;
  assign tmp6359 = l1 ? tmp6098 : tmp6076;
  assign tmp6358 = ~(s0 ? 1 : tmp6359);
  assign tmp6357 = ~(s1 ? tmp6123 : tmp6358);
  assign tmp6354 = s2 ? tmp6355 : tmp6357;
  assign tmp6361 = s0 ? tmp6097 : tmp6123;
  assign tmp6363 = ~(l1 ? tmp6120 : tmp6078);
  assign tmp6362 = ~(s0 ? tmp6079 : tmp6363);
  assign tmp6360 = ~(s1 ? tmp6361 : tmp6362);
  assign tmp6353 = ~(s3 ? tmp6354 : tmp6360);
  assign tmp6339 = s4 ? tmp6340 : tmp6353;
  assign tmp6332 = s5 ? tmp6333 : tmp6339;
  assign tmp6366 = s6 ? tmp6115 : tmp6332;
  assign tmp6372 = s1 ? tmp6343 : tmp6092;
  assign tmp6373 = s1 ? tmp6335 : tmp6346;
  assign tmp6371 = s2 ? tmp6372 : tmp6373;
  assign tmp6375 = s1 ? 1 : tmp6123;
  assign tmp6376 = ~(s1 ? tmp6351 : tmp6102);
  assign tmp6374 = s2 ? tmp6375 : tmp6376;
  assign tmp6370 = s3 ? tmp6371 : tmp6374;
  assign tmp6380 = ~(l1 ? tmp6098 : tmp6076);
  assign tmp6379 = ~(s1 ? tmp6123 : tmp6380);
  assign tmp6378 = s2 ? tmp6355 : tmp6379;
  assign tmp6381 = ~(s1 ? tmp6123 : tmp6338);
  assign tmp6377 = ~(s3 ? tmp6378 : tmp6381);
  assign tmp6369 = s4 ? tmp6370 : tmp6377;
  assign tmp6368 = s5 ? tmp6333 : tmp6369;
  assign tmp6367 = s6 ? tmp6368 : tmp6115;
  assign tmp6365 = s7 ? tmp6366 : tmp6367;
  assign tmp6387 = s2 ? tmp6342 : tmp6373;
  assign tmp6386 = s3 ? tmp6387 : tmp6347;
  assign tmp6385 = s4 ? tmp6386 : tmp6377;
  assign tmp6384 = s5 ? tmp6333 : tmp6385;
  assign tmp6383 = s6 ? tmp6115 : tmp6384;
  assign tmp6388 = s6 ? tmp6384 : tmp6368;
  assign tmp6382 = s7 ? tmp6383 : tmp6388;
  assign tmp6364 = s8 ? tmp6365 : tmp6382;
  assign tmp6331 = s9 ? tmp6332 : tmp6364;
  assign tmp6392 = s6 ? tmp6332 : tmp6368;
  assign tmp6391 = s7 ? tmp6366 : tmp6392;
  assign tmp6390 = s8 ? tmp6365 : tmp6391;
  assign tmp6389 = s9 ? tmp6332 : tmp6390;
  assign tmp6330 = s10 ? tmp6331 : tmp6389;
  assign tmp6264 = s11 ? tmp6265 : tmp6330;
  assign tmp6067 = s12 ? tmp6068 : tmp6264;
  assign tmp6401 = ~(l2 ? 1 : 0);
  assign tmp6400 = l1 ? tmp6120 : tmp6401;
  assign tmp6402 = l1 ? tmp6076 : tmp6401;
  assign tmp6399 = s1 ? tmp6400 : tmp6402;
  assign tmp6404 = s0 ? tmp6402 : tmp6202;
  assign tmp6406 = l1 ? tmp6076 : tmp6075;
  assign tmp6405 = s0 ? tmp6402 : tmp6406;
  assign tmp6403 = s1 ? tmp6404 : tmp6405;
  assign tmp6398 = s2 ? tmp6399 : tmp6403;
  assign tmp6410 = s1 ? tmp6402 : tmp6213;
  assign tmp6412 = s0 ? tmp6402 : tmp6213;
  assign tmp6411 = s1 ? tmp6400 : tmp6412;
  assign tmp6409 = s2 ? tmp6410 : tmp6411;
  assign tmp6414 = s1 ? tmp6216 : tmp6125;
  assign tmp6415 = ~(s1 ? tmp6218 : tmp6152);
  assign tmp6413 = ~(s2 ? tmp6414 : tmp6415);
  assign tmp6408 = s3 ? tmp6409 : tmp6413;
  assign tmp6420 = ~(l1 ? tmp6077 : tmp6120);
  assign tmp6419 = s0 ? tmp6152 : tmp6420;
  assign tmp6418 = s1 ? tmp6075 : tmp6419;
  assign tmp6421 = s1 ? tmp6402 : tmp6406;
  assign tmp6417 = s2 ? tmp6418 : tmp6421;
  assign tmp6424 = l1 ? tmp6077 : tmp6101;
  assign tmp6425 = ~(l1 ? tmp6076 : tmp6075);
  assign tmp6423 = s1 ? tmp6424 : tmp6425;
  assign tmp6426 = ~(l1 ? 1 : tmp6075);
  assign tmp6422 = ~(s2 ? tmp6423 : tmp6426);
  assign tmp6416 = s3 ? tmp6417 : tmp6422;
  assign tmp6407 = s4 ? tmp6408 : tmp6416;
  assign tmp6397 = s5 ? tmp6398 : tmp6407;
  assign tmp6430 = ~(s5 ? tmp6398 : tmp6407);
  assign tmp6429 = s6 ? tmp6115 : tmp6430;
  assign tmp6435 = l1 ? tmp6098 : tmp6101;
  assign tmp6434 = s1 ? tmp6435 : tmp6424;
  assign tmp6437 = s0 ? tmp6424 : tmp6077;
  assign tmp6439 = l1 ? tmp6077 : tmp6127;
  assign tmp6438 = s0 ? tmp6424 : tmp6439;
  assign tmp6436 = s1 ? tmp6437 : tmp6438;
  assign tmp6433 = s2 ? tmp6434 : tmp6436;
  assign tmp6443 = s1 ? tmp6424 : tmp6092;
  assign tmp6445 = s0 ? tmp6424 : tmp6092;
  assign tmp6444 = s1 ? tmp6435 : tmp6445;
  assign tmp6442 = s2 ? tmp6443 : tmp6444;
  assign tmp6448 = ~(l1 ? tmp6092 : tmp6127);
  assign tmp6447 = ~(s1 ? tmp6218 : tmp6448);
  assign tmp6446 = s2 ? tmp6414 : tmp6447;
  assign tmp6441 = s3 ? tmp6442 : tmp6446;
  assign tmp6451 = s1 ? tmp6075 : tmp6420;
  assign tmp6452 = ~(s1 ? tmp6424 : tmp6425);
  assign tmp6450 = s2 ? tmp6451 : tmp6452;
  assign tmp6453 = ~(s1 ? tmp6424 : tmp6439);
  assign tmp6449 = ~(s3 ? tmp6450 : tmp6453);
  assign tmp6440 = s4 ? tmp6441 : tmp6449;
  assign tmp6432 = s5 ? tmp6433 : tmp6440;
  assign tmp6431 = s6 ? tmp6432 : tmp6115;
  assign tmp6428 = s7 ? tmp6429 : tmp6431;
  assign tmp6458 = s3 ? tmp6417 : tmp6452;
  assign tmp6457 = s4 ? tmp6408 : tmp6458;
  assign tmp6456 = ~(s5 ? tmp6398 : tmp6457);
  assign tmp6455 = s6 ? tmp6115 : tmp6456;
  assign tmp6460 = s5 ? tmp6398 : tmp6457;
  assign tmp6461 = ~(s5 ? tmp6433 : tmp6440);
  assign tmp6459 = ~(s6 ? tmp6460 : tmp6461);
  assign tmp6454 = s7 ? tmp6455 : tmp6459;
  assign tmp6427 = ~(s8 ? tmp6428 : tmp6454);
  assign tmp6396 = s9 ? tmp6397 : tmp6427;
  assign tmp6465 = ~(s6 ? tmp6397 : tmp6461);
  assign tmp6464 = s7 ? tmp6429 : tmp6465;
  assign tmp6463 = ~(s8 ? tmp6428 : tmp6464);
  assign tmp6462 = s9 ? tmp6397 : tmp6463;
  assign tmp6395 = s10 ? tmp6396 : tmp6462;
  assign tmp6466 = ~(s10 ? tmp6070 : tmp6189);
  assign tmp6394 = s11 ? tmp6395 : tmp6466;
  assign tmp6473 = l1 ? 1 : tmp6401;
  assign tmp6474 = l1 ? tmp6075 : tmp6401;
  assign tmp6472 = s1 ? tmp6473 : tmp6474;
  assign tmp6477 = l1 ? tmp6075 : tmp6201;
  assign tmp6476 = s0 ? tmp6474 : tmp6477;
  assign tmp6478 = s0 ? tmp6402 : tmp6075;
  assign tmp6475 = s1 ? tmp6476 : tmp6478;
  assign tmp6471 = s2 ? tmp6472 : tmp6475;
  assign tmp6483 = s0 ? tmp6402 : tmp6474;
  assign tmp6482 = s1 ? tmp6483 : tmp6209;
  assign tmp6485 = s0 ? tmp6473 : tmp6079;
  assign tmp6486 = s0 ? tmp6474 : tmp6213;
  assign tmp6484 = s1 ? tmp6485 : tmp6486;
  assign tmp6481 = s2 ? tmp6482 : tmp6484;
  assign tmp6488 = s1 ? tmp6216 : tmp6119;
  assign tmp6490 = s0 ? tmp6120 : tmp6087;
  assign tmp6489 = s1 ? tmp6490 : tmp6426;
  assign tmp6487 = ~(s2 ? tmp6488 : tmp6489);
  assign tmp6480 = s3 ? tmp6481 : tmp6487;
  assign tmp6495 = ~(l1 ? tmp6101 : tmp6120);
  assign tmp6494 = s0 ? tmp6152 : tmp6495;
  assign tmp6493 = s1 ? tmp6075 : tmp6494;
  assign tmp6496 = s1 ? tmp6474 : tmp6075;
  assign tmp6492 = s2 ? tmp6493 : tmp6496;
  assign tmp6498 = s1 ? tmp6101 : tmp6127;
  assign tmp6499 = ~(s1 ? tmp6152 : tmp6153);
  assign tmp6497 = ~(s2 ? tmp6498 : tmp6499);
  assign tmp6491 = s3 ? tmp6492 : tmp6497;
  assign tmp6479 = s4 ? tmp6480 : tmp6491;
  assign tmp6470 = s5 ? tmp6471 : tmp6479;
  assign tmp6503 = ~(s5 ? tmp6471 : tmp6479);
  assign tmp6502 = s6 ? tmp6115 : tmp6503;
  assign tmp6508 = l1 ? tmp6092 : tmp6101;
  assign tmp6507 = s1 ? tmp6508 : tmp6101;
  assign tmp6511 = l1 ? tmp6101 : tmp6077;
  assign tmp6510 = s0 ? tmp6101 : tmp6511;
  assign tmp6513 = l1 ? tmp6101 : tmp6127;
  assign tmp6512 = s0 ? tmp6424 : tmp6513;
  assign tmp6509 = s1 ? tmp6510 : tmp6512;
  assign tmp6506 = s2 ? tmp6507 : tmp6509;
  assign tmp6518 = s0 ? tmp6424 : tmp6101;
  assign tmp6517 = s1 ? tmp6518 : tmp6092;
  assign tmp6520 = s0 ? tmp6101 : tmp6092;
  assign tmp6519 = s1 ? tmp6508 : tmp6520;
  assign tmp6516 = s2 ? tmp6517 : tmp6519;
  assign tmp6523 = l1 ? tmp6092 : tmp6127;
  assign tmp6522 = s1 ? tmp6490 : tmp6523;
  assign tmp6521 = s2 ? tmp6488 : tmp6522;
  assign tmp6515 = s3 ? tmp6516 : tmp6521;
  assign tmp6526 = s1 ? tmp6075 : tmp6495;
  assign tmp6527 = ~(s1 ? tmp6101 : tmp6127);
  assign tmp6525 = s2 ? tmp6526 : tmp6527;
  assign tmp6529 = s1 ? tmp6101 : tmp6513;
  assign tmp6528 = ~(s2 ? tmp6529 : tmp6120);
  assign tmp6524 = ~(s3 ? tmp6525 : tmp6528);
  assign tmp6514 = s4 ? tmp6515 : tmp6524;
  assign tmp6505 = s5 ? tmp6506 : tmp6514;
  assign tmp6504 = s6 ? tmp6505 : tmp6115;
  assign tmp6501 = s7 ? tmp6502 : tmp6504;
  assign tmp6536 = s1 ? tmp6473 : tmp6486;
  assign tmp6535 = s2 ? tmp6482 : tmp6536;
  assign tmp6534 = s3 ? tmp6535 : tmp6487;
  assign tmp6537 = s3 ? tmp6492 : tmp6527;
  assign tmp6533 = s4 ? tmp6534 : tmp6537;
  assign tmp6532 = ~(s5 ? tmp6471 : tmp6533);
  assign tmp6531 = s6 ? tmp6115 : tmp6532;
  assign tmp6543 = s1 ? tmp6518 : tmp6133;
  assign tmp6542 = s2 ? tmp6543 : tmp6519;
  assign tmp6541 = s3 ? tmp6542 : tmp6521;
  assign tmp6545 = s2 ? tmp6493 : tmp6527;
  assign tmp6546 = ~(s1 ? tmp6101 : tmp6513);
  assign tmp6544 = ~(s3 ? tmp6545 : tmp6546);
  assign tmp6540 = s4 ? tmp6541 : tmp6544;
  assign tmp6539 = s5 ? tmp6506 : tmp6540;
  assign tmp6549 = ~(s3 ? tmp6525 : tmp6546);
  assign tmp6548 = s4 ? tmp6515 : tmp6549;
  assign tmp6547 = s5 ? tmp6506 : tmp6548;
  assign tmp6538 = s6 ? tmp6539 : tmp6547;
  assign tmp6530 = s7 ? tmp6531 : tmp6538;
  assign tmp6500 = ~(s8 ? tmp6501 : tmp6530);
  assign tmp6469 = s9 ? tmp6470 : tmp6500;
  assign tmp6559 = s0 ? tmp6508 : tmp6134;
  assign tmp6558 = s1 ? tmp6559 : tmp6520;
  assign tmp6557 = s2 ? tmp6543 : tmp6558;
  assign tmp6556 = s3 ? tmp6557 : tmp6521;
  assign tmp6561 = ~(s2 ? tmp6529 : tmp6499);
  assign tmp6560 = ~(s3 ? tmp6545 : tmp6561);
  assign tmp6555 = s4 ? tmp6556 : tmp6560;
  assign tmp6554 = s5 ? tmp6506 : tmp6555;
  assign tmp6553 = s6 ? tmp6554 : tmp6505;
  assign tmp6552 = s7 ? tmp6502 : tmp6553;
  assign tmp6551 = ~(s8 ? tmp6501 : tmp6552);
  assign tmp6550 = s9 ? tmp6470 : tmp6551;
  assign tmp6468 = s10 ? tmp6469 : tmp6550;
  assign tmp6568 = s1 ? tmp6132 : tmp6087;
  assign tmp6569 = s1 ? tmp6118 : tmp6137;
  assign tmp6567 = s2 ? tmp6568 : tmp6569;
  assign tmp6571 = s1 ? tmp6351 : tmp6145;
  assign tmp6570 = ~(s2 ? tmp6139 : tmp6571);
  assign tmp6566 = s3 ? tmp6567 : tmp6570;
  assign tmp6574 = s1 ? tmp6075 : tmp6151;
  assign tmp6573 = s2 ? tmp6574 : tmp6154;
  assign tmp6576 = s1 ? tmp6161 : tmp6126;
  assign tmp6578 = ~(l1 ? tmp6092 : tmp6120);
  assign tmp6577 = ~(s1 ? tmp6152 : tmp6578);
  assign tmp6575 = ~(s2 ? tmp6576 : tmp6577);
  assign tmp6572 = ~(s3 ? tmp6573 : tmp6575);
  assign tmp6565 = s4 ? tmp6566 : tmp6572;
  assign tmp6564 = s5 ? tmp6116 : tmp6565;
  assign tmp6581 = s6 ? tmp6115 : tmp6564;
  assign tmp6587 = s1 ? tmp6132 : tmp6092;
  assign tmp6586 = s2 ? tmp6587 : tmp6569;
  assign tmp6589 = s1 ? 1 : tmp6119;
  assign tmp6590 = ~(s1 ? tmp6351 : tmp6145);
  assign tmp6588 = s2 ? tmp6589 : tmp6590;
  assign tmp6585 = s3 ? tmp6586 : tmp6588;
  assign tmp6593 = s1 ? tmp6075 : tmp6153;
  assign tmp6595 = ~(l1 ? tmp6098 : tmp6075);
  assign tmp6594 = ~(s1 ? tmp6119 : tmp6595);
  assign tmp6592 = s2 ? tmp6593 : tmp6594;
  assign tmp6596 = ~(s1 ? tmp6119 : tmp6126);
  assign tmp6591 = ~(s3 ? tmp6592 : tmp6596);
  assign tmp6584 = s4 ? tmp6585 : tmp6591;
  assign tmp6583 = s5 ? tmp6116 : tmp6584;
  assign tmp6582 = s6 ? tmp6583 : tmp6115;
  assign tmp6580 = s7 ? tmp6581 : tmp6582;
  assign tmp6603 = ~(s1 ? tmp6155 : tmp6595);
  assign tmp6602 = s2 ? tmp6574 : tmp6603;
  assign tmp6601 = ~(s3 ? tmp6602 : tmp6596);
  assign tmp6600 = s4 ? tmp6566 : tmp6601;
  assign tmp6599 = s5 ? tmp6116 : tmp6600;
  assign tmp6598 = s6 ? tmp6115 : tmp6599;
  assign tmp6607 = s3 ? tmp6586 : tmp6570;
  assign tmp6606 = s4 ? tmp6607 : tmp6601;
  assign tmp6605 = s5 ? tmp6116 : tmp6606;
  assign tmp6604 = s6 ? tmp6605 : tmp6583;
  assign tmp6597 = s7 ? tmp6598 : tmp6604;
  assign tmp6579 = s8 ? tmp6580 : tmp6597;
  assign tmp6563 = s9 ? tmp6564 : tmp6579;
  assign tmp6613 = s4 ? tmp6607 : tmp6572;
  assign tmp6612 = s5 ? tmp6116 : tmp6613;
  assign tmp6611 = s6 ? tmp6612 : tmp6583;
  assign tmp6610 = s7 ? tmp6581 : tmp6611;
  assign tmp6609 = s8 ? tmp6580 : tmp6610;
  assign tmp6608 = s9 ? tmp6564 : tmp6609;
  assign tmp6562 = ~(s10 ? tmp6563 : tmp6608);
  assign tmp6467 = s11 ? tmp6468 : tmp6562;
  assign tmp6393 = ~(s12 ? tmp6394 : tmp6467);
  assign tmp6066 = s13 ? tmp6067 : tmp6393;
  assign tmp6624 = s1 ? tmp6202 : tmp6213;
  assign tmp6623 = s2 ? tmp6624 : tmp6256;
  assign tmp6622 = s3 ? tmp6623 : tmp6214;
  assign tmp6621 = s4 ? tmp6622 : tmp6220;
  assign tmp6620 = s5 ? tmp6198 : tmp6621;
  assign tmp6626 = s7 ? tmp6114 : tmp6230;
  assign tmp6634 = s0 ? tmp6213 : tmp6079;
  assign tmp6633 = s1 ? tmp6202 : tmp6634;
  assign tmp6632 = s2 ? tmp6633 : tmp6210;
  assign tmp6637 = s0 ? 1 : tmp6223;
  assign tmp6636 = s1 ? tmp6637 : tmp6096;
  assign tmp6640 = ~(l1 ? tmp6120 : tmp6088);
  assign tmp6639 = s0 ? tmp6120 : tmp6640;
  assign tmp6641 = ~(s0 ? tmp6079 : tmp6219);
  assign tmp6638 = ~(s1 ? tmp6639 : tmp6641);
  assign tmp6635 = s2 ? tmp6636 : tmp6638;
  assign tmp6631 = s3 ? tmp6632 : tmp6635;
  assign tmp6645 = s0 ? tmp6150 : tmp6106;
  assign tmp6646 = s0 ? tmp6152 : tmp6223;
  assign tmp6644 = s1 ? tmp6645 : tmp6646;
  assign tmp6649 = ~(l1 ? tmp6076 : tmp6201);
  assign tmp6648 = s0 ? tmp6156 : tmp6649;
  assign tmp6650 = ~(s0 ? 1 : tmp6076);
  assign tmp6647 = ~(s1 ? tmp6648 : tmp6650);
  assign tmp6643 = s2 ? tmp6644 : tmp6647;
  assign tmp6653 = s0 ? tmp6097 : tmp6077;
  assign tmp6654 = ~(s0 ? tmp6079 : tmp6076);
  assign tmp6652 = s1 ? tmp6653 : tmp6654;
  assign tmp6651 = ~(s2 ? tmp6652 : tmp6164);
  assign tmp6642 = s3 ? tmp6643 : tmp6651;
  assign tmp6630 = s4 ? tmp6631 : tmp6642;
  assign tmp6629 = s5 ? tmp6198 : tmp6630;
  assign tmp6628 = s6 ? tmp6629 : tmp6620;
  assign tmp6655 = ~(s6 ? tmp6183 : tmp6231);
  assign tmp6627 = ~(s7 ? tmp6628 : tmp6655);
  assign tmp6625 = ~(s8 ? tmp6626 : tmp6627);
  assign tmp6619 = s9 ? tmp6620 : tmp6625;
  assign tmp6659 = ~(s6 ? tmp6071 : tmp6231);
  assign tmp6658 = ~(s7 ? tmp6628 : tmp6659);
  assign tmp6657 = ~(s8 ? tmp6626 : tmp6658);
  assign tmp6656 = s9 ? tmp6620 : tmp6657;
  assign tmp6618 = s10 ? tmp6619 : tmp6656;
  assign tmp6664 = s6 ? tmp6258 : tmp6259;
  assign tmp6663 = ~(s7 ? tmp6628 : tmp6664);
  assign tmp6662 = ~(s8 ? tmp6227 : tmp6663);
  assign tmp6661 = s9 ? tmp6620 : tmp6662;
  assign tmp6668 = s6 ? tmp6197 : tmp6259;
  assign tmp6667 = ~(s7 ? tmp6628 : tmp6668);
  assign tmp6666 = ~(s8 ? tmp6227 : tmp6667);
  assign tmp6665 = s9 ? tmp6620 : tmp6666;
  assign tmp6660 = s10 ? tmp6661 : tmp6665;
  assign tmp6617 = s11 ? tmp6618 : tmp6660;
  assign tmp6673 = s7 ? tmp6300 : tmp6230;
  assign tmp6675 = ~(s6 ? tmp6319 : tmp6231);
  assign tmp6674 = ~(s7 ? tmp6628 : tmp6675);
  assign tmp6672 = ~(s8 ? tmp6673 : tmp6674);
  assign tmp6671 = s9 ? tmp6620 : tmp6672;
  assign tmp6679 = ~(s6 ? tmp6267 : tmp6231);
  assign tmp6678 = ~(s7 ? tmp6628 : tmp6679);
  assign tmp6677 = ~(s8 ? tmp6673 : tmp6678);
  assign tmp6676 = s9 ? tmp6620 : tmp6677;
  assign tmp6670 = s10 ? tmp6671 : tmp6676;
  assign tmp6685 = l1 ? 1 : tmp6201;
  assign tmp6684 = s1 ? tmp6685 : tmp6477;
  assign tmp6687 = s0 ? tmp6202 : tmp6106;
  assign tmp6686 = s1 ? tmp6477 : tmp6687;
  assign tmp6683 = s2 ? tmp6684 : tmp6686;
  assign tmp6692 = s0 ? tmp6202 : tmp6477;
  assign tmp6691 = s1 ? tmp6692 : tmp6213;
  assign tmp6694 = s0 ? tmp6477 : tmp6213;
  assign tmp6693 = s1 ? tmp6685 : tmp6694;
  assign tmp6690 = s2 ? tmp6691 : tmp6693;
  assign tmp6696 = s1 ? tmp6216 : tmp6123;
  assign tmp6697 = ~(s1 ? tmp6213 : tmp6219);
  assign tmp6695 = ~(s2 ? tmp6696 : tmp6697);
  assign tmp6689 = s3 ? tmp6690 : tmp6695;
  assign tmp6701 = ~(l1 ? tmp6101 : 1);
  assign tmp6700 = s1 ? tmp6106 : tmp6701;
  assign tmp6702 = s1 ? tmp6477 : tmp6106;
  assign tmp6699 = s2 ? tmp6700 : tmp6702;
  assign tmp6704 = ~(l1 ? tmp6075 : tmp6076);
  assign tmp6703 = ~(s1 ? tmp6511 : tmp6704);
  assign tmp6698 = s3 ? tmp6699 : tmp6703;
  assign tmp6688 = s4 ? tmp6689 : tmp6698;
  assign tmp6682 = s5 ? tmp6683 : tmp6688;
  assign tmp6711 = l1 ? tmp6092 : tmp6077;
  assign tmp6710 = s1 ? tmp6711 : tmp6511;
  assign tmp6714 = l1 ? tmp6101 : tmp6078;
  assign tmp6713 = s0 ? tmp6077 : tmp6714;
  assign tmp6712 = s1 ? tmp6511 : tmp6713;
  assign tmp6709 = s2 ? tmp6710 : tmp6712;
  assign tmp6719 = s0 ? tmp6077 : tmp6511;
  assign tmp6718 = s1 ? tmp6719 : tmp6092;
  assign tmp6721 = s0 ? tmp6511 : tmp6092;
  assign tmp6720 = s1 ? tmp6711 : tmp6721;
  assign tmp6717 = s2 ? tmp6718 : tmp6720;
  assign tmp6723 = ~(s1 ? tmp6213 : tmp6246);
  assign tmp6722 = s2 ? tmp6696 : tmp6723;
  assign tmp6716 = s3 ? tmp6717 : tmp6722;
  assign tmp6725 = s2 ? tmp6700 : tmp6703;
  assign tmp6726 = ~(s1 ? tmp6511 : tmp6714);
  assign tmp6724 = ~(s3 ? tmp6725 : tmp6726);
  assign tmp6715 = s4 ? tmp6716 : tmp6724;
  assign tmp6708 = s5 ? tmp6709 : tmp6715;
  assign tmp6707 = s6 ? tmp6708 : tmp6115;
  assign tmp6706 = s7 ? tmp6366 : tmp6707;
  assign tmp6729 = ~(s5 ? tmp6683 : tmp6688);
  assign tmp6728 = s6 ? tmp6115 : tmp6729;
  assign tmp6730 = s6 ? tmp6384 : tmp6708;
  assign tmp6727 = s7 ? tmp6728 : tmp6730;
  assign tmp6705 = ~(s8 ? tmp6706 : tmp6727);
  assign tmp6681 = s9 ? tmp6682 : tmp6705;
  assign tmp6734 = s6 ? tmp6332 : tmp6708;
  assign tmp6733 = s7 ? tmp6728 : tmp6734;
  assign tmp6732 = ~(s8 ? tmp6706 : tmp6733);
  assign tmp6731 = s9 ? tmp6682 : tmp6732;
  assign tmp6680 = s10 ? tmp6681 : tmp6731;
  assign tmp6669 = s11 ? tmp6670 : tmp6680;
  assign tmp6616 = s12 ? tmp6617 : tmp6669;
  assign tmp6740 = s7 ? tmp6429 : tmp6230;
  assign tmp6742 = s6 ? tmp6460 : tmp6259;
  assign tmp6741 = ~(s7 ? tmp6628 : tmp6742);
  assign tmp6739 = ~(s8 ? tmp6740 : tmp6741);
  assign tmp6738 = s9 ? tmp6620 : tmp6739;
  assign tmp6746 = s6 ? tmp6397 : tmp6259;
  assign tmp6745 = ~(s7 ? tmp6628 : tmp6746);
  assign tmp6744 = ~(s8 ? tmp6740 : tmp6745);
  assign tmp6743 = s9 ? tmp6620 : tmp6744;
  assign tmp6737 = s10 ? tmp6738 : tmp6743;
  assign tmp6736 = s11 ? tmp6737 : tmp6618;
  assign tmp6751 = s7 ? tmp6502 : tmp6707;
  assign tmp6754 = s5 ? tmp6471 : tmp6533;
  assign tmp6755 = ~(s5 ? tmp6709 : tmp6715);
  assign tmp6753 = ~(s6 ? tmp6754 : tmp6755);
  assign tmp6752 = s7 ? tmp6728 : tmp6753;
  assign tmp6750 = ~(s8 ? tmp6751 : tmp6752);
  assign tmp6749 = s9 ? tmp6682 : tmp6750;
  assign tmp6759 = ~(s6 ? tmp6470 : tmp6755);
  assign tmp6758 = s7 ? tmp6728 : tmp6759;
  assign tmp6757 = ~(s8 ? tmp6751 : tmp6758);
  assign tmp6756 = s9 ? tmp6682 : tmp6757;
  assign tmp6748 = s10 ? tmp6749 : tmp6756;
  assign tmp6763 = s7 ? tmp6581 : tmp6707;
  assign tmp6765 = s6 ? tmp6599 : tmp6708;
  assign tmp6764 = s7 ? tmp6728 : tmp6765;
  assign tmp6762 = ~(s8 ? tmp6763 : tmp6764);
  assign tmp6761 = s9 ? tmp6682 : tmp6762;
  assign tmp6769 = s6 ? tmp6564 : tmp6708;
  assign tmp6768 = s7 ? tmp6728 : tmp6769;
  assign tmp6767 = ~(s8 ? tmp6763 : tmp6768);
  assign tmp6766 = s9 ? tmp6682 : tmp6767;
  assign tmp6760 = s10 ? tmp6761 : tmp6766;
  assign tmp6747 = s11 ? tmp6748 : tmp6760;
  assign tmp6735 = s12 ? tmp6736 : tmp6747;
  assign tmp6615 = s13 ? tmp6616 : tmp6735;
  assign tmp6782 = s1 ? tmp6095 : tmp6134;
  assign tmp6781 = ~(s2 ? tmp6782 : tmp6099);
  assign tmp6780 = s3 ? tmp6171 : tmp6781;
  assign tmp6783 = ~(s3 ? tmp6104 : tmp6180);
  assign tmp6779 = s4 ? tmp6780 : tmp6783;
  assign tmp6778 = s5 ? tmp6072 : tmp6779;
  assign tmp6777 = s6 ? tmp6778 : tmp6115;
  assign tmp6776 = s7 ? tmp6114 : tmp6777;
  assign tmp6787 = s4 ? tmp6780 : tmp6176;
  assign tmp6786 = s5 ? tmp6072 : tmp6787;
  assign tmp6785 = s6 ? tmp6186 : tmp6786;
  assign tmp6784 = s7 ? tmp6182 : tmp6785;
  assign tmp6775 = s8 ? tmp6776 : tmp6784;
  assign tmp6774 = s9 ? tmp6071 : tmp6775;
  assign tmp6791 = s6 ? tmp6193 : tmp6778;
  assign tmp6790 = s7 ? tmp6114 : tmp6791;
  assign tmp6789 = s8 ? tmp6776 : tmp6790;
  assign tmp6788 = s9 ? tmp6071 : tmp6789;
  assign tmp6773 = s10 ? tmp6774 : tmp6788;
  assign tmp6801 = s1 ? tmp6077 : tmp6133;
  assign tmp6803 = s0 ? tmp6234 : tmp6134;
  assign tmp6802 = s1 ? tmp6803 : tmp6243;
  assign tmp6800 = s2 ? tmp6801 : tmp6802;
  assign tmp6799 = s3 ? tmp6800 : tmp6244;
  assign tmp6798 = s4 ? tmp6799 : tmp6247;
  assign tmp6797 = s5 ? tmp6232 : tmp6798;
  assign tmp6796 = s6 ? tmp6797 : tmp6115;
  assign tmp6795 = s7 ? tmp6228 : tmp6796;
  assign tmp6809 = s2 ? tmp6801 : tmp6242;
  assign tmp6808 = s3 ? tmp6809 : tmp6244;
  assign tmp6807 = s4 ? tmp6808 : tmp6247;
  assign tmp6806 = ~(s5 ? tmp6232 : tmp6807);
  assign tmp6805 = ~(s6 ? tmp6258 : tmp6806);
  assign tmp6804 = s7 ? tmp6251 : tmp6805;
  assign tmp6794 = ~(s8 ? tmp6795 : tmp6804);
  assign tmp6793 = s9 ? tmp6197 : tmp6794;
  assign tmp6814 = ~(s5 ? tmp6232 : tmp6798);
  assign tmp6813 = ~(s6 ? tmp6197 : tmp6814);
  assign tmp6812 = s7 ? tmp6228 : tmp6813;
  assign tmp6811 = ~(s8 ? tmp6795 : tmp6812);
  assign tmp6810 = s9 ? tmp6197 : tmp6811;
  assign tmp6792 = ~(s10 ? tmp6793 : tmp6810);
  assign tmp6772 = s11 ? tmp6773 : tmp6792;
  assign tmp6825 = s1 ? tmp6149 : tmp6290;
  assign tmp6824 = s2 ? tmp6825 : tmp6314;
  assign tmp6827 = s1 ? tmp6125 : tmp6274;
  assign tmp6828 = ~(l1 ? 1 : tmp6098);
  assign tmp6826 = ~(s2 ? tmp6827 : tmp6828);
  assign tmp6823 = ~(s3 ? tmp6824 : tmp6826);
  assign tmp6822 = s4 ? tmp6304 : tmp6823;
  assign tmp6821 = s5 ? tmp6268 : tmp6822;
  assign tmp6820 = s6 ? tmp6821 : tmp6115;
  assign tmp6819 = s7 ? tmp6300 : tmp6820;
  assign tmp6833 = ~(s3 ? tmp6824 : tmp6316);
  assign tmp6832 = s4 ? tmp6304 : tmp6833;
  assign tmp6831 = s5 ? tmp6268 : tmp6832;
  assign tmp6830 = s6 ? tmp6319 : tmp6831;
  assign tmp6829 = s7 ? tmp6318 : tmp6830;
  assign tmp6818 = s8 ? tmp6819 : tmp6829;
  assign tmp6817 = s9 ? tmp6267 : tmp6818;
  assign tmp6837 = s6 ? tmp6267 : tmp6821;
  assign tmp6836 = s7 ? tmp6300 : tmp6837;
  assign tmp6835 = s8 ? tmp6819 : tmp6836;
  assign tmp6834 = s9 ? tmp6267 : tmp6835;
  assign tmp6816 = s10 ? tmp6817 : tmp6834;
  assign tmp6847 = ~(s1 ? tmp6351 : tmp6352);
  assign tmp6846 = s2 ? tmp6375 : tmp6847;
  assign tmp6845 = s3 ? tmp6371 : tmp6846;
  assign tmp6849 = ~(s1 ? tmp6123 : tmp6362);
  assign tmp6848 = ~(s3 ? tmp6378 : tmp6849);
  assign tmp6844 = s4 ? tmp6845 : tmp6848;
  assign tmp6843 = s5 ? tmp6333 : tmp6844;
  assign tmp6842 = s6 ? tmp6843 : tmp6115;
  assign tmp6841 = s7 ? tmp6366 : tmp6842;
  assign tmp6853 = s4 ? tmp6845 : tmp6377;
  assign tmp6852 = s5 ? tmp6333 : tmp6853;
  assign tmp6851 = s6 ? tmp6384 : tmp6852;
  assign tmp6850 = s7 ? tmp6383 : tmp6851;
  assign tmp6840 = s8 ? tmp6841 : tmp6850;
  assign tmp6839 = s9 ? tmp6332 : tmp6840;
  assign tmp6857 = s6 ? tmp6332 : tmp6843;
  assign tmp6856 = s7 ? tmp6366 : tmp6857;
  assign tmp6855 = s8 ? tmp6841 : tmp6856;
  assign tmp6854 = s9 ? tmp6332 : tmp6855;
  assign tmp6838 = s10 ? tmp6839 : tmp6854;
  assign tmp6815 = s11 ? tmp6816 : tmp6838;
  assign tmp6771 = s12 ? tmp6772 : tmp6815;
  assign tmp6868 = s2 ? tmp6418 : tmp6452;
  assign tmp6870 = s1 ? tmp6424 : tmp6439;
  assign tmp6869 = ~(s2 ? tmp6870 : tmp6426);
  assign tmp6867 = ~(s3 ? tmp6868 : tmp6869);
  assign tmp6866 = s4 ? tmp6441 : tmp6867;
  assign tmp6865 = s5 ? tmp6433 : tmp6866;
  assign tmp6864 = s6 ? tmp6865 : tmp6115;
  assign tmp6863 = s7 ? tmp6429 : tmp6864;
  assign tmp6875 = ~(s3 ? tmp6868 : tmp6453);
  assign tmp6874 = s4 ? tmp6441 : tmp6875;
  assign tmp6873 = ~(s5 ? tmp6433 : tmp6874);
  assign tmp6872 = ~(s6 ? tmp6460 : tmp6873);
  assign tmp6871 = s7 ? tmp6455 : tmp6872;
  assign tmp6862 = ~(s8 ? tmp6863 : tmp6871);
  assign tmp6861 = s9 ? tmp6397 : tmp6862;
  assign tmp6880 = ~(s5 ? tmp6433 : tmp6866);
  assign tmp6879 = ~(s6 ? tmp6397 : tmp6880);
  assign tmp6878 = s7 ? tmp6429 : tmp6879;
  assign tmp6877 = ~(s8 ? tmp6863 : tmp6878);
  assign tmp6876 = s9 ? tmp6397 : tmp6877;
  assign tmp6860 = s10 ? tmp6861 : tmp6876;
  assign tmp6890 = s1 ? 1 : tmp6111;
  assign tmp6889 = s2 ? tmp6890 : tmp6175;
  assign tmp6888 = s3 ? tmp6171 : tmp6889;
  assign tmp6891 = ~(s3 ? tmp6177 : tmp6110);
  assign tmp6887 = s4 ? tmp6888 : tmp6891;
  assign tmp6886 = s5 ? tmp6072 : tmp6887;
  assign tmp6885 = s6 ? tmp6886 : tmp6115;
  assign tmp6884 = s7 ? tmp6114 : tmp6885;
  assign tmp6892 = s7 ? tmp6182 : tmp6186;
  assign tmp6883 = s8 ? tmp6884 : tmp6892;
  assign tmp6882 = s9 ? tmp6071 : tmp6883;
  assign tmp6895 = s7 ? tmp6114 : tmp6193;
  assign tmp6894 = s8 ? tmp6884 : tmp6895;
  assign tmp6893 = s9 ? tmp6071 : tmp6894;
  assign tmp6881 = ~(s10 ? tmp6882 : tmp6893);
  assign tmp6859 = s11 ? tmp6860 : tmp6881;
  assign tmp6905 = s2 ? tmp6593 : tmp6603;
  assign tmp6907 = s1 ? tmp6119 : tmp6126;
  assign tmp6906 = ~(s2 ? tmp6907 : tmp6156);
  assign tmp6904 = ~(s3 ? tmp6905 : tmp6906);
  assign tmp6903 = s4 ? tmp6585 : tmp6904;
  assign tmp6902 = s5 ? tmp6116 : tmp6903;
  assign tmp6901 = s6 ? tmp6902 : tmp6115;
  assign tmp6900 = s7 ? tmp6581 : tmp6901;
  assign tmp6912 = ~(s3 ? tmp6905 : tmp6596);
  assign tmp6911 = s4 ? tmp6585 : tmp6912;
  assign tmp6910 = s5 ? tmp6116 : tmp6911;
  assign tmp6909 = s6 ? tmp6605 : tmp6910;
  assign tmp6908 = s7 ? tmp6598 : tmp6909;
  assign tmp6899 = s8 ? tmp6900 : tmp6908;
  assign tmp6898 = s9 ? tmp6564 : tmp6899;
  assign tmp6916 = s6 ? tmp6612 : tmp6902;
  assign tmp6915 = s7 ? tmp6581 : tmp6916;
  assign tmp6914 = s8 ? tmp6900 : tmp6915;
  assign tmp6913 = s9 ? tmp6564 : tmp6914;
  assign tmp6897 = ~(s10 ? tmp6898 : tmp6913);
  assign tmp6896 = s11 ? tmp6468 : tmp6897;
  assign tmp6858 = ~(s12 ? tmp6859 : tmp6896);
  assign tmp6770 = ~(s13 ? tmp6771 : tmp6858);
  assign tmp6614 = ~(s15 ? tmp6615 : tmp6770);
  assign tmp6065 = s16 ? tmp6066 : tmp6614;
  assign s2n = tmp6065;

  assign tmp6927 = l3 ? 1 : 0;
  assign tmp6926 = l2 ? 1 : tmp6927;
  assign tmp6929 = ~(l3 ? 1 : 0);
  assign tmp6928 = ~(l2 ? tmp6927 : tmp6929);
  assign tmp6925 = l1 ? tmp6926 : tmp6928;
  assign tmp6933 = ~(l2 ? tmp6927 : 0);
  assign tmp6932 = l1 ? tmp6926 : tmp6933;
  assign tmp6931 = s0 ? tmp6925 : tmp6932;
  assign tmp6935 = l1 ? tmp6927 : tmp6928;
  assign tmp6934 = s0 ? tmp6935 : tmp6925;
  assign tmp6930 = s1 ? tmp6931 : tmp6934;
  assign tmp6924 = s2 ? tmp6925 : tmp6930;
  assign tmp6939 = s1 ? tmp6934 : tmp6933;
  assign tmp6942 = l1 ? tmp6927 : 0;
  assign tmp6941 = s0 ? tmp6925 : tmp6942;
  assign tmp6940 = s1 ? tmp6925 : tmp6941;
  assign tmp6938 = s2 ? tmp6939 : tmp6940;
  assign tmp6947 = l2 ? 1 : tmp6929;
  assign tmp6946 = l1 ? tmp6947 : tmp6933;
  assign tmp6948 = ~(l2 ? tmp6927 : 1);
  assign tmp6945 = s0 ? tmp6946 : tmp6948;
  assign tmp6949 = ~(s0 ? 1 : tmp6926);
  assign tmp6944 = s1 ? tmp6945 : tmp6949;
  assign tmp6951 = l1 ? 1 : tmp6926;
  assign tmp6950 = ~(s1 ? tmp6932 : tmp6951);
  assign tmp6943 = ~(s2 ? tmp6944 : tmp6950);
  assign tmp6937 = s3 ? tmp6938 : tmp6943;
  assign tmp6955 = l2 ? tmp6927 : 1;
  assign tmp6957 = l2 ? tmp6927 : tmp6929;
  assign tmp6956 = l1 ? tmp6957 : 1;
  assign tmp6954 = s1 ? tmp6955 : tmp6956;
  assign tmp6960 = l1 ? tmp6957 : tmp6955;
  assign tmp6959 = ~(s0 ? tmp6946 : tmp6960);
  assign tmp6958 = ~(s1 ? tmp6925 : tmp6959);
  assign tmp6953 = s2 ? tmp6954 : tmp6958;
  assign tmp6962 = s0 ? 1 : tmp6925;
  assign tmp6961 = ~(s1 ? tmp6962 : tmp6925);
  assign tmp6952 = ~(s3 ? tmp6953 : tmp6961);
  assign tmp6936 = s4 ? tmp6937 : tmp6952;
  assign tmp6923 = s5 ? tmp6924 : tmp6936;
  assign tmp6970 = ~(l2 ? 1 : tmp6927);
  assign tmp6969 = l1 ? 1 : tmp6970;
  assign tmp6971 = l1 ? tmp6955 : tmp6970;
  assign tmp6968 = s1 ? tmp6969 : tmp6971;
  assign tmp6974 = l1 ? 1 : tmp6929;
  assign tmp6973 = s0 ? tmp6971 : tmp6974;
  assign tmp6976 = l1 ? tmp6927 : tmp6970;
  assign tmp6975 = s0 ? tmp6976 : tmp6971;
  assign tmp6972 = s1 ? tmp6973 : tmp6975;
  assign tmp6967 = s2 ? tmp6968 : tmp6972;
  assign tmp6983 = l2 ? tmp6927 : 0;
  assign tmp6984 = ~(l2 ? 1 : tmp6929);
  assign tmp6982 = ~(l1 ? tmp6983 : tmp6984);
  assign tmp6981 = s0 ? tmp6974 : tmp6982;
  assign tmp6980 = s1 ? tmp6975 : tmp6981;
  assign tmp6986 = s0 ? tmp6969 : tmp6982;
  assign tmp6987 = s0 ? tmp6971 : tmp6942;
  assign tmp6985 = s1 ? tmp6986 : tmp6987;
  assign tmp6979 = s2 ? tmp6980 : tmp6985;
  assign tmp6991 = l1 ? 1 : tmp6947;
  assign tmp6990 = ~(s0 ? 1 : tmp6991);
  assign tmp6989 = s1 ? tmp6945 : tmp6990;
  assign tmp6995 = l2 ? 1 : 0;
  assign tmp6994 = l1 ? tmp6926 : tmp6995;
  assign tmp6993 = s0 ? tmp6994 : tmp6974;
  assign tmp6997 = l1 ? tmp6926 : tmp6947;
  assign tmp6998 = l1 ? 1 : tmp6957;
  assign tmp6996 = s0 ? tmp6997 : tmp6998;
  assign tmp6992 = ~(s1 ? tmp6993 : tmp6996);
  assign tmp6988 = ~(s2 ? tmp6989 : tmp6992);
  assign tmp6978 = s3 ? tmp6979 : tmp6988;
  assign tmp7004 = ~(l2 ? 1 : 0);
  assign tmp7003 = l1 ? tmp6983 : tmp7004;
  assign tmp7002 = s0 ? tmp7003 : tmp6951;
  assign tmp7006 = l1 ? tmp6995 : tmp6926;
  assign tmp7005 = s0 ? tmp6955 : tmp7006;
  assign tmp7001 = s1 ? tmp7002 : tmp7005;
  assign tmp7009 = ~(l1 ? tmp6955 : tmp6970);
  assign tmp7008 = s0 ? tmp6956 : tmp7009;
  assign tmp7010 = s0 ? tmp6946 : tmp7006;
  assign tmp7007 = s1 ? tmp7008 : tmp7010;
  assign tmp7000 = s2 ? tmp7001 : tmp7007;
  assign tmp7014 = l1 ? tmp6955 : tmp6929;
  assign tmp7013 = s0 ? 1 : tmp7014;
  assign tmp7015 = s0 ? tmp6997 : tmp6971;
  assign tmp7012 = s1 ? tmp7013 : tmp7015;
  assign tmp7017 = s0 ? tmp7003 : tmp6955;
  assign tmp7019 = ~(l1 ? tmp6957 : 1);
  assign tmp7018 = ~(s0 ? tmp6994 : tmp7019);
  assign tmp7016 = ~(s1 ? tmp7017 : tmp7018);
  assign tmp7011 = ~(s2 ? tmp7012 : tmp7016);
  assign tmp6999 = ~(s3 ? tmp7000 : tmp7011);
  assign tmp6977 = s4 ? tmp6978 : tmp6999;
  assign tmp6966 = s5 ? tmp6967 : tmp6977;
  assign tmp6965 = s6 ? tmp6966 : tmp6923;
  assign tmp7024 = l1 ? tmp6926 : tmp6984;
  assign tmp7025 = l1 ? tmp6927 : tmp6984;
  assign tmp7023 = s1 ? tmp7024 : tmp7025;
  assign tmp7027 = s0 ? tmp7025 : tmp6932;
  assign tmp7026 = s1 ? tmp7027 : tmp7025;
  assign tmp7022 = s2 ? tmp7023 : tmp7026;
  assign tmp7032 = l1 ? 1 : tmp6933;
  assign tmp7031 = s1 ? tmp7025 : tmp7032;
  assign tmp7034 = s0 ? tmp7025 : tmp6942;
  assign tmp7033 = s1 ? tmp7024 : tmp7034;
  assign tmp7030 = s2 ? tmp7031 : tmp7033;
  assign tmp7036 = s1 ? tmp6955 : tmp6926;
  assign tmp7038 = l1 ? 1 : tmp6927;
  assign tmp7037 = s1 ? tmp6932 : tmp7038;
  assign tmp7035 = s2 ? tmp7036 : tmp7037;
  assign tmp7029 = s3 ? tmp7030 : tmp7035;
  assign tmp7042 = l1 ? tmp6947 : 1;
  assign tmp7041 = s1 ? 1 : tmp7042;
  assign tmp7044 = ~(l1 ? tmp6947 : 1);
  assign tmp7043 = ~(s1 ? tmp7025 : tmp7044);
  assign tmp7040 = s2 ? tmp7041 : tmp7043;
  assign tmp7045 = ~(s1 ? tmp6935 : tmp7025);
  assign tmp7039 = ~(s3 ? tmp7040 : tmp7045);
  assign tmp7028 = s4 ? tmp7029 : tmp7039;
  assign tmp7021 = s5 ? tmp7022 : tmp7028;
  assign tmp7020 = s6 ? tmp7021 : tmp6966;
  assign tmp6964 = s7 ? tmp6965 : tmp7020;
  assign tmp7053 = ~(l1 ? tmp6957 : tmp6955);
  assign tmp7052 = ~(s1 ? tmp6925 : tmp7053);
  assign tmp7051 = s2 ? tmp6954 : tmp7052;
  assign tmp7054 = ~(l1 ? tmp6926 : tmp6928);
  assign tmp7050 = ~(s3 ? tmp7051 : tmp7054);
  assign tmp7049 = s4 ? tmp6937 : tmp7050;
  assign tmp7048 = s5 ? tmp6924 : tmp7049;
  assign tmp7047 = s6 ? tmp6966 : tmp7048;
  assign tmp7060 = ~(s1 ? tmp6932 : tmp7038);
  assign tmp7059 = ~(s2 ? tmp6944 : tmp7060);
  assign tmp7058 = s3 ? tmp7030 : tmp7059;
  assign tmp7057 = s4 ? tmp7058 : tmp7039;
  assign tmp7056 = s5 ? tmp7022 : tmp7057;
  assign tmp7055 = s6 ? tmp7056 : tmp7021;
  assign tmp7046 = s7 ? tmp7047 : tmp7055;
  assign tmp6963 = s8 ? tmp6964 : tmp7046;
  assign tmp6922 = s9 ? tmp6923 : tmp6963;
  assign tmp7070 = ~(s0 ? tmp6946 : tmp7042);
  assign tmp7069 = ~(s1 ? tmp7025 : tmp7070);
  assign tmp7068 = s2 ? tmp7041 : tmp7069;
  assign tmp7072 = s0 ? 1 : tmp6935;
  assign tmp7071 = ~(s1 ? tmp7072 : tmp7025);
  assign tmp7067 = ~(s3 ? tmp7068 : tmp7071);
  assign tmp7066 = s4 ? tmp7058 : tmp7067;
  assign tmp7065 = s5 ? tmp7022 : tmp7066;
  assign tmp7064 = s6 ? tmp7065 : tmp7021;
  assign tmp7063 = s7 ? tmp6965 : tmp7064;
  assign tmp7062 = s8 ? tmp6964 : tmp7063;
  assign tmp7061 = s9 ? tmp6923 : tmp7062;
  assign tmp6921 = s10 ? tmp6922 : tmp7061;
  assign tmp7079 = l1 ? tmp6955 : tmp6927;
  assign tmp7078 = s0 ? tmp6955 : tmp7079;
  assign tmp7081 = l1 ? 1 : tmp6955;
  assign tmp7080 = s0 ? tmp7081 : tmp6955;
  assign tmp7077 = s1 ? tmp7078 : tmp7080;
  assign tmp7076 = s2 ? tmp6955 : tmp7077;
  assign tmp7086 = ~(s0 ? tmp6974 : tmp6982);
  assign tmp7085 = s1 ? tmp6955 : tmp7086;
  assign tmp7089 = l1 ? tmp6983 : tmp6984;
  assign tmp7088 = s0 ? tmp6955 : tmp7089;
  assign tmp7090 = s0 ? tmp6955 : 1;
  assign tmp7087 = s1 ? tmp7088 : tmp7090;
  assign tmp7084 = s2 ? tmp7085 : tmp7087;
  assign tmp7092 = s1 ? tmp7042 : tmp6994;
  assign tmp7094 = l1 ? tmp6995 : tmp6929;
  assign tmp7095 = ~(l1 ? tmp6927 : tmp7004);
  assign tmp7093 = s1 ? tmp7094 : tmp7095;
  assign tmp7091 = ~(s2 ? tmp7092 : tmp7093);
  assign tmp7083 = s3 ? tmp7084 : tmp7091;
  assign tmp7099 = l1 ? tmp6955 : 1;
  assign tmp7098 = s1 ? tmp6955 : tmp7099;
  assign tmp7097 = s2 ? tmp7098 : tmp6955;
  assign tmp7101 = l1 ? tmp6995 : tmp6948;
  assign tmp7100 = ~(s1 ? tmp7101 : tmp6948);
  assign tmp7096 = s3 ? tmp7097 : tmp7100;
  assign tmp7082 = s4 ? tmp7083 : tmp7096;
  assign tmp7075 = s5 ? tmp7076 : tmp7082;
  assign tmp7105 = ~(s5 ? tmp7076 : tmp7082);
  assign tmp7104 = s6 ? tmp6966 : tmp7105;
  assign tmp7109 = l1 ? tmp6995 : 0;
  assign tmp7111 = s0 ? tmp7109 : tmp7094;
  assign tmp7113 = l1 ? tmp6983 : 0;
  assign tmp7112 = s0 ? tmp7113 : tmp7109;
  assign tmp7110 = s1 ? tmp7111 : tmp7112;
  assign tmp7108 = s2 ? tmp7109 : tmp7110;
  assign tmp7117 = s1 ? tmp7109 : tmp6974;
  assign tmp7119 = s0 ? tmp7109 : tmp7113;
  assign tmp7118 = s1 ? tmp7109 : tmp7119;
  assign tmp7116 = s2 ? tmp7117 : tmp7118;
  assign tmp7122 = l1 ? tmp6947 : tmp6955;
  assign tmp7121 = s1 ? tmp7122 : tmp6994;
  assign tmp7124 = l1 ? tmp6947 : tmp6983;
  assign tmp7123 = s1 ? tmp7094 : tmp7124;
  assign tmp7120 = s2 ? tmp7121 : tmp7123;
  assign tmp7115 = s3 ? tmp7116 : tmp7120;
  assign tmp7128 = ~(l1 ? tmp6955 : 1);
  assign tmp7127 = ~(s1 ? tmp7109 : tmp7128);
  assign tmp7126 = s2 ? tmp7099 : tmp7127;
  assign tmp7129 = ~(s1 ? tmp7101 : tmp7109);
  assign tmp7125 = ~(s3 ? tmp7126 : tmp7129);
  assign tmp7114 = s4 ? tmp7115 : tmp7125;
  assign tmp7107 = s5 ? tmp7108 : tmp7114;
  assign tmp7106 = s6 ? tmp7107 : tmp6966;
  assign tmp7103 = s7 ? tmp7104 : tmp7106;
  assign tmp7135 = s2 ? tmp7085 : tmp7090;
  assign tmp7134 = s3 ? tmp7135 : tmp7091;
  assign tmp7133 = s4 ? tmp7134 : tmp7096;
  assign tmp7132 = ~(s5 ? tmp7076 : tmp7133);
  assign tmp7131 = s6 ? tmp6966 : tmp7132;
  assign tmp7137 = s5 ? tmp7076 : tmp7133;
  assign tmp7138 = ~(s5 ? tmp7108 : tmp7114);
  assign tmp7136 = ~(s6 ? tmp7137 : tmp7138);
  assign tmp7130 = s7 ? tmp7131 : tmp7136;
  assign tmp7102 = ~(s8 ? tmp7103 : tmp7130);
  assign tmp7074 = s9 ? tmp7075 : tmp7102;
  assign tmp7142 = ~(s6 ? tmp7075 : tmp7138);
  assign tmp7141 = s7 ? tmp7104 : tmp7142;
  assign tmp7140 = ~(s8 ? tmp7103 : tmp7141);
  assign tmp7139 = s9 ? tmp7075 : tmp7140;
  assign tmp7073 = ~(s10 ? tmp7074 : tmp7139);
  assign tmp6920 = s11 ? tmp6921 : tmp7073;
  assign tmp7148 = l1 ? tmp6926 : tmp6970;
  assign tmp7151 = l1 ? tmp6926 : tmp6929;
  assign tmp7150 = s0 ? tmp7148 : tmp7151;
  assign tmp7152 = s0 ? tmp6976 : tmp7148;
  assign tmp7149 = s1 ? tmp7150 : tmp7152;
  assign tmp7147 = s2 ? tmp7148 : tmp7149;
  assign tmp7156 = s1 ? tmp7152 : tmp6981;
  assign tmp7158 = s0 ? tmp7148 : tmp6982;
  assign tmp7159 = s0 ? tmp7148 : tmp6942;
  assign tmp7157 = s1 ? tmp7158 : tmp7159;
  assign tmp7155 = s2 ? tmp7156 : tmp7157;
  assign tmp7162 = ~(s0 ? 1 : tmp6997);
  assign tmp7161 = s1 ? tmp6945 : tmp7162;
  assign tmp7163 = ~(s1 ? tmp7151 : tmp6998);
  assign tmp7160 = ~(s2 ? tmp7161 : tmp7163);
  assign tmp7154 = s3 ? tmp7155 : tmp7160;
  assign tmp7168 = l1 ? tmp6957 : tmp6926;
  assign tmp7167 = s0 ? tmp6955 : tmp7168;
  assign tmp7166 = s1 ? tmp7002 : tmp7167;
  assign tmp7170 = ~(s0 ? tmp6946 : tmp7168);
  assign tmp7169 = ~(s1 ? tmp7148 : tmp7170);
  assign tmp7165 = s2 ? tmp7166 : tmp7169;
  assign tmp7173 = s0 ? 1 : tmp7151;
  assign tmp7172 = s1 ? tmp7173 : tmp7148;
  assign tmp7174 = ~(s0 ? tmp7003 : tmp6955);
  assign tmp7171 = ~(s2 ? tmp7172 : tmp7174);
  assign tmp7164 = ~(s3 ? tmp7165 : tmp7171);
  assign tmp7153 = s4 ? tmp7154 : tmp7164;
  assign tmp7146 = s5 ? tmp7147 : tmp7153;
  assign tmp7177 = s6 ? tmp6966 : tmp7146;
  assign tmp7181 = s1 ? tmp7148 : tmp6976;
  assign tmp7183 = s0 ? tmp6976 : tmp7151;
  assign tmp7182 = s1 ? tmp7183 : tmp6976;
  assign tmp7180 = s2 ? tmp7181 : tmp7182;
  assign tmp7187 = s1 ? tmp6976 : tmp6974;
  assign tmp7189 = s0 ? tmp6976 : tmp6942;
  assign tmp7188 = s1 ? tmp7148 : tmp7189;
  assign tmp7186 = s2 ? tmp7187 : tmp7188;
  assign tmp7191 = s1 ? tmp6955 : tmp6997;
  assign tmp7192 = s1 ? tmp7151 : tmp6998;
  assign tmp7190 = s2 ? tmp7191 : tmp7192;
  assign tmp7185 = s3 ? tmp7186 : tmp7190;
  assign tmp7196 = l1 ? tmp6947 : tmp6926;
  assign tmp7195 = s1 ? tmp6951 : tmp7196;
  assign tmp7198 = ~(l1 ? tmp6947 : tmp6926);
  assign tmp7197 = ~(s1 ? tmp6976 : tmp7198);
  assign tmp7194 = s2 ? tmp7195 : tmp7197;
  assign tmp7200 = l1 ? tmp6927 : tmp6929;
  assign tmp7199 = ~(s1 ? tmp7200 : tmp6976);
  assign tmp7193 = ~(s3 ? tmp7194 : tmp7199);
  assign tmp7184 = s4 ? tmp7185 : tmp7193;
  assign tmp7179 = s5 ? tmp7180 : tmp7184;
  assign tmp7178 = s6 ? tmp7179 : tmp6966;
  assign tmp7176 = s7 ? tmp7177 : tmp7178;
  assign tmp7207 = s1 ? tmp7148 : tmp7159;
  assign tmp7206 = s2 ? tmp7156 : tmp7207;
  assign tmp7205 = s3 ? tmp7206 : tmp7160;
  assign tmp7211 = ~(l1 ? tmp6957 : tmp6926);
  assign tmp7210 = ~(s1 ? tmp7148 : tmp7211);
  assign tmp7209 = s2 ? tmp7166 : tmp7210;
  assign tmp7212 = ~(s1 ? tmp7151 : tmp7148);
  assign tmp7208 = ~(s3 ? tmp7209 : tmp7212);
  assign tmp7204 = s4 ? tmp7205 : tmp7208;
  assign tmp7203 = s5 ? tmp7147 : tmp7204;
  assign tmp7202 = s6 ? tmp6966 : tmp7203;
  assign tmp7218 = s1 ? tmp6976 : tmp6981;
  assign tmp7217 = s2 ? tmp7218 : tmp7188;
  assign tmp7216 = s3 ? tmp7217 : tmp7160;
  assign tmp7222 = s0 ? tmp6955 : tmp7196;
  assign tmp7221 = s1 ? tmp7002 : tmp7222;
  assign tmp7220 = s2 ? tmp7221 : tmp7197;
  assign tmp7219 = ~(s3 ? tmp7220 : tmp7199);
  assign tmp7215 = s4 ? tmp7216 : tmp7219;
  assign tmp7214 = s5 ? tmp7180 : tmp7215;
  assign tmp7213 = s6 ? tmp7214 : tmp7179;
  assign tmp7201 = s7 ? tmp7202 : tmp7213;
  assign tmp7175 = s8 ? tmp7176 : tmp7201;
  assign tmp7145 = s9 ? tmp7146 : tmp7175;
  assign tmp7231 = s1 ? tmp7158 : tmp7189;
  assign tmp7230 = s2 ? tmp7218 : tmp7231;
  assign tmp7229 = s3 ? tmp7230 : tmp7160;
  assign tmp7235 = ~(s0 ? tmp6946 : tmp7196);
  assign tmp7234 = ~(s1 ? tmp6976 : tmp7235);
  assign tmp7233 = s2 ? tmp7221 : tmp7234;
  assign tmp7238 = s0 ? 1 : tmp7200;
  assign tmp7237 = s1 ? tmp7238 : tmp6976;
  assign tmp7236 = ~(s2 ? tmp7237 : tmp7174);
  assign tmp7232 = ~(s3 ? tmp7233 : tmp7236);
  assign tmp7228 = s4 ? tmp7229 : tmp7232;
  assign tmp7227 = s5 ? tmp7180 : tmp7228;
  assign tmp7226 = s6 ? tmp7227 : tmp7179;
  assign tmp7225 = s7 ? tmp7177 : tmp7226;
  assign tmp7224 = s8 ? tmp7176 : tmp7225;
  assign tmp7223 = s9 ? tmp7146 : tmp7224;
  assign tmp7144 = s10 ? tmp7145 : tmp7223;
  assign tmp7244 = l1 ? 1 : tmp6948;
  assign tmp7245 = l1 ? tmp6955 : tmp6948;
  assign tmp7243 = s1 ? tmp7244 : tmp7245;
  assign tmp7247 = s0 ? tmp7245 : tmp6974;
  assign tmp7249 = l1 ? tmp6927 : tmp6948;
  assign tmp7248 = s0 ? tmp7249 : tmp7245;
  assign tmp7246 = s1 ? tmp7247 : tmp7248;
  assign tmp7242 = s2 ? tmp7243 : tmp7246;
  assign tmp7253 = s1 ? tmp7248 : tmp6981;
  assign tmp7255 = s0 ? tmp7244 : tmp6982;
  assign tmp7256 = s0 ? tmp7245 : tmp6942;
  assign tmp7254 = s1 ? tmp7255 : tmp7256;
  assign tmp7252 = s2 ? tmp7253 : tmp7254;
  assign tmp7260 = l1 ? 1 : tmp6995;
  assign tmp7259 = ~(s0 ? 1 : tmp7260);
  assign tmp7258 = s1 ? tmp6945 : tmp7259;
  assign tmp7262 = s0 ? tmp6997 : tmp7260;
  assign tmp7261 = ~(s1 ? tmp6974 : tmp7262);
  assign tmp7257 = ~(s2 ? tmp7258 : tmp7261);
  assign tmp7251 = s3 ? tmp7252 : tmp7257;
  assign tmp7266 = l1 ? tmp6995 : 1;
  assign tmp7265 = s1 ? tmp7081 : tmp7266;
  assign tmp7269 = l1 ? tmp6995 : tmp6955;
  assign tmp7268 = ~(s0 ? tmp6946 : tmp7269);
  assign tmp7267 = ~(s1 ? tmp7245 : tmp7268);
  assign tmp7264 = s2 ? tmp7265 : tmp7267;
  assign tmp7271 = s0 ? 1 : tmp7245;
  assign tmp7272 = s0 ? tmp6997 : tmp7245;
  assign tmp7270 = ~(s1 ? tmp7271 : tmp7272);
  assign tmp7263 = ~(s3 ? tmp7264 : tmp7270);
  assign tmp7250 = s4 ? tmp7251 : tmp7263;
  assign tmp7241 = s5 ? tmp7242 : tmp7250;
  assign tmp7275 = s6 ? tmp6966 : tmp7241;
  assign tmp7280 = l1 ? 1 : 0;
  assign tmp7281 = l1 ? tmp6955 : 0;
  assign tmp7279 = s1 ? tmp7280 : tmp7281;
  assign tmp7283 = s0 ? tmp7281 : tmp6974;
  assign tmp7284 = s0 ? tmp6942 : tmp7281;
  assign tmp7282 = s1 ? tmp7283 : tmp7284;
  assign tmp7278 = s2 ? tmp7279 : tmp7282;
  assign tmp7288 = s1 ? tmp7284 : tmp6974;
  assign tmp7290 = s0 ? tmp7281 : tmp6942;
  assign tmp7289 = s1 ? tmp7280 : tmp7290;
  assign tmp7287 = s2 ? tmp7288 : tmp7289;
  assign tmp7292 = s1 ? tmp6955 : tmp7260;
  assign tmp7294 = l1 ? 1 : tmp6983;
  assign tmp7293 = s1 ? tmp6974 : tmp7294;
  assign tmp7291 = s2 ? tmp7292 : tmp7293;
  assign tmp7286 = s3 ? tmp7287 : tmp7291;
  assign tmp7297 = s1 ? 1 : tmp7266;
  assign tmp7299 = ~(l1 ? tmp6995 : 1);
  assign tmp7298 = ~(s1 ? tmp7281 : tmp7299);
  assign tmp7296 = s2 ? tmp7297 : tmp7298;
  assign tmp7300 = ~(s1 ? tmp7245 : tmp7281);
  assign tmp7295 = ~(s3 ? tmp7296 : tmp7300);
  assign tmp7285 = s4 ? tmp7286 : tmp7295;
  assign tmp7277 = s5 ? tmp7278 : tmp7285;
  assign tmp7276 = s6 ? tmp7277 : tmp6966;
  assign tmp7274 = s7 ? tmp7275 : tmp7276;
  assign tmp7307 = s1 ? tmp7244 : tmp7256;
  assign tmp7306 = s2 ? tmp7253 : tmp7307;
  assign tmp7305 = s3 ? tmp7306 : tmp7257;
  assign tmp7311 = ~(l1 ? tmp6995 : tmp6955);
  assign tmp7310 = ~(s1 ? tmp7245 : tmp7311);
  assign tmp7309 = s2 ? tmp7265 : tmp7310;
  assign tmp7312 = ~(l1 ? tmp6955 : tmp6948);
  assign tmp7308 = ~(s3 ? tmp7309 : tmp7312);
  assign tmp7304 = s4 ? tmp7305 : tmp7308;
  assign tmp7303 = s5 ? tmp7242 : tmp7304;
  assign tmp7302 = s6 ? tmp6966 : tmp7303;
  assign tmp7318 = s1 ? tmp7284 : tmp6981;
  assign tmp7317 = s2 ? tmp7318 : tmp7289;
  assign tmp7321 = s0 ? tmp6997 : tmp7294;
  assign tmp7320 = ~(s1 ? tmp6974 : tmp7321);
  assign tmp7319 = ~(s2 ? tmp7258 : tmp7320);
  assign tmp7316 = s3 ? tmp7317 : tmp7319;
  assign tmp7315 = s4 ? tmp7316 : tmp7295;
  assign tmp7314 = s5 ? tmp7278 : tmp7315;
  assign tmp7313 = s6 ? tmp7314 : tmp7277;
  assign tmp7301 = s7 ? tmp7302 : tmp7313;
  assign tmp7273 = s8 ? tmp7274 : tmp7301;
  assign tmp7240 = s9 ? tmp7241 : tmp7273;
  assign tmp7331 = s0 ? tmp7280 : tmp6982;
  assign tmp7330 = s1 ? tmp7331 : tmp7290;
  assign tmp7329 = s2 ? tmp7318 : tmp7330;
  assign tmp7328 = s3 ? tmp7329 : tmp7319;
  assign tmp7335 = ~(s0 ? tmp6946 : tmp7266);
  assign tmp7334 = ~(s1 ? tmp7281 : tmp7335);
  assign tmp7333 = s2 ? tmp7297 : tmp7334;
  assign tmp7337 = s0 ? tmp6997 : tmp7281;
  assign tmp7336 = ~(s1 ? tmp7271 : tmp7337);
  assign tmp7332 = ~(s3 ? tmp7333 : tmp7336);
  assign tmp7327 = s4 ? tmp7328 : tmp7332;
  assign tmp7326 = s5 ? tmp7278 : tmp7327;
  assign tmp7325 = s6 ? tmp7326 : tmp7277;
  assign tmp7324 = s7 ? tmp7275 : tmp7325;
  assign tmp7323 = s8 ? tmp7274 : tmp7324;
  assign tmp7322 = s9 ? tmp7241 : tmp7323;
  assign tmp7239 = s10 ? tmp7240 : tmp7322;
  assign tmp7143 = s11 ? tmp7144 : tmp7239;
  assign tmp6919 = s12 ? tmp6920 : tmp7143;
  assign tmp7344 = l1 ? tmp6955 : tmp6995;
  assign tmp7347 = l1 ? tmp6955 : tmp6983;
  assign tmp7346 = s0 ? tmp7344 : tmp7347;
  assign tmp7348 = s0 ? tmp7260 : tmp7344;
  assign tmp7345 = s1 ? tmp7346 : tmp7348;
  assign tmp7343 = s2 ? tmp7344 : tmp7345;
  assign tmp7352 = s1 ? tmp7348 : tmp6983;
  assign tmp7353 = s0 ? tmp7344 : 1;
  assign tmp7351 = s2 ? tmp7352 : tmp7353;
  assign tmp7356 = l1 ? tmp6926 : 1;
  assign tmp7355 = s1 ? tmp7042 : tmp7356;
  assign tmp7358 = l1 ? tmp6995 : tmp6933;
  assign tmp7359 = ~(l1 ? tmp6927 : tmp6948);
  assign tmp7357 = s1 ? tmp7358 : tmp7359;
  assign tmp7354 = ~(s2 ? tmp7355 : tmp7357);
  assign tmp7350 = s3 ? tmp7351 : tmp7354;
  assign tmp7364 = l1 ? tmp6955 : tmp6926;
  assign tmp7363 = s0 ? tmp6955 : tmp7364;
  assign tmp7362 = s1 ? tmp6951 : tmp7363;
  assign tmp7365 = s1 ? tmp7344 : tmp7364;
  assign tmp7361 = s2 ? tmp7362 : tmp7365;
  assign tmp7368 = ~(l1 ? tmp6955 : tmp6995);
  assign tmp7367 = s1 ? tmp7358 : tmp7368;
  assign tmp7366 = ~(s2 ? tmp7367 : tmp6948);
  assign tmp7360 = s3 ? tmp7361 : tmp7366;
  assign tmp7349 = s4 ? tmp7350 : tmp7360;
  assign tmp7342 = s5 ? tmp7343 : tmp7349;
  assign tmp7372 = ~(s5 ? tmp7343 : tmp7349);
  assign tmp7371 = s6 ? tmp6966 : tmp7372;
  assign tmp7377 = l1 ? tmp6995 : tmp7004;
  assign tmp7376 = s1 ? tmp7377 : tmp7003;
  assign tmp7379 = s0 ? tmp7003 : tmp7358;
  assign tmp7378 = s1 ? tmp7379 : tmp7003;
  assign tmp7375 = s2 ? tmp7376 : tmp7378;
  assign tmp7383 = s1 ? tmp7003 : tmp7032;
  assign tmp7385 = s0 ? tmp7003 : tmp7113;
  assign tmp7384 = s1 ? tmp7377 : tmp7385;
  assign tmp7382 = s2 ? tmp7383 : tmp7384;
  assign tmp7387 = s1 ? tmp6960 : tmp7356;
  assign tmp7388 = s1 ? tmp7358 : tmp7122;
  assign tmp7386 = s2 ? tmp7387 : tmp7388;
  assign tmp7381 = s3 ? tmp7382 : tmp7386;
  assign tmp7392 = ~(l1 ? 1 : tmp6926);
  assign tmp7391 = ~(s1 ? tmp7003 : tmp7392);
  assign tmp7390 = s2 ? tmp6951 : tmp7391;
  assign tmp7394 = l1 ? tmp6983 : tmp6933;
  assign tmp7393 = ~(s1 ? tmp7394 : tmp7003);
  assign tmp7389 = ~(s3 ? tmp7390 : tmp7393);
  assign tmp7380 = s4 ? tmp7381 : tmp7389;
  assign tmp7374 = s5 ? tmp7375 : tmp7380;
  assign tmp7373 = s6 ? tmp7374 : tmp6966;
  assign tmp7370 = s7 ? tmp7371 : tmp7373;
  assign tmp7400 = ~(s1 ? tmp7358 : tmp7368);
  assign tmp7399 = s3 ? tmp7361 : tmp7400;
  assign tmp7398 = s4 ? tmp7350 : tmp7399;
  assign tmp7397 = ~(s5 ? tmp7343 : tmp7398);
  assign tmp7396 = s6 ? tmp6966 : tmp7397;
  assign tmp7402 = s5 ? tmp7343 : tmp7398;
  assign tmp7403 = ~(s5 ? tmp7375 : tmp7380);
  assign tmp7401 = ~(s6 ? tmp7402 : tmp7403);
  assign tmp7395 = s7 ? tmp7396 : tmp7401;
  assign tmp7369 = ~(s8 ? tmp7370 : tmp7395);
  assign tmp7341 = s9 ? tmp7342 : tmp7369;
  assign tmp7407 = ~(s6 ? tmp7342 : tmp7403);
  assign tmp7406 = s7 ? tmp7371 : tmp7407;
  assign tmp7405 = ~(s8 ? tmp7370 : tmp7406);
  assign tmp7404 = s9 ? tmp7342 : tmp7405;
  assign tmp7340 = s10 ? tmp7341 : tmp7404;
  assign tmp7408 = ~(s10 ? tmp6922 : tmp7061);
  assign tmp7339 = s11 ? tmp7340 : tmp7408;
  assign tmp7415 = l1 ? tmp6927 : tmp6926;
  assign tmp7414 = s1 ? tmp7415 : tmp6926;
  assign tmp7417 = s0 ? tmp6926 : tmp6927;
  assign tmp7418 = s0 ? tmp6951 : tmp6926;
  assign tmp7416 = s1 ? tmp7417 : tmp7418;
  assign tmp7413 = s2 ? tmp7414 : tmp7416;
  assign tmp7422 = s1 ? tmp7418 : tmp7086;
  assign tmp7424 = s0 ? tmp7415 : tmp7089;
  assign tmp7425 = s0 ? tmp6926 : 1;
  assign tmp7423 = s1 ? tmp7424 : tmp7425;
  assign tmp7421 = s2 ? tmp7422 : tmp7423;
  assign tmp7427 = s1 ? tmp7042 : tmp6991;
  assign tmp7430 = l1 ? tmp6947 : tmp6929;
  assign tmp7429 = s0 ? tmp6994 : tmp7430;
  assign tmp7431 = ~(l1 ? tmp6927 : tmp6928);
  assign tmp7428 = s1 ? tmp7429 : tmp7431;
  assign tmp7426 = ~(s2 ? tmp7427 : tmp7428);
  assign tmp7420 = s3 ? tmp7421 : tmp7426;
  assign tmp7435 = s0 ? tmp6955 : tmp6926;
  assign tmp7434 = s1 ? tmp6951 : tmp7435;
  assign tmp7433 = s2 ? tmp7434 : tmp6926;
  assign tmp7438 = l1 ? tmp6957 : tmp6929;
  assign tmp7437 = s1 ? tmp7438 : tmp6970;
  assign tmp7440 = ~(l1 ? tmp6926 : tmp6995);
  assign tmp7439 = ~(s1 ? tmp6955 : tmp7440);
  assign tmp7436 = ~(s2 ? tmp7437 : tmp7439);
  assign tmp7432 = s3 ? tmp7433 : tmp7436;
  assign tmp7419 = s4 ? tmp7420 : tmp7432;
  assign tmp7412 = s5 ? tmp7413 : tmp7419;
  assign tmp7444 = ~(s5 ? tmp7413 : tmp7419);
  assign tmp7443 = s6 ? tmp6966 : tmp7444;
  assign tmp7449 = l1 ? tmp6947 : tmp6970;
  assign tmp7450 = l1 ? tmp6957 : tmp6970;
  assign tmp7448 = s1 ? tmp7449 : tmp7450;
  assign tmp7452 = s0 ? tmp7450 : tmp7430;
  assign tmp7454 = l1 ? tmp6983 : tmp6970;
  assign tmp7453 = s0 ? tmp7454 : tmp7450;
  assign tmp7451 = s1 ? tmp7452 : tmp7453;
  assign tmp7447 = s2 ? tmp7448 : tmp7451;
  assign tmp7458 = s1 ? tmp7453 : tmp6974;
  assign tmp7460 = s0 ? tmp7450 : tmp7113;
  assign tmp7459 = s1 ? tmp7449 : tmp7460;
  assign tmp7457 = s2 ? tmp7458 : tmp7459;
  assign tmp7462 = s1 ? tmp6960 : tmp6991;
  assign tmp7464 = l1 ? tmp6947 : tmp6957;
  assign tmp7463 = s1 ? tmp7429 : tmp7464;
  assign tmp7461 = s2 ? tmp7462 : tmp7463;
  assign tmp7456 = s3 ? tmp7457 : tmp7461;
  assign tmp7467 = s1 ? tmp6951 : tmp6926;
  assign tmp7468 = ~(s1 ? tmp7450 : tmp6970);
  assign tmp7466 = s2 ? tmp7467 : tmp7468;
  assign tmp7470 = s1 ? tmp7438 : tmp7450;
  assign tmp7469 = ~(s2 ? tmp7470 : tmp6994);
  assign tmp7465 = ~(s3 ? tmp7466 : tmp7469);
  assign tmp7455 = s4 ? tmp7456 : tmp7465;
  assign tmp7446 = s5 ? tmp7447 : tmp7455;
  assign tmp7445 = s6 ? tmp7446 : tmp6966;
  assign tmp7442 = s7 ? tmp7443 : tmp7445;
  assign tmp7477 = s1 ? tmp7415 : tmp7425;
  assign tmp7476 = s2 ? tmp7422 : tmp7477;
  assign tmp7475 = s3 ? tmp7476 : tmp7426;
  assign tmp7479 = ~(s1 ? tmp7438 : tmp6970);
  assign tmp7478 = s3 ? tmp7433 : tmp7479;
  assign tmp7474 = s4 ? tmp7475 : tmp7478;
  assign tmp7473 = ~(s5 ? tmp7413 : tmp7474);
  assign tmp7472 = s6 ? tmp6966 : tmp7473;
  assign tmp7485 = s1 ? tmp7453 : tmp6981;
  assign tmp7484 = s2 ? tmp7485 : tmp7459;
  assign tmp7483 = s3 ? tmp7484 : tmp7461;
  assign tmp7487 = s2 ? tmp7434 : tmp7468;
  assign tmp7488 = ~(s1 ? tmp7438 : tmp7450);
  assign tmp7486 = ~(s3 ? tmp7487 : tmp7488);
  assign tmp7482 = s4 ? tmp7483 : tmp7486;
  assign tmp7481 = s5 ? tmp7447 : tmp7482;
  assign tmp7491 = ~(s3 ? tmp7466 : tmp7488);
  assign tmp7490 = s4 ? tmp7456 : tmp7491;
  assign tmp7489 = s5 ? tmp7447 : tmp7490;
  assign tmp7480 = s6 ? tmp7481 : tmp7489;
  assign tmp7471 = s7 ? tmp7472 : tmp7480;
  assign tmp7441 = ~(s8 ? tmp7442 : tmp7471);
  assign tmp7411 = s9 ? tmp7412 : tmp7441;
  assign tmp7501 = s0 ? tmp7449 : tmp6982;
  assign tmp7500 = s1 ? tmp7501 : tmp7460;
  assign tmp7499 = s2 ? tmp7485 : tmp7500;
  assign tmp7498 = s3 ? tmp7499 : tmp7461;
  assign tmp7503 = ~(s2 ? tmp7470 : tmp7439);
  assign tmp7502 = ~(s3 ? tmp7487 : tmp7503);
  assign tmp7497 = s4 ? tmp7498 : tmp7502;
  assign tmp7496 = s5 ? tmp7447 : tmp7497;
  assign tmp7495 = s6 ? tmp7496 : tmp7446;
  assign tmp7494 = s7 ? tmp7443 : tmp7495;
  assign tmp7493 = ~(s8 ? tmp7442 : tmp7494);
  assign tmp7492 = s9 ? tmp7412 : tmp7493;
  assign tmp7410 = s10 ? tmp7411 : tmp7492;
  assign tmp7509 = l1 ? 1 : tmp7004;
  assign tmp7510 = l1 ? tmp6955 : tmp7004;
  assign tmp7508 = s1 ? tmp7509 : tmp7510;
  assign tmp7512 = s0 ? tmp7510 : tmp7032;
  assign tmp7514 = l1 ? tmp6927 : tmp7004;
  assign tmp7513 = s0 ? tmp7514 : tmp7510;
  assign tmp7511 = s1 ? tmp7512 : tmp7513;
  assign tmp7507 = s2 ? tmp7508 : tmp7511;
  assign tmp7518 = s1 ? tmp7513 : tmp6933;
  assign tmp7520 = s0 ? tmp7510 : tmp6942;
  assign tmp7519 = s1 ? tmp7509 : tmp7520;
  assign tmp7517 = s2 ? tmp7518 : tmp7519;
  assign tmp7522 = s1 ? tmp6945 : 0;
  assign tmp7523 = ~(s1 ? tmp7032 : tmp7081);
  assign tmp7521 = ~(s2 ? tmp7522 : tmp7523);
  assign tmp7516 = s3 ? tmp7517 : tmp7521;
  assign tmp7526 = s1 ? tmp6951 : tmp7005;
  assign tmp7529 = ~(l1 ? tmp6955 : tmp7004);
  assign tmp7528 = s0 ? tmp6956 : tmp7529;
  assign tmp7527 = s1 ? tmp7528 : tmp7010;
  assign tmp7525 = s2 ? tmp7526 : tmp7527;
  assign tmp7533 = l1 ? tmp6955 : tmp6933;
  assign tmp7532 = s0 ? 1 : tmp7533;
  assign tmp7531 = s1 ? tmp7532 : tmp7510;
  assign tmp7534 = ~(s1 ? tmp6955 : tmp6956);
  assign tmp7530 = ~(s2 ? tmp7531 : tmp7534);
  assign tmp7524 = ~(s3 ? tmp7525 : tmp7530);
  assign tmp7515 = s4 ? tmp7516 : tmp7524;
  assign tmp7506 = s5 ? tmp7507 : tmp7515;
  assign tmp7537 = s6 ? tmp6966 : tmp7506;
  assign tmp7543 = s1 ? tmp7513 : tmp7032;
  assign tmp7542 = s2 ? tmp7543 : tmp7519;
  assign tmp7545 = s1 ? tmp6955 : 1;
  assign tmp7546 = s1 ? tmp7032 : tmp7081;
  assign tmp7544 = s2 ? tmp7545 : tmp7546;
  assign tmp7541 = s3 ? tmp7542 : tmp7544;
  assign tmp7549 = s1 ? tmp6951 : tmp7006;
  assign tmp7551 = ~(l1 ? tmp6995 : tmp6926);
  assign tmp7550 = ~(s1 ? tmp7510 : tmp7551);
  assign tmp7548 = s2 ? tmp7549 : tmp7550;
  assign tmp7552 = ~(s1 ? tmp7533 : tmp7510);
  assign tmp7547 = ~(s3 ? tmp7548 : tmp7552);
  assign tmp7540 = s4 ? tmp7541 : tmp7547;
  assign tmp7539 = s5 ? tmp7507 : tmp7540;
  assign tmp7538 = s6 ? tmp7539 : tmp6966;
  assign tmp7536 = s7 ? tmp7537 : tmp7538;
  assign tmp7559 = s1 ? tmp7528 : tmp7006;
  assign tmp7558 = s2 ? tmp7526 : tmp7559;
  assign tmp7557 = ~(s3 ? tmp7558 : tmp7552);
  assign tmp7556 = s4 ? tmp7516 : tmp7557;
  assign tmp7555 = s5 ? tmp7507 : tmp7556;
  assign tmp7554 = s6 ? tmp6966 : tmp7555;
  assign tmp7563 = s3 ? tmp7542 : tmp7521;
  assign tmp7562 = s4 ? tmp7563 : tmp7557;
  assign tmp7561 = s5 ? tmp7507 : tmp7562;
  assign tmp7560 = s6 ? tmp7561 : tmp7539;
  assign tmp7553 = s7 ? tmp7554 : tmp7560;
  assign tmp7535 = s8 ? tmp7536 : tmp7553;
  assign tmp7505 = s9 ? tmp7506 : tmp7535;
  assign tmp7569 = s4 ? tmp7563 : tmp7524;
  assign tmp7568 = s5 ? tmp7507 : tmp7569;
  assign tmp7567 = s6 ? tmp7568 : tmp7539;
  assign tmp7566 = s7 ? tmp7537 : tmp7567;
  assign tmp7565 = s8 ? tmp7536 : tmp7566;
  assign tmp7564 = s9 ? tmp7506 : tmp7565;
  assign tmp7504 = ~(s10 ? tmp7505 : tmp7564);
  assign tmp7409 = s11 ? tmp7410 : tmp7504;
  assign tmp7338 = ~(s12 ? tmp7339 : tmp7409);
  assign tmp6918 = s13 ? tmp6919 : tmp7338;
  assign tmp7578 = l1 ? tmp6955 : tmp6957;
  assign tmp7580 = s0 ? tmp7578 : tmp7347;
  assign tmp7581 = s0 ? tmp6998 : tmp7578;
  assign tmp7579 = s1 ? tmp7580 : tmp7581;
  assign tmp7577 = s2 ? tmp7578 : tmp7579;
  assign tmp7585 = s1 ? tmp7578 : tmp6983;
  assign tmp7586 = s0 ? tmp7578 : 1;
  assign tmp7584 = s2 ? tmp7585 : tmp7586;
  assign tmp7588 = s1 ? tmp7042 : tmp6926;
  assign tmp7590 = ~(l1 ? tmp6927 : tmp6970);
  assign tmp7589 = s1 ? tmp7358 : tmp7590;
  assign tmp7587 = ~(s2 ? tmp7588 : tmp7589);
  assign tmp7583 = s3 ? tmp7584 : tmp7587;
  assign tmp7593 = s1 ? tmp7578 : tmp6955;
  assign tmp7592 = s2 ? tmp7098 : tmp7593;
  assign tmp7595 = l1 ? tmp6995 : tmp6928;
  assign tmp7596 = ~(l1 ? tmp6955 : tmp6957);
  assign tmp7594 = ~(s1 ? tmp7595 : tmp7596);
  assign tmp7591 = s3 ? tmp7592 : tmp7594;
  assign tmp7582 = s4 ? tmp7583 : tmp7591;
  assign tmp7576 = s5 ? tmp7577 : tmp7582;
  assign tmp7603 = l1 ? tmp6995 : tmp6984;
  assign tmp7602 = s1 ? tmp7603 : tmp7089;
  assign tmp7605 = s0 ? tmp7089 : tmp7358;
  assign tmp7604 = s1 ? tmp7605 : tmp7089;
  assign tmp7601 = s2 ? tmp7602 : tmp7604;
  assign tmp7609 = s1 ? tmp7089 : tmp7032;
  assign tmp7611 = s0 ? tmp7089 : tmp7113;
  assign tmp7610 = s1 ? tmp7603 : tmp7611;
  assign tmp7608 = s2 ? tmp7609 : tmp7610;
  assign tmp7613 = s1 ? tmp6960 : tmp6926;
  assign tmp7615 = l1 ? tmp6947 : tmp6927;
  assign tmp7614 = s1 ? tmp7358 : tmp7615;
  assign tmp7612 = s2 ? tmp7613 : tmp7614;
  assign tmp7607 = s3 ? tmp7608 : tmp7612;
  assign tmp7618 = ~(s1 ? tmp7089 : 0);
  assign tmp7617 = s2 ? 1 : tmp7618;
  assign tmp7620 = l1 ? tmp6983 : tmp6928;
  assign tmp7619 = ~(s1 ? tmp7620 : tmp7089);
  assign tmp7616 = ~(s3 ? tmp7617 : tmp7619);
  assign tmp7606 = s4 ? tmp7607 : tmp7616;
  assign tmp7600 = s5 ? tmp7601 : tmp7606;
  assign tmp7599 = s6 ? tmp7600 : tmp6966;
  assign tmp7598 = s7 ? tmp6965 : tmp7599;
  assign tmp7628 = s0 ? tmp6983 : tmp7089;
  assign tmp7627 = s1 ? tmp7578 : tmp7628;
  assign tmp7630 = s0 ? tmp7578 : tmp7089;
  assign tmp7629 = s1 ? tmp7630 : tmp7586;
  assign tmp7626 = s2 ? tmp7627 : tmp7629;
  assign tmp7633 = s0 ? tmp6946 : tmp7044;
  assign tmp7632 = s1 ? tmp7633 : tmp6949;
  assign tmp7635 = s0 ? tmp6994 : tmp7358;
  assign tmp7636 = s0 ? tmp6997 : tmp7590;
  assign tmp7634 = ~(s1 ? tmp7635 : tmp7636);
  assign tmp7631 = s2 ? tmp7632 : tmp7634;
  assign tmp7625 = s3 ? tmp7626 : tmp7631;
  assign tmp7640 = s0 ? tmp6955 : tmp7099;
  assign tmp7639 = s1 ? tmp7017 : tmp7640;
  assign tmp7642 = s0 ? tmp6956 : tmp7578;
  assign tmp7643 = s0 ? tmp6946 : tmp6955;
  assign tmp7641 = s1 ? tmp7642 : tmp7643;
  assign tmp7638 = s2 ? tmp7639 : tmp7641;
  assign tmp7646 = s0 ? 1 : tmp7595;
  assign tmp7647 = s0 ? tmp6997 : tmp7596;
  assign tmp7645 = s1 ? tmp7646 : tmp7647;
  assign tmp7644 = ~(s2 ? tmp7645 : tmp7016);
  assign tmp7637 = s3 ? tmp7638 : tmp7644;
  assign tmp7624 = s4 ? tmp7625 : tmp7637;
  assign tmp7623 = s5 ? tmp7577 : tmp7624;
  assign tmp7622 = s6 ? tmp7623 : tmp7576;
  assign tmp7648 = ~(s6 ? tmp7048 : tmp7600);
  assign tmp7621 = ~(s7 ? tmp7622 : tmp7648);
  assign tmp7597 = ~(s8 ? tmp7598 : tmp7621);
  assign tmp7575 = s9 ? tmp7576 : tmp7597;
  assign tmp7652 = ~(s6 ? tmp6923 : tmp7600);
  assign tmp7651 = ~(s7 ? tmp7622 : tmp7652);
  assign tmp7650 = ~(s8 ? tmp7598 : tmp7651);
  assign tmp7649 = s9 ? tmp7576 : tmp7650;
  assign tmp7574 = s10 ? tmp7575 : tmp7649;
  assign tmp7661 = s0 ? tmp7603 : tmp7358;
  assign tmp7662 = s0 ? tmp7089 : tmp7603;
  assign tmp7660 = s1 ? tmp7661 : tmp7662;
  assign tmp7659 = s2 ? tmp7603 : tmp7660;
  assign tmp7666 = s1 ? tmp7603 : tmp7032;
  assign tmp7668 = s0 ? tmp7603 : tmp7113;
  assign tmp7667 = s1 ? tmp7603 : tmp7668;
  assign tmp7665 = s2 ? tmp7666 : tmp7667;
  assign tmp7670 = s1 ? tmp7122 : tmp6926;
  assign tmp7669 = s2 ? tmp7670 : tmp7614;
  assign tmp7664 = s3 ? tmp7665 : tmp7669;
  assign tmp7673 = ~(s1 ? tmp7603 : tmp7128);
  assign tmp7672 = s2 ? tmp7099 : tmp7673;
  assign tmp7674 = ~(s1 ? tmp7595 : tmp7603);
  assign tmp7671 = ~(s3 ? tmp7672 : tmp7674);
  assign tmp7663 = s4 ? tmp7664 : tmp7671;
  assign tmp7658 = s5 ? tmp7659 : tmp7663;
  assign tmp7657 = s6 ? tmp7658 : tmp6966;
  assign tmp7656 = s7 ? tmp7104 : tmp7657;
  assign tmp7677 = ~(s5 ? tmp7659 : tmp7663);
  assign tmp7676 = s6 ? tmp7137 : tmp7677;
  assign tmp7675 = ~(s7 ? tmp7622 : tmp7676);
  assign tmp7655 = ~(s8 ? tmp7656 : tmp7675);
  assign tmp7654 = s9 ? tmp7576 : tmp7655;
  assign tmp7681 = s6 ? tmp7075 : tmp7677;
  assign tmp7680 = ~(s7 ? tmp7622 : tmp7681);
  assign tmp7679 = ~(s8 ? tmp7656 : tmp7680);
  assign tmp7678 = s9 ? tmp7576 : tmp7679;
  assign tmp7653 = s10 ? tmp7654 : tmp7678;
  assign tmp7573 = s11 ? tmp7574 : tmp7653;
  assign tmp7686 = s7 ? tmp7177 : tmp7599;
  assign tmp7688 = ~(s6 ? tmp7203 : tmp7600);
  assign tmp7687 = ~(s7 ? tmp7622 : tmp7688);
  assign tmp7685 = ~(s8 ? tmp7686 : tmp7687);
  assign tmp7684 = s9 ? tmp7576 : tmp7685;
  assign tmp7692 = ~(s6 ? tmp7146 : tmp7600);
  assign tmp7691 = ~(s7 ? tmp7622 : tmp7692);
  assign tmp7690 = ~(s8 ? tmp7686 : tmp7691);
  assign tmp7689 = s9 ? tmp7576 : tmp7690;
  assign tmp7683 = s10 ? tmp7684 : tmp7689;
  assign tmp7698 = l1 ? tmp6927 : tmp6957;
  assign tmp7699 = l1 ? tmp6926 : tmp6957;
  assign tmp7697 = s1 ? tmp7698 : tmp7699;
  assign tmp7702 = l1 ? tmp6927 : tmp6983;
  assign tmp7701 = s0 ? tmp7699 : tmp7702;
  assign tmp7703 = s0 ? tmp6998 : tmp7699;
  assign tmp7700 = s1 ? tmp7701 : tmp7703;
  assign tmp7696 = s2 ? tmp7697 : tmp7700;
  assign tmp7707 = s1 ? tmp7703 : tmp6983;
  assign tmp7709 = s0 ? tmp7699 : 1;
  assign tmp7708 = s1 ? tmp7698 : tmp7709;
  assign tmp7706 = s2 ? tmp7707 : tmp7708;
  assign tmp7711 = s1 ? tmp7042 : tmp6951;
  assign tmp7712 = s1 ? tmp6946 : tmp7590;
  assign tmp7710 = ~(s2 ? tmp7711 : tmp7712);
  assign tmp7705 = s3 ? tmp7706 : tmp7710;
  assign tmp7715 = s1 ? tmp6955 : tmp7356;
  assign tmp7717 = l1 ? tmp6926 : tmp6955;
  assign tmp7716 = s1 ? tmp7699 : tmp7717;
  assign tmp7714 = s2 ? tmp7715 : tmp7716;
  assign tmp7719 = l1 ? tmp6957 : tmp6928;
  assign tmp7720 = ~(l1 ? tmp6926 : tmp6957);
  assign tmp7718 = ~(s1 ? tmp7719 : tmp7720);
  assign tmp7713 = s3 ? tmp7714 : tmp7718;
  assign tmp7704 = s4 ? tmp7705 : tmp7713;
  assign tmp7695 = s5 ? tmp7696 : tmp7704;
  assign tmp7727 = l1 ? tmp6947 : tmp6984;
  assign tmp7728 = l1 ? tmp6957 : tmp6984;
  assign tmp7726 = s1 ? tmp7727 : tmp7728;
  assign tmp7730 = s0 ? tmp7728 : tmp6946;
  assign tmp7731 = s0 ? tmp7089 : tmp7728;
  assign tmp7729 = s1 ? tmp7730 : tmp7731;
  assign tmp7725 = s2 ? tmp7726 : tmp7729;
  assign tmp7735 = s1 ? tmp7731 : tmp7032;
  assign tmp7737 = s0 ? tmp7728 : tmp7113;
  assign tmp7736 = s1 ? tmp7727 : tmp7737;
  assign tmp7734 = s2 ? tmp7735 : tmp7736;
  assign tmp7739 = s1 ? tmp6960 : tmp6951;
  assign tmp7740 = s1 ? tmp6946 : tmp7615;
  assign tmp7738 = s2 ? tmp7739 : tmp7740;
  assign tmp7733 = s3 ? tmp7734 : tmp7738;
  assign tmp7743 = s1 ? 1 : tmp7356;
  assign tmp7745 = ~(l1 ? tmp6926 : 1);
  assign tmp7744 = ~(s1 ? tmp7728 : tmp7745);
  assign tmp7742 = s2 ? tmp7743 : tmp7744;
  assign tmp7746 = ~(s1 ? tmp7719 : tmp7728);
  assign tmp7741 = ~(s3 ? tmp7742 : tmp7746);
  assign tmp7732 = s4 ? tmp7733 : tmp7741;
  assign tmp7724 = s5 ? tmp7725 : tmp7732;
  assign tmp7723 = s6 ? tmp7724 : tmp6966;
  assign tmp7722 = s7 ? tmp7275 : tmp7723;
  assign tmp7749 = ~(s5 ? tmp7696 : tmp7704);
  assign tmp7748 = s6 ? tmp6966 : tmp7749;
  assign tmp7750 = s6 ? tmp7303 : tmp7724;
  assign tmp7747 = s7 ? tmp7748 : tmp7750;
  assign tmp7721 = ~(s8 ? tmp7722 : tmp7747);
  assign tmp7694 = s9 ? tmp7695 : tmp7721;
  assign tmp7754 = s6 ? tmp7241 : tmp7724;
  assign tmp7753 = s7 ? tmp7748 : tmp7754;
  assign tmp7752 = ~(s8 ? tmp7722 : tmp7753);
  assign tmp7751 = s9 ? tmp7695 : tmp7752;
  assign tmp7693 = s10 ? tmp7694 : tmp7751;
  assign tmp7682 = s11 ? tmp7683 : tmp7693;
  assign tmp7572 = s12 ? tmp7573 : tmp7682;
  assign tmp7760 = s7 ? tmp7371 : tmp7599;
  assign tmp7763 = ~(s5 ? tmp7601 : tmp7606);
  assign tmp7762 = s6 ? tmp7402 : tmp7763;
  assign tmp7761 = ~(s7 ? tmp7622 : tmp7762);
  assign tmp7759 = ~(s8 ? tmp7760 : tmp7761);
  assign tmp7758 = s9 ? tmp7576 : tmp7759;
  assign tmp7767 = s6 ? tmp7342 : tmp7763;
  assign tmp7766 = ~(s7 ? tmp7622 : tmp7767);
  assign tmp7765 = ~(s8 ? tmp7760 : tmp7766);
  assign tmp7764 = s9 ? tmp7576 : tmp7765;
  assign tmp7757 = s10 ? tmp7758 : tmp7764;
  assign tmp7756 = s11 ? tmp7757 : tmp7574;
  assign tmp7772 = s7 ? tmp7443 : tmp7723;
  assign tmp7775 = s5 ? tmp7413 : tmp7474;
  assign tmp7776 = ~(s5 ? tmp7725 : tmp7732);
  assign tmp7774 = ~(s6 ? tmp7775 : tmp7776);
  assign tmp7773 = s7 ? tmp7748 : tmp7774;
  assign tmp7771 = ~(s8 ? tmp7772 : tmp7773);
  assign tmp7770 = s9 ? tmp7695 : tmp7771;
  assign tmp7780 = ~(s6 ? tmp7412 : tmp7776);
  assign tmp7779 = s7 ? tmp7748 : tmp7780;
  assign tmp7778 = ~(s8 ? tmp7772 : tmp7779);
  assign tmp7777 = s9 ? tmp7695 : tmp7778;
  assign tmp7769 = s10 ? tmp7770 : tmp7777;
  assign tmp7784 = s7 ? tmp7537 : tmp7723;
  assign tmp7786 = s6 ? tmp7555 : tmp7724;
  assign tmp7785 = s7 ? tmp7748 : tmp7786;
  assign tmp7783 = ~(s8 ? tmp7784 : tmp7785);
  assign tmp7782 = s9 ? tmp7695 : tmp7783;
  assign tmp7790 = s6 ? tmp7506 : tmp7724;
  assign tmp7789 = s7 ? tmp7748 : tmp7790;
  assign tmp7788 = ~(s8 ? tmp7784 : tmp7789);
  assign tmp7787 = s9 ? tmp7695 : tmp7788;
  assign tmp7781 = s10 ? tmp7782 : tmp7787;
  assign tmp7768 = s11 ? tmp7769 : tmp7781;
  assign tmp7755 = s12 ? tmp7756 : tmp7768;
  assign tmp7571 = s13 ? tmp7572 : tmp7755;
  assign tmp7803 = s1 ? tmp6945 : tmp6970;
  assign tmp7802 = ~(s2 ? tmp7803 : tmp7060);
  assign tmp7801 = s3 ? tmp7030 : tmp7802;
  assign tmp7804 = ~(s3 ? tmp7068 : tmp7045);
  assign tmp7800 = s4 ? tmp7801 : tmp7804;
  assign tmp7799 = s5 ? tmp7022 : tmp7800;
  assign tmp7798 = s6 ? tmp7799 : tmp6966;
  assign tmp7797 = s7 ? tmp6965 : tmp7798;
  assign tmp7808 = s4 ? tmp7801 : tmp7039;
  assign tmp7807 = s5 ? tmp7022 : tmp7808;
  assign tmp7806 = s6 ? tmp7056 : tmp7807;
  assign tmp7805 = s7 ? tmp7047 : tmp7806;
  assign tmp7796 = s8 ? tmp7797 : tmp7805;
  assign tmp7795 = s9 ? tmp6923 : tmp7796;
  assign tmp7812 = s6 ? tmp7065 : tmp7799;
  assign tmp7811 = s7 ? tmp6965 : tmp7812;
  assign tmp7810 = s8 ? tmp7797 : tmp7811;
  assign tmp7809 = s9 ? tmp6923 : tmp7810;
  assign tmp7794 = s10 ? tmp7795 : tmp7809;
  assign tmp7822 = s1 ? tmp7109 : tmp6981;
  assign tmp7824 = s0 ? tmp7109 : tmp6982;
  assign tmp7823 = s1 ? tmp7824 : tmp7119;
  assign tmp7821 = s2 ? tmp7822 : tmp7823;
  assign tmp7820 = s3 ? tmp7821 : tmp7120;
  assign tmp7819 = s4 ? tmp7820 : tmp7125;
  assign tmp7818 = s5 ? tmp7108 : tmp7819;
  assign tmp7817 = s6 ? tmp7818 : tmp6966;
  assign tmp7816 = s7 ? tmp7104 : tmp7817;
  assign tmp7830 = s2 ? tmp7822 : tmp7118;
  assign tmp7829 = s3 ? tmp7830 : tmp7120;
  assign tmp7828 = s4 ? tmp7829 : tmp7125;
  assign tmp7827 = ~(s5 ? tmp7108 : tmp7828);
  assign tmp7826 = ~(s6 ? tmp7137 : tmp7827);
  assign tmp7825 = s7 ? tmp7131 : tmp7826;
  assign tmp7815 = ~(s8 ? tmp7816 : tmp7825);
  assign tmp7814 = s9 ? tmp7075 : tmp7815;
  assign tmp7835 = ~(s5 ? tmp7108 : tmp7819);
  assign tmp7834 = ~(s6 ? tmp7075 : tmp7835);
  assign tmp7833 = s7 ? tmp7104 : tmp7834;
  assign tmp7832 = ~(s8 ? tmp7816 : tmp7833);
  assign tmp7831 = s9 ? tmp7075 : tmp7832;
  assign tmp7813 = ~(s10 ? tmp7814 : tmp7831);
  assign tmp7793 = s11 ? tmp7794 : tmp7813;
  assign tmp7846 = s1 ? tmp7002 : tmp7196;
  assign tmp7845 = s2 ? tmp7846 : tmp7197;
  assign tmp7848 = s1 ? tmp7200 : tmp6976;
  assign tmp7849 = ~(l1 ? tmp6983 : tmp7004);
  assign tmp7847 = ~(s2 ? tmp7848 : tmp7849);
  assign tmp7844 = ~(s3 ? tmp7845 : tmp7847);
  assign tmp7843 = s4 ? tmp7185 : tmp7844;
  assign tmp7842 = s5 ? tmp7180 : tmp7843;
  assign tmp7841 = s6 ? tmp7842 : tmp6966;
  assign tmp7840 = s7 ? tmp7177 : tmp7841;
  assign tmp7854 = ~(s3 ? tmp7845 : tmp7199);
  assign tmp7853 = s4 ? tmp7185 : tmp7854;
  assign tmp7852 = s5 ? tmp7180 : tmp7853;
  assign tmp7851 = s6 ? tmp7214 : tmp7852;
  assign tmp7850 = s7 ? tmp7202 : tmp7851;
  assign tmp7839 = s8 ? tmp7840 : tmp7850;
  assign tmp7838 = s9 ? tmp7146 : tmp7839;
  assign tmp7858 = s6 ? tmp7227 : tmp7842;
  assign tmp7857 = s7 ? tmp7177 : tmp7858;
  assign tmp7856 = s8 ? tmp7840 : tmp7857;
  assign tmp7855 = s9 ? tmp7146 : tmp7856;
  assign tmp7837 = s10 ? tmp7838 : tmp7855;
  assign tmp7868 = s1 ? tmp6974 : tmp7321;
  assign tmp7867 = s2 ? tmp7292 : tmp7868;
  assign tmp7866 = s3 ? tmp7287 : tmp7867;
  assign tmp7870 = ~(s1 ? tmp7245 : tmp7337);
  assign tmp7869 = ~(s3 ? tmp7296 : tmp7870);
  assign tmp7865 = s4 ? tmp7866 : tmp7869;
  assign tmp7864 = s5 ? tmp7278 : tmp7865;
  assign tmp7863 = s6 ? tmp7864 : tmp6966;
  assign tmp7862 = s7 ? tmp7275 : tmp7863;
  assign tmp7874 = s4 ? tmp7866 : tmp7295;
  assign tmp7873 = s5 ? tmp7278 : tmp7874;
  assign tmp7872 = s6 ? tmp7314 : tmp7873;
  assign tmp7871 = s7 ? tmp7302 : tmp7872;
  assign tmp7861 = s8 ? tmp7862 : tmp7871;
  assign tmp7860 = s9 ? tmp7241 : tmp7861;
  assign tmp7878 = s6 ? tmp7326 : tmp7864;
  assign tmp7877 = s7 ? tmp7275 : tmp7878;
  assign tmp7876 = s8 ? tmp7862 : tmp7877;
  assign tmp7875 = s9 ? tmp7241 : tmp7876;
  assign tmp7859 = s10 ? tmp7860 : tmp7875;
  assign tmp7836 = s11 ? tmp7837 : tmp7859;
  assign tmp7792 = s12 ? tmp7793 : tmp7836;
  assign tmp7891 = s0 ? tmp6955 : tmp6951;
  assign tmp7890 = s1 ? tmp6951 : tmp7891;
  assign tmp7889 = s2 ? tmp7890 : tmp7391;
  assign tmp7893 = s1 ? tmp7394 : tmp7003;
  assign tmp7892 = ~(s2 ? tmp7893 : tmp6948);
  assign tmp7888 = ~(s3 ? tmp7889 : tmp7892);
  assign tmp7887 = s4 ? tmp7381 : tmp7888;
  assign tmp7886 = s5 ? tmp7375 : tmp7887;
  assign tmp7885 = s6 ? tmp7886 : tmp6966;
  assign tmp7884 = s7 ? tmp7371 : tmp7885;
  assign tmp7898 = ~(s3 ? tmp7889 : tmp7393);
  assign tmp7897 = s4 ? tmp7381 : tmp7898;
  assign tmp7896 = ~(s5 ? tmp7375 : tmp7897);
  assign tmp7895 = ~(s6 ? tmp7402 : tmp7896);
  assign tmp7894 = s7 ? tmp7396 : tmp7895;
  assign tmp7883 = ~(s8 ? tmp7884 : tmp7894);
  assign tmp7882 = s9 ? tmp7342 : tmp7883;
  assign tmp7903 = ~(s5 ? tmp7375 : tmp7887);
  assign tmp7902 = ~(s6 ? tmp7342 : tmp7903);
  assign tmp7901 = s7 ? tmp7371 : tmp7902;
  assign tmp7900 = ~(s8 ? tmp7884 : tmp7901);
  assign tmp7899 = s9 ? tmp7342 : tmp7900;
  assign tmp7881 = s10 ? tmp7882 : tmp7899;
  assign tmp7914 = s0 ? 1 : tmp6926;
  assign tmp7913 = s1 ? tmp6955 : tmp7914;
  assign tmp7912 = s2 ? tmp7913 : tmp7037;
  assign tmp7911 = s3 ? tmp7030 : tmp7912;
  assign tmp7915 = ~(s3 ? tmp7040 : tmp7071);
  assign tmp7910 = s4 ? tmp7911 : tmp7915;
  assign tmp7909 = s5 ? tmp7022 : tmp7910;
  assign tmp7908 = s6 ? tmp7909 : tmp6966;
  assign tmp7907 = s7 ? tmp6965 : tmp7908;
  assign tmp7919 = s4 ? tmp7911 : tmp7039;
  assign tmp7918 = s5 ? tmp7022 : tmp7919;
  assign tmp7917 = s6 ? tmp7056 : tmp7918;
  assign tmp7916 = s7 ? tmp7047 : tmp7917;
  assign tmp7906 = s8 ? tmp7907 : tmp7916;
  assign tmp7905 = s9 ? tmp6923 : tmp7906;
  assign tmp7923 = s6 ? tmp7065 : tmp7909;
  assign tmp7922 = s7 ? tmp6965 : tmp7923;
  assign tmp7921 = s8 ? tmp7907 : tmp7922;
  assign tmp7920 = s9 ? tmp6923 : tmp7921;
  assign tmp7904 = ~(s10 ? tmp7905 : tmp7920);
  assign tmp7880 = s11 ? tmp7881 : tmp7904;
  assign tmp7933 = s2 ? tmp7549 : tmp7559;
  assign tmp7935 = s1 ? tmp7533 : tmp7510;
  assign tmp7934 = ~(s2 ? tmp7935 : tmp7019);
  assign tmp7932 = ~(s3 ? tmp7933 : tmp7934);
  assign tmp7931 = s4 ? tmp7541 : tmp7932;
  assign tmp7930 = s5 ? tmp7507 : tmp7931;
  assign tmp7929 = s6 ? tmp7930 : tmp6966;
  assign tmp7928 = s7 ? tmp7537 : tmp7929;
  assign tmp7940 = ~(s3 ? tmp7933 : tmp7552);
  assign tmp7939 = s4 ? tmp7541 : tmp7940;
  assign tmp7938 = s5 ? tmp7507 : tmp7939;
  assign tmp7937 = s6 ? tmp7561 : tmp7938;
  assign tmp7936 = s7 ? tmp7554 : tmp7937;
  assign tmp7927 = s8 ? tmp7928 : tmp7936;
  assign tmp7926 = s9 ? tmp7506 : tmp7927;
  assign tmp7944 = s6 ? tmp7568 : tmp7930;
  assign tmp7943 = s7 ? tmp7537 : tmp7944;
  assign tmp7942 = s8 ? tmp7928 : tmp7943;
  assign tmp7941 = s9 ? tmp7506 : tmp7942;
  assign tmp7925 = ~(s10 ? tmp7926 : tmp7941);
  assign tmp7924 = s11 ? tmp7410 : tmp7925;
  assign tmp7879 = ~(s12 ? tmp7880 : tmp7924);
  assign tmp7791 = ~(s13 ? tmp7792 : tmp7879);
  assign tmp7570 = ~(s15 ? tmp7571 : tmp7791);
  assign tmp6917 = s16 ? tmp6918 : tmp7570;
  assign s1n = tmp6917;

  assign tmp7956 = l3 ? 1 : 0;
  assign tmp7955 = l2 ? 1 : tmp7956;
  assign tmp7957 = l2 ? tmp7956 : 0;
  assign tmp7954 = l1 ? tmp7955 : tmp7957;
  assign tmp7958 = l1 ? tmp7956 : tmp7957;
  assign tmp7953 = s1 ? tmp7954 : tmp7958;
  assign tmp7961 = l1 ? 1 : tmp7957;
  assign tmp7960 = s0 ? tmp7961 : tmp7958;
  assign tmp7959 = s1 ? tmp7958 : tmp7960;
  assign tmp7952 = s2 ? tmp7953 : tmp7959;
  assign tmp7967 = l1 ? tmp7955 : 0;
  assign tmp7966 = s0 ? tmp7967 : tmp7958;
  assign tmp7969 = ~(l2 ? tmp7956 : 0);
  assign tmp7968 = ~(l1 ? 1 : tmp7969);
  assign tmp7965 = s1 ? tmp7966 : tmp7968;
  assign tmp7972 = l1 ? 1 : tmp7969;
  assign tmp7971 = s0 ? tmp7958 : tmp7972;
  assign tmp7970 = s1 ? tmp7954 : tmp7971;
  assign tmp7964 = s2 ? tmp7965 : tmp7970;
  assign tmp7975 = s0 ? tmp7972 : 1;
  assign tmp7978 = l2 ? tmp7956 : 1;
  assign tmp7977 = l1 ? tmp7978 : 1;
  assign tmp7976 = s0 ? tmp7977 : 0;
  assign tmp7974 = s1 ? tmp7975 : tmp7976;
  assign tmp7982 = ~(l3 ? 1 : 0);
  assign tmp7981 = l2 ? 1 : tmp7982;
  assign tmp7980 = l1 ? tmp7955 : tmp7981;
  assign tmp7983 = l1 ? tmp7956 : 0;
  assign tmp7979 = s1 ? tmp7980 : tmp7983;
  assign tmp7973 = s2 ? tmp7974 : tmp7979;
  assign tmp7963 = s3 ? tmp7964 : tmp7973;
  assign tmp7987 = l1 ? tmp7981 : 1;
  assign tmp7986 = s1 ? 1 : tmp7987;
  assign tmp7990 = ~(l1 ? tmp7981 : 1);
  assign tmp7989 = s0 ? tmp7972 : tmp7990;
  assign tmp7988 = ~(s1 ? tmp7958 : tmp7989);
  assign tmp7985 = s2 ? tmp7986 : tmp7988;
  assign tmp7993 = ~(l1 ? tmp7981 : tmp7969);
  assign tmp7992 = s0 ? tmp7977 : tmp7993;
  assign tmp7991 = ~(s1 ? tmp7992 : tmp7958);
  assign tmp7984 = ~(s3 ? tmp7985 : tmp7991);
  assign tmp7962 = s4 ? tmp7963 : tmp7984;
  assign tmp7951 = s5 ? tmp7952 : tmp7962;
  assign tmp8002 = ~(l2 ? 1 : tmp7982);
  assign tmp8001 = l1 ? tmp7978 : tmp8002;
  assign tmp8000 = s0 ? tmp7972 : tmp8001;
  assign tmp7999 = s1 ? tmp8000 : tmp7975;
  assign tmp7998 = s2 ? tmp7972 : tmp7999;
  assign tmp8008 = l1 ? tmp7955 : tmp7969;
  assign tmp8007 = s0 ? tmp8008 : tmp7972;
  assign tmp8009 = l1 ? tmp7957 : tmp8002;
  assign tmp8006 = s1 ? tmp8007 : tmp8009;
  assign tmp8011 = s0 ? tmp7972 : tmp8009;
  assign tmp8010 = s1 ? tmp8011 : tmp7972;
  assign tmp8005 = s2 ? tmp8006 : tmp8010;
  assign tmp8016 = l2 ? 1 : 0;
  assign tmp8015 = ~(l1 ? tmp7955 : tmp8016);
  assign tmp8014 = s0 ? tmp7977 : tmp8015;
  assign tmp8013 = s1 ? tmp7975 : tmp8014;
  assign tmp8018 = s0 ? tmp7980 : tmp7968;
  assign tmp8020 = l1 ? tmp7956 : tmp7969;
  assign tmp8019 = ~(s0 ? tmp7972 : tmp8020);
  assign tmp8017 = ~(s1 ? tmp8018 : tmp8019);
  assign tmp8012 = s2 ? tmp8013 : tmp8017;
  assign tmp8004 = s3 ? tmp8005 : tmp8012;
  assign tmp8026 = ~(l2 ? tmp7956 : tmp7982);
  assign tmp8025 = l1 ? tmp7956 : tmp8026;
  assign tmp8027 = ~(l1 ? tmp7978 : tmp7956);
  assign tmp8024 = s0 ? tmp8025 : tmp8027;
  assign tmp8029 = l1 ? 1 : tmp7978;
  assign tmp8030 = l1 ? tmp7957 : tmp7955;
  assign tmp8028 = ~(s0 ? tmp8029 : tmp8030);
  assign tmp8023 = s1 ? tmp8024 : tmp8028;
  assign tmp8033 = l1 ? tmp8016 : 1;
  assign tmp8032 = s0 ? tmp8033 : tmp7968;
  assign tmp8035 = ~(l1 ? tmp7957 : tmp7956);
  assign tmp8034 = ~(s0 ? tmp7972 : tmp8035);
  assign tmp8031 = ~(s1 ? tmp8032 : tmp8034);
  assign tmp8022 = s2 ? tmp8023 : tmp8031;
  assign tmp8039 = ~(l1 ? tmp7957 : tmp8016);
  assign tmp8038 = s0 ? tmp7977 : tmp8039;
  assign tmp8037 = s1 ? tmp8038 : tmp7975;
  assign tmp8042 = ~(l1 ? 1 : tmp7978);
  assign tmp8041 = s0 ? tmp8025 : tmp8042;
  assign tmp8043 = ~(s0 ? tmp7980 : tmp8033);
  assign tmp8040 = s1 ? tmp8041 : tmp8043;
  assign tmp8036 = s2 ? tmp8037 : tmp8040;
  assign tmp8021 = s3 ? tmp8022 : tmp8036;
  assign tmp8003 = s4 ? tmp8004 : tmp8021;
  assign tmp7997 = s5 ? tmp7998 : tmp8003;
  assign tmp7996 = s6 ? tmp7997 : tmp7951;
  assign tmp8048 = ~(l2 ? tmp7956 : 1);
  assign tmp8047 = l1 ? tmp7955 : tmp8048;
  assign tmp8050 = s0 ? tmp8047 : tmp7983;
  assign tmp8052 = l1 ? 1 : tmp8048;
  assign tmp8053 = l1 ? tmp7955 : tmp8016;
  assign tmp8051 = s0 ? tmp8052 : tmp8053;
  assign tmp8049 = s1 ? tmp8050 : tmp8051;
  assign tmp8046 = s2 ? tmp8047 : tmp8049;
  assign tmp8058 = l1 ? tmp7957 : 0;
  assign tmp8057 = s1 ? tmp8047 : tmp8058;
  assign tmp8060 = s0 ? tmp8047 : tmp7972;
  assign tmp8059 = s1 ? tmp8047 : tmp8060;
  assign tmp8056 = s2 ? tmp8057 : tmp8059;
  assign tmp8062 = s1 ? 1 : 0;
  assign tmp8064 = l1 ? tmp7955 : tmp7982;
  assign tmp8065 = l1 ? tmp7956 : tmp8048;
  assign tmp8063 = s1 ? tmp8064 : tmp8065;
  assign tmp8061 = s2 ? tmp8062 : tmp8063;
  assign tmp8055 = s3 ? tmp8056 : tmp8061;
  assign tmp8070 = l2 ? tmp7956 : tmp7982;
  assign tmp8069 = l1 ? tmp8070 : 1;
  assign tmp8068 = s1 ? tmp7978 : tmp8069;
  assign tmp8072 = ~(l1 ? tmp8070 : tmp7978);
  assign tmp8071 = ~(s1 ? tmp8047 : tmp8072);
  assign tmp8067 = s2 ? tmp8068 : tmp8071;
  assign tmp8073 = s1 ? tmp8069 : tmp8015;
  assign tmp8066 = ~(s3 ? tmp8067 : tmp8073);
  assign tmp8054 = s4 ? tmp8055 : tmp8066;
  assign tmp8045 = s5 ? tmp8046 : tmp8054;
  assign tmp8044 = s6 ? tmp8045 : tmp7997;
  assign tmp7995 = s7 ? tmp7996 : tmp8044;
  assign tmp8080 = ~(s1 ? tmp7958 : tmp7990);
  assign tmp8079 = s2 ? tmp7986 : tmp8080;
  assign tmp8082 = l1 ? tmp7981 : tmp7969;
  assign tmp8083 = ~(l1 ? tmp7956 : tmp7957);
  assign tmp8081 = s1 ? tmp8082 : tmp8083;
  assign tmp8078 = ~(s3 ? tmp8079 : tmp8081);
  assign tmp8077 = s4 ? tmp7963 : tmp8078;
  assign tmp8076 = s5 ? tmp7952 : tmp8077;
  assign tmp8075 = s6 ? tmp7997 : tmp8076;
  assign tmp8088 = s2 ? tmp7974 : tmp8063;
  assign tmp8087 = s3 ? tmp8056 : tmp8088;
  assign tmp8086 = s4 ? tmp8087 : tmp8066;
  assign tmp8085 = s5 ? tmp8046 : tmp8086;
  assign tmp8084 = s6 ? tmp8085 : tmp8045;
  assign tmp8074 = s7 ? tmp8075 : tmp8084;
  assign tmp7994 = s8 ? tmp7995 : tmp8074;
  assign tmp7950 = s9 ? tmp7951 : tmp7994;
  assign tmp8098 = s0 ? tmp7972 : tmp8072;
  assign tmp8097 = ~(s1 ? tmp8047 : tmp8098);
  assign tmp8096 = s2 ? tmp8068 : tmp8097;
  assign tmp8101 = ~(l1 ? tmp8070 : 1);
  assign tmp8100 = s0 ? tmp7977 : tmp8101;
  assign tmp8099 = ~(s1 ? tmp8100 : tmp8053);
  assign tmp8095 = ~(s3 ? tmp8096 : tmp8099);
  assign tmp8094 = s4 ? tmp8087 : tmp8095;
  assign tmp8093 = s5 ? tmp8046 : tmp8094;
  assign tmp8092 = s6 ? tmp8093 : tmp8045;
  assign tmp8091 = s7 ? tmp7996 : tmp8092;
  assign tmp8090 = s8 ? tmp7995 : tmp8091;
  assign tmp8089 = s9 ? tmp7951 : tmp8090;
  assign tmp7949 = s10 ? tmp7950 : tmp8089;
  assign tmp8107 = l1 ? tmp7978 : tmp7981;
  assign tmp8108 = l1 ? 1 : tmp7981;
  assign tmp8106 = s1 ? tmp8107 : tmp8108;
  assign tmp8111 = l1 ? tmp7956 : tmp7981;
  assign tmp8112 = l1 ? 1 : tmp7982;
  assign tmp8110 = s0 ? tmp8111 : tmp8112;
  assign tmp8109 = s1 ? tmp8108 : tmp8110;
  assign tmp8105 = s2 ? tmp8106 : tmp8109;
  assign tmp8117 = ~(l1 ? tmp7957 : tmp8002);
  assign tmp8116 = s1 ? tmp8108 : tmp8117;
  assign tmp8119 = s0 ? tmp8107 : tmp8117;
  assign tmp8120 = s0 ? tmp8108 : tmp7983;
  assign tmp8118 = s1 ? tmp8119 : tmp8120;
  assign tmp8115 = s2 ? tmp8116 : tmp8118;
  assign tmp8123 = l1 ? tmp8070 : tmp7978;
  assign tmp8124 = ~(l1 ? 1 : tmp7981);
  assign tmp8122 = s1 ? tmp8123 : tmp8124;
  assign tmp8126 = l1 ? tmp8016 : tmp7969;
  assign tmp8125 = s1 ? tmp8126 : tmp8124;
  assign tmp8121 = ~(s2 ? tmp8122 : tmp8125);
  assign tmp8114 = s3 ? tmp8115 : tmp8121;
  assign tmp8129 = s1 ? tmp8108 : 1;
  assign tmp8128 = s2 ? 1 : tmp8129;
  assign tmp8130 = s1 ? tmp8108 : tmp8112;
  assign tmp8127 = s3 ? tmp8128 : tmp8130;
  assign tmp8113 = s4 ? tmp8114 : tmp8127;
  assign tmp8104 = s5 ? tmp8105 : tmp8113;
  assign tmp8134 = ~(s5 ? tmp8105 : tmp8113);
  assign tmp8133 = s6 ? tmp7997 : tmp8134;
  assign tmp8139 = l1 ? tmp8016 : tmp8026;
  assign tmp8140 = l1 ? tmp7957 : tmp8026;
  assign tmp8138 = s1 ? tmp8139 : tmp8140;
  assign tmp8142 = s0 ? tmp8140 : tmp8009;
  assign tmp8144 = l1 ? tmp7981 : tmp8026;
  assign tmp8143 = s0 ? tmp8144 : tmp8030;
  assign tmp8141 = s1 ? tmp8142 : tmp8143;
  assign tmp8137 = s2 ? tmp8138 : tmp8141;
  assign tmp8148 = s1 ? tmp8140 : tmp8009;
  assign tmp8150 = s0 ? tmp8140 : tmp8082;
  assign tmp8149 = s1 ? tmp8139 : tmp8150;
  assign tmp8147 = s2 ? tmp8148 : tmp8149;
  assign tmp8152 = s1 ? tmp8069 : tmp8124;
  assign tmp8153 = s1 ? tmp8126 : tmp8140;
  assign tmp8151 = s2 ? tmp8152 : tmp8153;
  assign tmp8146 = s3 ? tmp8147 : tmp8151;
  assign tmp8156 = s1 ? tmp8029 : 1;
  assign tmp8157 = ~(s1 ? tmp8140 : tmp8042);
  assign tmp8155 = s2 ? tmp8156 : tmp8157;
  assign tmp8159 = ~(l1 ? tmp7957 : tmp7955);
  assign tmp8158 = s1 ? tmp8108 : tmp8159;
  assign tmp8154 = ~(s3 ? tmp8155 : tmp8158);
  assign tmp8145 = s4 ? tmp8146 : tmp8154;
  assign tmp8136 = s5 ? tmp8137 : tmp8145;
  assign tmp8135 = s6 ? tmp8136 : tmp7997;
  assign tmp8132 = s7 ? tmp8133 : tmp8135;
  assign tmp8166 = s1 ? tmp8107 : tmp8120;
  assign tmp8165 = s2 ? tmp8116 : tmp8166;
  assign tmp8164 = s3 ? tmp8165 : tmp8121;
  assign tmp8163 = s4 ? tmp8164 : tmp8127;
  assign tmp8162 = ~(s5 ? tmp8105 : tmp8163);
  assign tmp8161 = s6 ? tmp7997 : tmp8162;
  assign tmp8168 = s5 ? tmp8105 : tmp8163;
  assign tmp8169 = ~(s5 ? tmp8137 : tmp8145);
  assign tmp8167 = ~(s6 ? tmp8168 : tmp8169);
  assign tmp8160 = s7 ? tmp8161 : tmp8167;
  assign tmp8131 = ~(s8 ? tmp8132 : tmp8160);
  assign tmp8103 = s9 ? tmp8104 : tmp8131;
  assign tmp8173 = ~(s6 ? tmp8104 : tmp8169);
  assign tmp8172 = s7 ? tmp8133 : tmp8173;
  assign tmp8171 = ~(s8 ? tmp8132 : tmp8172);
  assign tmp8170 = s9 ? tmp8104 : tmp8171;
  assign tmp8102 = ~(s10 ? tmp8103 : tmp8170);
  assign tmp7948 = s11 ? tmp7949 : tmp8102;
  assign tmp8179 = s1 ? tmp8008 : tmp8020;
  assign tmp8182 = l1 ? tmp7956 : tmp8002;
  assign tmp8181 = s0 ? tmp8020 : tmp8182;
  assign tmp8184 = l1 ? tmp7956 : 1;
  assign tmp8183 = s0 ? tmp7972 : tmp8184;
  assign tmp8180 = s1 ? tmp8181 : tmp8183;
  assign tmp8178 = s2 ? tmp8179 : tmp8180;
  assign tmp8189 = s0 ? tmp8008 : tmp8020;
  assign tmp8188 = s1 ? tmp8189 : tmp8009;
  assign tmp8191 = s0 ? tmp8008 : tmp8009;
  assign tmp8192 = s0 ? tmp8020 : tmp7972;
  assign tmp8190 = s1 ? tmp8191 : tmp8192;
  assign tmp8187 = s2 ? tmp8188 : tmp8190;
  assign tmp8196 = ~(l1 ? 1 : tmp8016);
  assign tmp8195 = s0 ? tmp7977 : tmp8196;
  assign tmp8194 = s1 ? tmp7975 : tmp8195;
  assign tmp8193 = s2 ? tmp8194 : tmp8179;
  assign tmp8186 = s3 ? tmp8187 : tmp8193;
  assign tmp8201 = l1 ? tmp7981 : tmp7955;
  assign tmp8200 = ~(s0 ? tmp8029 : tmp8201);
  assign tmp8199 = s1 ? tmp8024 : tmp8200;
  assign tmp8204 = ~(l1 ? tmp7981 : tmp7956);
  assign tmp8203 = s0 ? tmp7972 : tmp8204;
  assign tmp8202 = s1 ? tmp8020 : tmp8203;
  assign tmp8198 = s2 ? tmp8199 : tmp8202;
  assign tmp8208 = ~(l1 ? tmp7981 : tmp8016);
  assign tmp8207 = s0 ? tmp7977 : tmp8208;
  assign tmp8206 = s1 ? tmp8207 : tmp8184;
  assign tmp8205 = s2 ? tmp8206 : tmp8041;
  assign tmp8197 = s3 ? tmp8198 : tmp8205;
  assign tmp8185 = s4 ? tmp8186 : tmp8197;
  assign tmp8177 = s5 ? tmp8178 : tmp8185;
  assign tmp8211 = s6 ? tmp7997 : tmp8177;
  assign tmp8216 = s0 ? tmp8008 : tmp8182;
  assign tmp8218 = l1 ? tmp7955 : 1;
  assign tmp8217 = s0 ? tmp7972 : tmp8218;
  assign tmp8215 = s1 ? tmp8216 : tmp8217;
  assign tmp8214 = s2 ? tmp8008 : tmp8215;
  assign tmp8222 = s1 ? tmp8008 : tmp8009;
  assign tmp8223 = s1 ? tmp8008 : tmp8007;
  assign tmp8221 = s2 ? tmp8222 : tmp8223;
  assign tmp8225 = s1 ? 1 : tmp8196;
  assign tmp8224 = s2 ? tmp8225 : tmp8179;
  assign tmp8220 = s3 ? tmp8221 : tmp8224;
  assign tmp8229 = l1 ? tmp7978 : tmp7956;
  assign tmp8230 = l1 ? tmp8070 : tmp7955;
  assign tmp8228 = s1 ? tmp8229 : tmp8230;
  assign tmp8232 = ~(l1 ? tmp8070 : tmp7956);
  assign tmp8231 = ~(s1 ? tmp8008 : tmp8232);
  assign tmp8227 = s2 ? tmp8228 : tmp8231;
  assign tmp8234 = l1 ? tmp8070 : tmp8016;
  assign tmp8235 = ~(l1 ? tmp7955 : 1);
  assign tmp8233 = s1 ? tmp8234 : tmp8235;
  assign tmp8226 = ~(s3 ? tmp8227 : tmp8233);
  assign tmp8219 = s4 ? tmp8220 : tmp8226;
  assign tmp8213 = s5 ? tmp8214 : tmp8219;
  assign tmp8212 = s6 ? tmp8213 : tmp7997;
  assign tmp8210 = s7 ? tmp8211 : tmp8212;
  assign tmp8242 = s1 ? tmp8008 : tmp8192;
  assign tmp8241 = s2 ? tmp8188 : tmp8242;
  assign tmp8240 = s3 ? tmp8241 : tmp8193;
  assign tmp8245 = s1 ? tmp8020 : tmp8204;
  assign tmp8244 = s2 ? tmp8199 : tmp8245;
  assign tmp8247 = l1 ? tmp7981 : tmp8016;
  assign tmp8248 = ~(l1 ? tmp7956 : 1);
  assign tmp8246 = ~(s1 ? tmp8247 : tmp8248);
  assign tmp8243 = s3 ? tmp8244 : tmp8246;
  assign tmp8239 = s4 ? tmp8240 : tmp8243;
  assign tmp8238 = s5 ? tmp8178 : tmp8239;
  assign tmp8237 = s6 ? tmp7997 : tmp8238;
  assign tmp8252 = s3 ? tmp8221 : tmp8193;
  assign tmp8256 = ~(s0 ? tmp8029 : tmp8230);
  assign tmp8255 = s1 ? tmp8024 : tmp8256;
  assign tmp8257 = s1 ? tmp8008 : tmp8232;
  assign tmp8254 = s2 ? tmp8255 : tmp8257;
  assign tmp8258 = ~(s1 ? tmp8234 : tmp8235);
  assign tmp8253 = s3 ? tmp8254 : tmp8258;
  assign tmp8251 = s4 ? tmp8252 : tmp8253;
  assign tmp8250 = s5 ? tmp8214 : tmp8251;
  assign tmp8249 = s6 ? tmp8250 : tmp8213;
  assign tmp8236 = s7 ? tmp8237 : tmp8249;
  assign tmp8209 = s8 ? tmp8210 : tmp8236;
  assign tmp8176 = s9 ? tmp8177 : tmp8209;
  assign tmp8267 = s1 ? tmp8191 : tmp8007;
  assign tmp8266 = s2 ? tmp8222 : tmp8267;
  assign tmp8265 = s3 ? tmp8266 : tmp8193;
  assign tmp8271 = s0 ? tmp7972 : tmp8232;
  assign tmp8270 = s1 ? tmp8008 : tmp8271;
  assign tmp8269 = s2 ? tmp8255 : tmp8270;
  assign tmp8275 = ~(l1 ? tmp8070 : tmp8016);
  assign tmp8274 = s0 ? tmp7977 : tmp8275;
  assign tmp8273 = s1 ? tmp8274 : tmp8218;
  assign tmp8272 = s2 ? tmp8273 : tmp8041;
  assign tmp8268 = s3 ? tmp8269 : tmp8272;
  assign tmp8264 = s4 ? tmp8265 : tmp8268;
  assign tmp8263 = s5 ? tmp8214 : tmp8264;
  assign tmp8262 = s6 ? tmp8263 : tmp8213;
  assign tmp8261 = s7 ? tmp8211 : tmp8262;
  assign tmp8260 = s8 ? tmp8210 : tmp8261;
  assign tmp8259 = s9 ? tmp8177 : tmp8260;
  assign tmp8175 = s10 ? tmp8176 : tmp8259;
  assign tmp8280 = l1 ? 1 : tmp8002;
  assign tmp8282 = s0 ? tmp8280 : tmp8001;
  assign tmp8284 = l1 ? 1 : tmp7956;
  assign tmp8283 = s0 ? tmp8280 : tmp8284;
  assign tmp8281 = s1 ? tmp8282 : tmp8283;
  assign tmp8279 = s2 ? tmp8280 : tmp8281;
  assign tmp8290 = l1 ? tmp7955 : tmp8002;
  assign tmp8289 = s0 ? tmp8290 : tmp8280;
  assign tmp8288 = s1 ? tmp8289 : tmp8009;
  assign tmp8292 = s0 ? tmp8280 : tmp8009;
  assign tmp8293 = s0 ? tmp8280 : tmp7972;
  assign tmp8291 = s1 ? tmp8292 : tmp8293;
  assign tmp8287 = s2 ? tmp8288 : tmp8291;
  assign tmp8297 = ~(l1 ? tmp7955 : tmp7981);
  assign tmp8296 = s0 ? tmp7977 : tmp8297;
  assign tmp8295 = s1 ? tmp7975 : tmp8296;
  assign tmp8299 = s0 ? tmp7972 : tmp8182;
  assign tmp8298 = s1 ? tmp7972 : tmp8299;
  assign tmp8294 = s2 ? tmp8295 : tmp8298;
  assign tmp8286 = s3 ? tmp8287 : tmp8294;
  assign tmp8303 = l1 ? tmp7957 : 1;
  assign tmp8302 = s1 ? tmp7977 : tmp8303;
  assign tmp8306 = ~(l1 ? tmp7957 : 1);
  assign tmp8305 = s0 ? tmp7972 : tmp8306;
  assign tmp8304 = ~(s1 ? tmp8280 : tmp8305);
  assign tmp8301 = s2 ? tmp8302 : tmp8304;
  assign tmp8309 = ~(l1 ? tmp7957 : tmp7981);
  assign tmp8308 = s0 ? tmp7977 : tmp8309;
  assign tmp8310 = s0 ? tmp7972 : tmp8284;
  assign tmp8307 = ~(s1 ? tmp8308 : tmp8310);
  assign tmp8300 = ~(s3 ? tmp8301 : tmp8307);
  assign tmp8285 = s4 ? tmp8286 : tmp8300;
  assign tmp8278 = s5 ? tmp8279 : tmp8285;
  assign tmp8313 = s6 ? tmp7997 : tmp8278;
  assign tmp8317 = l1 ? 1 : tmp8026;
  assign tmp8319 = s0 ? tmp8317 : tmp8001;
  assign tmp8321 = l1 ? 1 : tmp7955;
  assign tmp8320 = s0 ? tmp8317 : tmp8321;
  assign tmp8318 = s1 ? tmp8319 : tmp8320;
  assign tmp8316 = s2 ? tmp8317 : tmp8318;
  assign tmp8327 = l1 ? tmp7955 : tmp8026;
  assign tmp8326 = s0 ? tmp8327 : tmp8317;
  assign tmp8325 = s1 ? tmp8326 : tmp8009;
  assign tmp8329 = s0 ? tmp8317 : tmp7972;
  assign tmp8328 = s1 ? tmp8317 : tmp8329;
  assign tmp8324 = s2 ? tmp8325 : tmp8328;
  assign tmp8331 = s1 ? 1 : tmp8297;
  assign tmp8332 = s1 ? tmp7972 : tmp8025;
  assign tmp8330 = s2 ? tmp8331 : tmp8332;
  assign tmp8323 = s3 ? tmp8324 : tmp8330;
  assign tmp8335 = s1 ? tmp7978 : tmp8303;
  assign tmp8337 = ~(l1 ? tmp7957 : tmp7978);
  assign tmp8336 = ~(s1 ? tmp8317 : tmp8337);
  assign tmp8334 = s2 ? tmp8335 : tmp8336;
  assign tmp8339 = l1 ? tmp7957 : tmp7981;
  assign tmp8340 = ~(l1 ? 1 : tmp7955);
  assign tmp8338 = s1 ? tmp8339 : tmp8340;
  assign tmp8333 = ~(s3 ? tmp8334 : tmp8338);
  assign tmp8322 = s4 ? tmp8323 : tmp8333;
  assign tmp8315 = s5 ? tmp8316 : tmp8322;
  assign tmp8314 = s6 ? tmp8315 : tmp7997;
  assign tmp8312 = s7 ? tmp8313 : tmp8314;
  assign tmp8347 = s1 ? tmp8280 : tmp8293;
  assign tmp8346 = s2 ? tmp8288 : tmp8347;
  assign tmp8345 = s3 ? tmp8346 : tmp8294;
  assign tmp8350 = ~(s1 ? tmp8280 : tmp8306);
  assign tmp8349 = s2 ? tmp8302 : tmp8350;
  assign tmp8352 = ~(l1 ? 1 : tmp7956);
  assign tmp8351 = s1 ? tmp8339 : tmp8352;
  assign tmp8348 = ~(s3 ? tmp8349 : tmp8351);
  assign tmp8344 = s4 ? tmp8345 : tmp8348;
  assign tmp8343 = s5 ? tmp8279 : tmp8344;
  assign tmp8342 = s6 ? tmp7997 : tmp8343;
  assign tmp8359 = s0 ? tmp7972 : tmp8025;
  assign tmp8358 = s1 ? tmp7972 : tmp8359;
  assign tmp8357 = s2 ? tmp8295 : tmp8358;
  assign tmp8356 = s3 ? tmp8324 : tmp8357;
  assign tmp8355 = s4 ? tmp8356 : tmp8333;
  assign tmp8354 = s5 ? tmp8316 : tmp8355;
  assign tmp8353 = s6 ? tmp8354 : tmp8315;
  assign tmp8341 = s7 ? tmp8342 : tmp8353;
  assign tmp8311 = s8 ? tmp8312 : tmp8341;
  assign tmp8277 = s9 ? tmp8278 : tmp8311;
  assign tmp8369 = s0 ? tmp8317 : tmp8009;
  assign tmp8368 = s1 ? tmp8369 : tmp8329;
  assign tmp8367 = s2 ? tmp8325 : tmp8368;
  assign tmp8366 = s3 ? tmp8367 : tmp8357;
  assign tmp8373 = s0 ? tmp7972 : tmp8337;
  assign tmp8372 = ~(s1 ? tmp8317 : tmp8373);
  assign tmp8371 = s2 ? tmp8335 : tmp8372;
  assign tmp8375 = s0 ? tmp7972 : tmp8321;
  assign tmp8374 = ~(s1 ? tmp8308 : tmp8375);
  assign tmp8370 = ~(s3 ? tmp8371 : tmp8374);
  assign tmp8365 = s4 ? tmp8366 : tmp8370;
  assign tmp8364 = s5 ? tmp8316 : tmp8365;
  assign tmp8363 = s6 ? tmp8364 : tmp8315;
  assign tmp8362 = s7 ? tmp8313 : tmp8363;
  assign tmp8361 = s8 ? tmp8312 : tmp8362;
  assign tmp8360 = s9 ? tmp8278 : tmp8361;
  assign tmp8276 = s10 ? tmp8277 : tmp8360;
  assign tmp8174 = s11 ? tmp8175 : tmp8276;
  assign tmp7947 = s12 ? tmp7948 : tmp8174;
  assign tmp8382 = s1 ? tmp8001 : tmp8280;
  assign tmp8384 = s0 ? tmp8182 : tmp8280;
  assign tmp8383 = s1 ? tmp8293 : tmp8384;
  assign tmp8381 = s2 ? tmp8382 : tmp8383;
  assign tmp8389 = s0 ? tmp8229 : tmp8280;
  assign tmp8388 = s1 ? tmp8389 : tmp7972;
  assign tmp8391 = s0 ? tmp8280 : tmp7983;
  assign tmp8390 = s1 ? tmp8001 : tmp8391;
  assign tmp8387 = s2 ? tmp8388 : tmp8390;
  assign tmp8393 = s1 ? tmp8123 : tmp8340;
  assign tmp8395 = l1 ? tmp8016 : tmp7981;
  assign tmp8394 = s1 ? tmp8395 : tmp8352;
  assign tmp8392 = ~(s2 ? tmp8393 : tmp8394);
  assign tmp8386 = s3 ? tmp8387 : tmp8392;
  assign tmp8399 = s0 ? tmp8029 : tmp8321;
  assign tmp8398 = s1 ? tmp8229 : tmp8399;
  assign tmp8400 = s1 ? tmp8280 : tmp8284;
  assign tmp8397 = s2 ? tmp8398 : tmp8400;
  assign tmp8402 = s1 ? tmp8317 : tmp8280;
  assign tmp8401 = s2 ? tmp8402 : tmp8029;
  assign tmp8396 = s3 ? tmp8397 : tmp8401;
  assign tmp8385 = s4 ? tmp8386 : tmp8396;
  assign tmp8380 = s5 ? tmp8381 : tmp8385;
  assign tmp8406 = ~(s5 ? tmp8381 : tmp8385);
  assign tmp8405 = s6 ? tmp7997 : tmp8406;
  assign tmp8411 = s0 ? tmp8395 : tmp7957;
  assign tmp8412 = s0 ? tmp7981 : tmp8395;
  assign tmp8410 = s1 ? tmp8411 : tmp8412;
  assign tmp8409 = s2 ? tmp8395 : tmp8410;
  assign tmp8418 = l1 ? tmp8016 : tmp7982;
  assign tmp8417 = s0 ? tmp8418 : tmp8395;
  assign tmp8416 = s1 ? tmp8417 : tmp7957;
  assign tmp8420 = s0 ? tmp8395 : tmp7987;
  assign tmp8419 = s1 ? tmp8395 : tmp8420;
  assign tmp8415 = s2 ? tmp8416 : tmp8419;
  assign tmp8422 = s1 ? tmp7987 : tmp8340;
  assign tmp8424 = l1 ? tmp7957 : tmp7982;
  assign tmp8423 = s1 ? tmp8395 : tmp8424;
  assign tmp8421 = s2 ? tmp8422 : tmp8423;
  assign tmp8414 = s3 ? tmp8415 : tmp8421;
  assign tmp8428 = l1 ? tmp7978 : tmp7955;
  assign tmp8427 = s1 ? tmp8229 : tmp8428;
  assign tmp8429 = ~(s1 ? tmp8395 : tmp8027);
  assign tmp8426 = s2 ? tmp8427 : tmp8429;
  assign tmp8431 = l1 ? tmp7978 : tmp8026;
  assign tmp8432 = ~(l1 ? tmp8016 : tmp7981);
  assign tmp8430 = s1 ? tmp8431 : tmp8432;
  assign tmp8425 = ~(s3 ? tmp8426 : tmp8430);
  assign tmp8413 = s4 ? tmp8414 : tmp8425;
  assign tmp8408 = s5 ? tmp8409 : tmp8413;
  assign tmp8407 = s6 ? tmp8408 : tmp7997;
  assign tmp8404 = s7 ? tmp8405 : tmp8407;
  assign tmp8437 = s3 ? tmp8397 : tmp8402;
  assign tmp8436 = s4 ? tmp8386 : tmp8437;
  assign tmp8435 = ~(s5 ? tmp8381 : tmp8436);
  assign tmp8434 = s6 ? tmp7997 : tmp8435;
  assign tmp8439 = s5 ? tmp8381 : tmp8436;
  assign tmp8440 = ~(s5 ? tmp8409 : tmp8413);
  assign tmp8438 = ~(s6 ? tmp8439 : tmp8440);
  assign tmp8433 = s7 ? tmp8434 : tmp8438;
  assign tmp8403 = ~(s8 ? tmp8404 : tmp8433);
  assign tmp8379 = s9 ? tmp8380 : tmp8403;
  assign tmp8444 = ~(s6 ? tmp8380 : tmp8440);
  assign tmp8443 = s7 ? tmp8405 : tmp8444;
  assign tmp8442 = ~(s8 ? tmp8404 : tmp8443);
  assign tmp8441 = s9 ? tmp8380 : tmp8442;
  assign tmp8378 = s10 ? tmp8379 : tmp8441;
  assign tmp8445 = ~(s10 ? tmp7950 : tmp8089);
  assign tmp8377 = s11 ? tmp8378 : tmp8445;
  assign tmp8452 = s0 ? tmp7958 : tmp7980;
  assign tmp8453 = s0 ? tmp7958 : tmp7983;
  assign tmp8451 = s1 ? tmp8452 : tmp8453;
  assign tmp8450 = s2 ? tmp7958 : tmp8451;
  assign tmp8459 = l1 ? tmp7978 : tmp7957;
  assign tmp8458 = s0 ? tmp8459 : tmp7958;
  assign tmp8457 = s1 ? tmp8458 : tmp8117;
  assign tmp8461 = s0 ? tmp7958 : tmp8117;
  assign tmp8460 = s1 ? tmp8461 : tmp7958;
  assign tmp8456 = s2 ? tmp8457 : tmp8460;
  assign tmp8463 = s1 ? tmp8123 : tmp8015;
  assign tmp8465 = s0 ? tmp7980 : tmp7993;
  assign tmp8464 = ~(s1 ? tmp8465 : tmp7961);
  assign tmp8462 = ~(s2 ? tmp8463 : tmp8464);
  assign tmp8455 = s3 ? tmp8456 : tmp8462;
  assign tmp8470 = l1 ? tmp7956 : tmp7955;
  assign tmp8469 = s0 ? tmp8029 : tmp8470;
  assign tmp8468 = s1 ? tmp8229 : tmp8469;
  assign tmp8471 = s1 ? tmp7958 : tmp7956;
  assign tmp8467 = s2 ? tmp8468 : tmp8471;
  assign tmp8474 = l1 ? tmp7956 : tmp8016;
  assign tmp8473 = s1 ? tmp8474 : tmp7983;
  assign tmp8475 = s1 ? tmp8029 : tmp7980;
  assign tmp8472 = s2 ? tmp8473 : tmp8475;
  assign tmp8466 = s3 ? tmp8467 : tmp8472;
  assign tmp8454 = s4 ? tmp8455 : tmp8466;
  assign tmp8449 = s5 ? tmp8450 : tmp8454;
  assign tmp8479 = ~(s5 ? tmp8450 : tmp8454);
  assign tmp8478 = s6 ? tmp7997 : tmp8479;
  assign tmp8485 = l1 ? tmp8070 : tmp8002;
  assign tmp8484 = s0 ? tmp8082 : tmp8485;
  assign tmp8486 = s0 ? tmp8082 : tmp7987;
  assign tmp8483 = s1 ? tmp8484 : tmp8486;
  assign tmp8482 = s2 ? tmp8082 : tmp8483;
  assign tmp8491 = s0 ? tmp8126 : tmp8082;
  assign tmp8490 = s1 ? tmp8491 : tmp8009;
  assign tmp8489 = s2 ? tmp8490 : tmp8082;
  assign tmp8493 = s1 ? tmp7987 : tmp8015;
  assign tmp8495 = ~(l1 ? tmp7957 : tmp7969);
  assign tmp8494 = ~(s1 ? tmp8465 : tmp8495);
  assign tmp8492 = s2 ? tmp8493 : tmp8494;
  assign tmp8488 = s3 ? tmp8489 : tmp8492;
  assign tmp8498 = s1 ? tmp8229 : tmp8470;
  assign tmp8499 = ~(s1 ? tmp8082 : tmp7982);
  assign tmp8497 = s2 ? tmp8498 : tmp8499;
  assign tmp8501 = s1 ? tmp8474 : tmp7990;
  assign tmp8500 = s2 ? tmp8501 : tmp7980;
  assign tmp8496 = ~(s3 ? tmp8497 : tmp8500);
  assign tmp8487 = s4 ? tmp8488 : tmp8496;
  assign tmp8481 = s5 ? tmp8482 : tmp8487;
  assign tmp8480 = s6 ? tmp8481 : tmp7997;
  assign tmp8477 = s7 ? tmp8478 : tmp8480;
  assign tmp8507 = s2 ? tmp8457 : tmp7958;
  assign tmp8506 = s3 ? tmp8507 : tmp8462;
  assign tmp8508 = s3 ? tmp8467 : tmp8473;
  assign tmp8505 = s4 ? tmp8506 : tmp8508;
  assign tmp8504 = ~(s5 ? tmp8450 : tmp8505);
  assign tmp8503 = s6 ? tmp7997 : tmp8504;
  assign tmp8513 = s2 ? tmp8468 : tmp8499;
  assign tmp8512 = ~(s3 ? tmp8513 : tmp8501);
  assign tmp8511 = s4 ? tmp8488 : tmp8512;
  assign tmp8510 = s5 ? tmp8482 : tmp8511;
  assign tmp8516 = ~(s3 ? tmp8497 : tmp8501);
  assign tmp8515 = s4 ? tmp8488 : tmp8516;
  assign tmp8514 = s5 ? tmp8482 : tmp8515;
  assign tmp8509 = s6 ? tmp8510 : tmp8514;
  assign tmp8502 = s7 ? tmp8503 : tmp8509;
  assign tmp8476 = ~(s8 ? tmp8477 : tmp8502);
  assign tmp8448 = s9 ? tmp8449 : tmp8476;
  assign tmp8526 = s0 ? tmp8082 : tmp8009;
  assign tmp8525 = s1 ? tmp8526 : tmp8082;
  assign tmp8524 = s2 ? tmp8490 : tmp8525;
  assign tmp8523 = s3 ? tmp8524 : tmp8492;
  assign tmp8528 = s2 ? tmp8501 : tmp8475;
  assign tmp8527 = ~(s3 ? tmp8513 : tmp8528);
  assign tmp8522 = s4 ? tmp8523 : tmp8527;
  assign tmp8521 = s5 ? tmp8482 : tmp8522;
  assign tmp8520 = s6 ? tmp8521 : tmp8481;
  assign tmp8519 = s7 ? tmp8478 : tmp8520;
  assign tmp8518 = ~(s8 ? tmp8477 : tmp8519);
  assign tmp8517 = s9 ? tmp8449 : tmp8518;
  assign tmp8447 = s10 ? tmp8448 : tmp8517;
  assign tmp8534 = s0 ? tmp8108 : tmp8459;
  assign tmp8533 = s1 ? tmp8534 : tmp8108;
  assign tmp8532 = s2 ? tmp8108 : tmp8533;
  assign tmp8539 = s0 ? tmp8064 : tmp8108;
  assign tmp8538 = s1 ? tmp8539 : tmp7968;
  assign tmp8541 = s0 ? tmp8108 : tmp7972;
  assign tmp8540 = s1 ? tmp8108 : tmp8541;
  assign tmp8537 = s2 ? tmp8538 : tmp8540;
  assign tmp8545 = ~(l2 ? 1 : tmp7956);
  assign tmp8544 = s0 ? tmp7977 : tmp8545;
  assign tmp8543 = s1 ? tmp7975 : tmp8544;
  assign tmp8547 = l1 ? tmp7956 : tmp7982;
  assign tmp8546 = s1 ? tmp8108 : tmp8547;
  assign tmp8542 = s2 ? tmp8543 : tmp8546;
  assign tmp8536 = s3 ? tmp8537 : tmp8542;
  assign tmp8551 = s0 ? tmp8029 : tmp8030;
  assign tmp8550 = s1 ? tmp8229 : tmp8551;
  assign tmp8553 = s0 ? tmp8033 : tmp8124;
  assign tmp8552 = s1 ? tmp8553 : tmp8034;
  assign tmp8549 = s2 ? tmp8550 : tmp8552;
  assign tmp8557 = ~(l1 ? tmp7957 : tmp8026);
  assign tmp8556 = s0 ? tmp7977 : tmp8557;
  assign tmp8555 = s1 ? tmp8556 : tmp8108;
  assign tmp8558 = ~(s1 ? tmp8029 : tmp8033);
  assign tmp8554 = ~(s2 ? tmp8555 : tmp8558);
  assign tmp8548 = ~(s3 ? tmp8549 : tmp8554);
  assign tmp8535 = s4 ? tmp8536 : tmp8548;
  assign tmp8531 = s5 ? tmp8532 : tmp8535;
  assign tmp8561 = s6 ? tmp7997 : tmp8531;
  assign tmp8567 = l1 ? tmp7978 : 0;
  assign tmp8566 = s0 ? tmp8112 : tmp8567;
  assign tmp8568 = s0 ? tmp8112 : tmp8108;
  assign tmp8565 = s1 ? tmp8566 : tmp8568;
  assign tmp8564 = s2 ? tmp8112 : tmp8565;
  assign tmp8573 = s0 ? tmp8064 : tmp8112;
  assign tmp8572 = s1 ? tmp8573 : tmp8058;
  assign tmp8575 = s0 ? tmp8112 : tmp7972;
  assign tmp8574 = s1 ? tmp8112 : tmp8575;
  assign tmp8571 = s2 ? tmp8572 : tmp8574;
  assign tmp8577 = s1 ? 1 : tmp8545;
  assign tmp8578 = s1 ? tmp8112 : tmp8547;
  assign tmp8576 = s2 ? tmp8577 : tmp8578;
  assign tmp8570 = s3 ? tmp8571 : tmp8576;
  assign tmp8581 = s1 ? tmp8229 : tmp8030;
  assign tmp8582 = ~(s1 ? tmp8112 : tmp8035);
  assign tmp8580 = s2 ? tmp8581 : tmp8582;
  assign tmp8583 = s1 ? tmp8030 : tmp8124;
  assign tmp8579 = ~(s3 ? tmp8580 : tmp8583);
  assign tmp8569 = s4 ? tmp8570 : tmp8579;
  assign tmp8563 = s5 ? tmp8564 : tmp8569;
  assign tmp8562 = s6 ? tmp8563 : tmp7997;
  assign tmp8560 = s7 ? tmp8561 : tmp8562;
  assign tmp8591 = l1 ? tmp7957 : tmp7956;
  assign tmp8590 = s1 ? tmp8553 : tmp8591;
  assign tmp8589 = s2 ? tmp8550 : tmp8590;
  assign tmp8592 = s1 ? tmp8140 : tmp8124;
  assign tmp8588 = ~(s3 ? tmp8589 : tmp8592);
  assign tmp8587 = s4 ? tmp8536 : tmp8588;
  assign tmp8586 = s5 ? tmp8532 : tmp8587;
  assign tmp8585 = s6 ? tmp7997 : tmp8586;
  assign tmp8597 = s2 ? tmp8543 : tmp8578;
  assign tmp8596 = s3 ? tmp8571 : tmp8597;
  assign tmp8602 = ~(l1 ? 1 : tmp7982);
  assign tmp8601 = s0 ? tmp8033 : tmp8602;
  assign tmp8600 = s1 ? tmp8601 : tmp8591;
  assign tmp8599 = s2 ? tmp8550 : tmp8600;
  assign tmp8598 = ~(s3 ? tmp8599 : tmp8583);
  assign tmp8595 = s4 ? tmp8596 : tmp8598;
  assign tmp8594 = s5 ? tmp8564 : tmp8595;
  assign tmp8593 = s6 ? tmp8594 : tmp8563;
  assign tmp8584 = s7 ? tmp8585 : tmp8593;
  assign tmp8559 = s8 ? tmp8560 : tmp8584;
  assign tmp8530 = s9 ? tmp8531 : tmp8559;
  assign tmp8611 = s1 ? tmp8601 : tmp8034;
  assign tmp8610 = s2 ? tmp8550 : tmp8611;
  assign tmp8614 = s0 ? tmp7977 : tmp8159;
  assign tmp8613 = s1 ? tmp8614 : tmp8108;
  assign tmp8612 = ~(s2 ? tmp8613 : tmp8558);
  assign tmp8609 = ~(s3 ? tmp8610 : tmp8612);
  assign tmp8608 = s4 ? tmp8596 : tmp8609;
  assign tmp8607 = s5 ? tmp8564 : tmp8608;
  assign tmp8606 = s6 ? tmp8607 : tmp8563;
  assign tmp8605 = s7 ? tmp8561 : tmp8606;
  assign tmp8604 = s8 ? tmp8560 : tmp8605;
  assign tmp8603 = s9 ? tmp8531 : tmp8604;
  assign tmp8529 = ~(s10 ? tmp8530 : tmp8603);
  assign tmp8446 = s11 ? tmp8447 : tmp8529;
  assign tmp8376 = ~(s12 ? tmp8377 : tmp8446);
  assign tmp7946 = s13 ? tmp7947 : tmp8376;
  assign tmp8624 = l1 ? tmp7978 : tmp7969;
  assign tmp8623 = s1 ? tmp8624 : tmp7972;
  assign tmp8625 = s1 ? tmp7972 : tmp8192;
  assign tmp8622 = s2 ? tmp8623 : tmp8625;
  assign tmp8630 = s0 ? 1 : tmp7972;
  assign tmp8629 = s1 ? tmp8630 : tmp7972;
  assign tmp8632 = s0 ? tmp7972 : tmp7983;
  assign tmp8631 = s1 ? tmp8624 : tmp8632;
  assign tmp8628 = s2 ? tmp8629 : tmp8631;
  assign tmp8634 = s1 ? tmp8123 : 0;
  assign tmp8635 = s1 ? tmp8395 : 0;
  assign tmp8633 = ~(s2 ? tmp8634 : tmp8635);
  assign tmp8627 = s3 ? tmp8628 : tmp8633;
  assign tmp8638 = s1 ? tmp7972 : 1;
  assign tmp8637 = s2 ? 1 : tmp8638;
  assign tmp8636 = s3 ? tmp8637 : tmp7972;
  assign tmp8626 = s4 ? tmp8627 : tmp8636;
  assign tmp8621 = s5 ? tmp8622 : tmp8626;
  assign tmp8644 = l1 ? tmp8016 : tmp8048;
  assign tmp8646 = s0 ? tmp8644 : tmp8058;
  assign tmp8648 = l1 ? tmp7981 : tmp8048;
  assign tmp8647 = s0 ? tmp8648 : tmp8016;
  assign tmp8645 = s1 ? tmp8646 : tmp8647;
  assign tmp8643 = s2 ? tmp8644 : tmp8645;
  assign tmp8652 = s1 ? tmp8644 : tmp8058;
  assign tmp8654 = s0 ? tmp8644 : tmp8082;
  assign tmp8653 = s1 ? tmp8644 : tmp8654;
  assign tmp8651 = s2 ? tmp8652 : tmp8653;
  assign tmp8656 = s1 ? tmp7987 : 0;
  assign tmp8658 = l1 ? tmp7957 : tmp8048;
  assign tmp8657 = s1 ? tmp8418 : tmp8658;
  assign tmp8655 = s2 ? tmp8656 : tmp8657;
  assign tmp8650 = s3 ? tmp8651 : tmp8655;
  assign tmp8661 = s1 ? tmp7978 : tmp7977;
  assign tmp8662 = ~(s1 ? tmp8644 : tmp8048);
  assign tmp8660 = s2 ? tmp8661 : tmp8662;
  assign tmp8664 = ~(l2 ? 1 : 0);
  assign tmp8663 = s1 ? tmp7977 : tmp8664;
  assign tmp8659 = ~(s3 ? tmp8660 : tmp8663);
  assign tmp8649 = s4 ? tmp8650 : tmp8659;
  assign tmp8642 = s5 ? tmp8643 : tmp8649;
  assign tmp8641 = s6 ? tmp8642 : tmp7997;
  assign tmp8640 = s7 ? tmp7996 : tmp8641;
  assign tmp8672 = s0 ? tmp7972 : tmp8117;
  assign tmp8671 = s1 ? tmp8630 : tmp8672;
  assign tmp8674 = s0 ? tmp8624 : tmp8117;
  assign tmp8673 = s1 ? tmp8674 : tmp8632;
  assign tmp8670 = s2 ? tmp8671 : tmp8673;
  assign tmp8677 = s0 ? tmp7972 : tmp8123;
  assign tmp8676 = s1 ? tmp8677 : tmp7976;
  assign tmp8679 = s0 ? tmp7980 : tmp8432;
  assign tmp8680 = ~(s0 ? tmp7972 : 0);
  assign tmp8678 = ~(s1 ? tmp8679 : tmp8680);
  assign tmp8675 = ~(s2 ? tmp8676 : tmp8678);
  assign tmp8669 = s3 ? tmp8670 : tmp8675;
  assign tmp8684 = s0 ? tmp8025 : 0;
  assign tmp8685 = ~(s0 ? tmp8029 : 1);
  assign tmp8683 = s1 ? tmp8684 : tmp8685;
  assign tmp8687 = s0 ? tmp8033 : tmp7972;
  assign tmp8686 = ~(s1 ? tmp8687 : tmp8680);
  assign tmp8682 = s2 ? tmp8683 : tmp8686;
  assign tmp8690 = s0 ? tmp7977 : tmp7968;
  assign tmp8691 = s0 ? tmp7972 : tmp7968;
  assign tmp8689 = s1 ? tmp8690 : tmp8691;
  assign tmp8688 = s2 ? tmp8689 : tmp8040;
  assign tmp8681 = ~(s3 ? tmp8682 : tmp8688);
  assign tmp8668 = s4 ? tmp8669 : tmp8681;
  assign tmp8667 = s5 ? tmp8622 : tmp8668;
  assign tmp8666 = s6 ? tmp8667 : tmp8621;
  assign tmp8692 = ~(s6 ? tmp8076 : tmp8642);
  assign tmp8665 = ~(s7 ? tmp8666 : tmp8692);
  assign tmp8639 = ~(s8 ? tmp8640 : tmp8665);
  assign tmp8620 = s9 ? tmp8621 : tmp8639;
  assign tmp8696 = ~(s6 ? tmp7951 : tmp8642);
  assign tmp8695 = ~(s7 ? tmp8666 : tmp8696);
  assign tmp8694 = ~(s8 ? tmp8640 : tmp8695);
  assign tmp8693 = s9 ? tmp8621 : tmp8694;
  assign tmp8619 = s10 ? tmp8620 : tmp8693;
  assign tmp8704 = s1 ? tmp8644 : tmp8658;
  assign tmp8706 = s0 ? tmp8658 : tmp8058;
  assign tmp8708 = l1 ? tmp7957 : tmp8016;
  assign tmp8707 = s0 ? tmp8648 : tmp8708;
  assign tmp8705 = s1 ? tmp8706 : tmp8707;
  assign tmp8703 = s2 ? tmp8704 : tmp8705;
  assign tmp8712 = s1 ? tmp8658 : tmp8058;
  assign tmp8714 = s0 ? tmp8658 : tmp8082;
  assign tmp8713 = s1 ? tmp8644 : tmp8714;
  assign tmp8711 = s2 ? tmp8712 : tmp8713;
  assign tmp8716 = s1 ? tmp8069 : 0;
  assign tmp8715 = s2 ? tmp8716 : tmp8657;
  assign tmp8710 = s3 ? tmp8711 : tmp8715;
  assign tmp8719 = ~(s1 ? tmp8658 : tmp8042);
  assign tmp8718 = s2 ? tmp8156 : tmp8719;
  assign tmp8720 = s1 ? 1 : tmp8039;
  assign tmp8717 = ~(s3 ? tmp8718 : tmp8720);
  assign tmp8709 = s4 ? tmp8710 : tmp8717;
  assign tmp8702 = s5 ? tmp8703 : tmp8709;
  assign tmp8701 = s6 ? tmp8702 : tmp7997;
  assign tmp8700 = s7 ? tmp8133 : tmp8701;
  assign tmp8723 = ~(s5 ? tmp8703 : tmp8709);
  assign tmp8722 = s6 ? tmp8168 : tmp8723;
  assign tmp8721 = ~(s7 ? tmp8666 : tmp8722);
  assign tmp8699 = ~(s8 ? tmp8700 : tmp8721);
  assign tmp8698 = s9 ? tmp8621 : tmp8699;
  assign tmp8727 = s6 ? tmp8104 : tmp8723;
  assign tmp8726 = ~(s7 ? tmp8666 : tmp8727);
  assign tmp8725 = ~(s8 ? tmp8700 : tmp8726);
  assign tmp8724 = s9 ? tmp8621 : tmp8725;
  assign tmp8697 = s10 ? tmp8698 : tmp8724;
  assign tmp8618 = s11 ? tmp8619 : tmp8697;
  assign tmp8732 = s7 ? tmp8211 : tmp8641;
  assign tmp8734 = ~(s6 ? tmp8238 : tmp8642);
  assign tmp8733 = ~(s7 ? tmp8666 : tmp8734);
  assign tmp8731 = ~(s8 ? tmp8732 : tmp8733);
  assign tmp8730 = s9 ? tmp8621 : tmp8731;
  assign tmp8738 = ~(s6 ? tmp8177 : tmp8642);
  assign tmp8737 = ~(s7 ? tmp8666 : tmp8738);
  assign tmp8736 = ~(s8 ? tmp8732 : tmp8737);
  assign tmp8735 = s9 ? tmp8621 : tmp8736;
  assign tmp8729 = s10 ? tmp8730 : tmp8735;
  assign tmp8744 = s0 ? tmp8020 : tmp8008;
  assign tmp8743 = s1 ? tmp8744 : tmp8020;
  assign tmp8742 = s2 ? tmp8020 : tmp8743;
  assign tmp8749 = s0 ? tmp7977 : tmp8020;
  assign tmp8748 = s1 ? tmp8749 : tmp7972;
  assign tmp8751 = s0 ? tmp8020 : tmp7983;
  assign tmp8750 = s1 ? tmp8020 : tmp8751;
  assign tmp8747 = s2 ? tmp8748 : tmp8750;
  assign tmp8753 = s1 ? tmp8123 : tmp8235;
  assign tmp8754 = s1 ? tmp7981 : 0;
  assign tmp8752 = ~(s2 ? tmp8753 : tmp8754);
  assign tmp8746 = s3 ? tmp8747 : tmp8752;
  assign tmp8757 = s1 ? 1 : tmp8184;
  assign tmp8758 = s1 ? tmp8020 : tmp8184;
  assign tmp8756 = s2 ? tmp8757 : tmp8758;
  assign tmp8755 = s3 ? tmp8756 : tmp8020;
  assign tmp8745 = s4 ? tmp8746 : tmp8755;
  assign tmp8741 = s5 ? tmp8742 : tmp8745;
  assign tmp8766 = l1 ? tmp8070 : 0;
  assign tmp8765 = s0 ? tmp8648 : tmp8766;
  assign tmp8767 = s0 ? tmp8648 : tmp8247;
  assign tmp8764 = s1 ? tmp8765 : tmp8767;
  assign tmp8763 = s2 ? tmp8648 : tmp8764;
  assign tmp8772 = s0 ? tmp8644 : tmp8648;
  assign tmp8771 = s1 ? tmp8772 : tmp8058;
  assign tmp8774 = s0 ? tmp8648 : tmp8082;
  assign tmp8773 = s1 ? tmp8648 : tmp8774;
  assign tmp8770 = s2 ? tmp8771 : tmp8773;
  assign tmp8776 = s1 ? tmp7987 : tmp8235;
  assign tmp8778 = l1 ? tmp7981 : tmp7982;
  assign tmp8777 = s1 ? tmp8778 : tmp8658;
  assign tmp8775 = s2 ? tmp8776 : tmp8777;
  assign tmp8769 = s3 ? tmp8770 : tmp8775;
  assign tmp8781 = s1 ? tmp7978 : tmp8184;
  assign tmp8783 = ~(l1 ? tmp7956 : tmp7978);
  assign tmp8782 = ~(s1 ? tmp8648 : tmp8783);
  assign tmp8780 = s2 ? tmp8781 : tmp8782;
  assign tmp8784 = s1 ? tmp8184 : tmp8208;
  assign tmp8779 = ~(s3 ? tmp8780 : tmp8784);
  assign tmp8768 = s4 ? tmp8769 : tmp8779;
  assign tmp8762 = s5 ? tmp8763 : tmp8768;
  assign tmp8761 = s6 ? tmp8762 : tmp7997;
  assign tmp8760 = s7 ? tmp8313 : tmp8761;
  assign tmp8787 = ~(s5 ? tmp8742 : tmp8745);
  assign tmp8786 = s6 ? tmp7997 : tmp8787;
  assign tmp8788 = s6 ? tmp8343 : tmp8762;
  assign tmp8785 = s7 ? tmp8786 : tmp8788;
  assign tmp8759 = ~(s8 ? tmp8760 : tmp8785);
  assign tmp8740 = s9 ? tmp8741 : tmp8759;
  assign tmp8792 = s6 ? tmp8278 : tmp8762;
  assign tmp8791 = s7 ? tmp8786 : tmp8792;
  assign tmp8790 = ~(s8 ? tmp8760 : tmp8791);
  assign tmp8789 = s9 ? tmp8741 : tmp8790;
  assign tmp8739 = s10 ? tmp8740 : tmp8789;
  assign tmp8728 = s11 ? tmp8729 : tmp8739;
  assign tmp8617 = s12 ? tmp8618 : tmp8728;
  assign tmp8803 = s0 ? tmp8016 : tmp7957;
  assign tmp8804 = s0 ? tmp8247 : tmp8016;
  assign tmp8802 = s1 ? tmp8803 : tmp8804;
  assign tmp8801 = s2 ? tmp8016 : tmp8802;
  assign tmp8809 = s0 ? tmp8644 : tmp8016;
  assign tmp8808 = s1 ? tmp8809 : tmp7957;
  assign tmp8811 = s0 ? tmp8016 : tmp7987;
  assign tmp8810 = s1 ? tmp8016 : tmp8811;
  assign tmp8807 = s2 ? tmp8808 : tmp8810;
  assign tmp8813 = s1 ? tmp8395 : tmp8658;
  assign tmp8812 = s2 ? tmp8656 : tmp8813;
  assign tmp8806 = s3 ? tmp8807 : tmp8812;
  assign tmp8816 = ~(s1 ? tmp8016 : tmp8048);
  assign tmp8815 = s2 ? tmp8661 : tmp8816;
  assign tmp8817 = s1 ? tmp8624 : tmp8664;
  assign tmp8814 = ~(s3 ? tmp8815 : tmp8817);
  assign tmp8805 = s4 ? tmp8806 : tmp8814;
  assign tmp8800 = s5 ? tmp8801 : tmp8805;
  assign tmp8799 = s6 ? tmp8800 : tmp7997;
  assign tmp8798 = s7 ? tmp8405 : tmp8799;
  assign tmp8820 = ~(s5 ? tmp8801 : tmp8805);
  assign tmp8819 = s6 ? tmp8439 : tmp8820;
  assign tmp8818 = ~(s7 ? tmp8666 : tmp8819);
  assign tmp8797 = ~(s8 ? tmp8798 : tmp8818);
  assign tmp8796 = s9 ? tmp8621 : tmp8797;
  assign tmp8824 = s6 ? tmp8380 : tmp8820;
  assign tmp8823 = ~(s7 ? tmp8666 : tmp8824);
  assign tmp8822 = ~(s8 ? tmp8798 : tmp8823);
  assign tmp8821 = s9 ? tmp8621 : tmp8822;
  assign tmp8795 = s10 ? tmp8796 : tmp8821;
  assign tmp8794 = s11 ? tmp8795 : tmp8619;
  assign tmp8829 = s7 ? tmp8478 : tmp8761;
  assign tmp8832 = s5 ? tmp8450 : tmp8505;
  assign tmp8833 = ~(s5 ? tmp8763 : tmp8768);
  assign tmp8831 = ~(s6 ? tmp8832 : tmp8833);
  assign tmp8830 = s7 ? tmp8786 : tmp8831;
  assign tmp8828 = ~(s8 ? tmp8829 : tmp8830);
  assign tmp8827 = s9 ? tmp8741 : tmp8828;
  assign tmp8837 = ~(s6 ? tmp8449 : tmp8833);
  assign tmp8836 = s7 ? tmp8786 : tmp8837;
  assign tmp8835 = ~(s8 ? tmp8829 : tmp8836);
  assign tmp8834 = s9 ? tmp8741 : tmp8835;
  assign tmp8826 = s10 ? tmp8827 : tmp8834;
  assign tmp8841 = s7 ? tmp8561 : tmp8761;
  assign tmp8843 = s6 ? tmp8586 : tmp8762;
  assign tmp8842 = s7 ? tmp8786 : tmp8843;
  assign tmp8840 = ~(s8 ? tmp8841 : tmp8842);
  assign tmp8839 = s9 ? tmp8741 : tmp8840;
  assign tmp8847 = s6 ? tmp8531 : tmp8762;
  assign tmp8846 = s7 ? tmp8786 : tmp8847;
  assign tmp8845 = ~(s8 ? tmp8841 : tmp8846);
  assign tmp8844 = s9 ? tmp8741 : tmp8845;
  assign tmp8838 = s10 ? tmp8839 : tmp8844;
  assign tmp8825 = s11 ? tmp8826 : tmp8838;
  assign tmp8793 = s12 ? tmp8794 : tmp8825;
  assign tmp8616 = s13 ? tmp8617 : tmp8793;
  assign tmp8860 = s1 ? tmp7975 : 0;
  assign tmp8859 = s2 ? tmp8860 : tmp8063;
  assign tmp8858 = s3 ? tmp8056 : tmp8859;
  assign tmp8861 = ~(s3 ? tmp8096 : tmp8073);
  assign tmp8857 = s4 ? tmp8858 : tmp8861;
  assign tmp8856 = s5 ? tmp8046 : tmp8857;
  assign tmp8855 = s6 ? tmp8856 : tmp7997;
  assign tmp8854 = s7 ? tmp7996 : tmp8855;
  assign tmp8865 = s4 ? tmp8858 : tmp8066;
  assign tmp8864 = s5 ? tmp8046 : tmp8865;
  assign tmp8863 = s6 ? tmp8085 : tmp8864;
  assign tmp8862 = s7 ? tmp8075 : tmp8863;
  assign tmp8853 = s8 ? tmp8854 : tmp8862;
  assign tmp8852 = s9 ? tmp7951 : tmp8853;
  assign tmp8869 = s6 ? tmp8093 : tmp8856;
  assign tmp8868 = s7 ? tmp7996 : tmp8869;
  assign tmp8867 = s8 ? tmp8854 : tmp8868;
  assign tmp8866 = s9 ? tmp7951 : tmp8867;
  assign tmp8851 = s10 ? tmp8852 : tmp8866;
  assign tmp8880 = s0 ? tmp8139 : tmp8009;
  assign tmp8879 = s1 ? tmp8880 : tmp8150;
  assign tmp8878 = s2 ? tmp8148 : tmp8879;
  assign tmp8877 = s3 ? tmp8878 : tmp8151;
  assign tmp8876 = s4 ? tmp8877 : tmp8154;
  assign tmp8875 = s5 ? tmp8137 : tmp8876;
  assign tmp8874 = s6 ? tmp8875 : tmp7997;
  assign tmp8873 = s7 ? tmp8133 : tmp8874;
  assign tmp8872 = ~(s8 ? tmp8873 : tmp8160);
  assign tmp8871 = s9 ? tmp8104 : tmp8872;
  assign tmp8885 = ~(s5 ? tmp8137 : tmp8876);
  assign tmp8884 = ~(s6 ? tmp8104 : tmp8885);
  assign tmp8883 = s7 ? tmp8133 : tmp8884;
  assign tmp8882 = ~(s8 ? tmp8873 : tmp8883);
  assign tmp8881 = s9 ? tmp8104 : tmp8882;
  assign tmp8870 = ~(s10 ? tmp8871 : tmp8881);
  assign tmp8850 = s11 ? tmp8851 : tmp8870;
  assign tmp8897 = ~(l1 ? tmp8070 : tmp7955);
  assign tmp8896 = s1 ? tmp8024 : tmp8897;
  assign tmp8895 = s2 ? tmp8896 : tmp8257;
  assign tmp8899 = ~(l1 ? tmp7956 : tmp8026);
  assign tmp8898 = ~(s2 ? tmp8233 : tmp8899);
  assign tmp8894 = s3 ? tmp8895 : tmp8898;
  assign tmp8893 = s4 ? tmp8220 : tmp8894;
  assign tmp8892 = s5 ? tmp8214 : tmp8893;
  assign tmp8891 = s6 ? tmp8892 : tmp7997;
  assign tmp8890 = s7 ? tmp8211 : tmp8891;
  assign tmp8904 = s3 ? tmp8895 : tmp8258;
  assign tmp8903 = s4 ? tmp8220 : tmp8904;
  assign tmp8902 = s5 ? tmp8214 : tmp8903;
  assign tmp8901 = s6 ? tmp8250 : tmp8902;
  assign tmp8900 = s7 ? tmp8237 : tmp8901;
  assign tmp8889 = s8 ? tmp8890 : tmp8900;
  assign tmp8888 = s9 ? tmp8177 : tmp8889;
  assign tmp8908 = s6 ? tmp8263 : tmp8892;
  assign tmp8907 = s7 ? tmp8211 : tmp8908;
  assign tmp8906 = s8 ? tmp8890 : tmp8907;
  assign tmp8905 = s9 ? tmp8177 : tmp8906;
  assign tmp8887 = s10 ? tmp8888 : tmp8905;
  assign tmp8917 = s2 ? tmp8331 : tmp8358;
  assign tmp8916 = s3 ? tmp8324 : tmp8917;
  assign tmp8920 = ~(s0 ? tmp7972 : tmp8321);
  assign tmp8919 = s1 ? tmp8339 : tmp8920;
  assign tmp8918 = ~(s3 ? tmp8334 : tmp8919);
  assign tmp8915 = s4 ? tmp8916 : tmp8918;
  assign tmp8914 = s5 ? tmp8316 : tmp8915;
  assign tmp8913 = s6 ? tmp8914 : tmp7997;
  assign tmp8912 = s7 ? tmp8313 : tmp8913;
  assign tmp8924 = s4 ? tmp8916 : tmp8333;
  assign tmp8923 = s5 ? tmp8316 : tmp8924;
  assign tmp8922 = s6 ? tmp8354 : tmp8923;
  assign tmp8921 = s7 ? tmp8342 : tmp8922;
  assign tmp8911 = s8 ? tmp8912 : tmp8921;
  assign tmp8910 = s9 ? tmp8278 : tmp8911;
  assign tmp8928 = s6 ? tmp8364 : tmp8914;
  assign tmp8927 = s7 ? tmp8313 : tmp8928;
  assign tmp8926 = s8 ? tmp8912 : tmp8927;
  assign tmp8925 = s9 ? tmp8278 : tmp8926;
  assign tmp8909 = s10 ? tmp8910 : tmp8925;
  assign tmp8886 = s11 ? tmp8887 : tmp8909;
  assign tmp8849 = s12 ? tmp8850 : tmp8886;
  assign tmp8941 = s0 ? tmp8029 : tmp8428;
  assign tmp8940 = s1 ? tmp8229 : tmp8941;
  assign tmp8939 = s2 ? tmp8940 : tmp8429;
  assign tmp8942 = s2 ? tmp8430 : tmp8029;
  assign tmp8938 = ~(s3 ? tmp8939 : tmp8942);
  assign tmp8937 = s4 ? tmp8414 : tmp8938;
  assign tmp8936 = s5 ? tmp8409 : tmp8937;
  assign tmp8935 = s6 ? tmp8936 : tmp7997;
  assign tmp8934 = s7 ? tmp8405 : tmp8935;
  assign tmp8947 = ~(s3 ? tmp8939 : tmp8430);
  assign tmp8946 = s4 ? tmp8414 : tmp8947;
  assign tmp8945 = ~(s5 ? tmp8409 : tmp8946);
  assign tmp8944 = ~(s6 ? tmp8439 : tmp8945);
  assign tmp8943 = s7 ? tmp8434 : tmp8944;
  assign tmp8933 = ~(s8 ? tmp8934 : tmp8943);
  assign tmp8932 = s9 ? tmp8380 : tmp8933;
  assign tmp8952 = ~(s5 ? tmp8409 : tmp8937);
  assign tmp8951 = ~(s6 ? tmp8380 : tmp8952);
  assign tmp8950 = s7 ? tmp8405 : tmp8951;
  assign tmp8949 = ~(s8 ? tmp8934 : tmp8950);
  assign tmp8948 = s9 ? tmp8380 : tmp8949;
  assign tmp8931 = s10 ? tmp8932 : tmp8948;
  assign tmp8962 = s1 ? 1 : tmp7976;
  assign tmp8961 = s2 ? tmp8962 : tmp8063;
  assign tmp8960 = s3 ? tmp8056 : tmp8961;
  assign tmp8963 = ~(s3 ? tmp8067 : tmp8099);
  assign tmp8959 = s4 ? tmp8960 : tmp8963;
  assign tmp8958 = s5 ? tmp8046 : tmp8959;
  assign tmp8957 = s6 ? tmp8958 : tmp7997;
  assign tmp8956 = s7 ? tmp7996 : tmp8957;
  assign tmp8967 = s4 ? tmp8960 : tmp8066;
  assign tmp8966 = s5 ? tmp8046 : tmp8967;
  assign tmp8965 = s6 ? tmp8085 : tmp8966;
  assign tmp8964 = s7 ? tmp8075 : tmp8965;
  assign tmp8955 = s8 ? tmp8956 : tmp8964;
  assign tmp8954 = s9 ? tmp7951 : tmp8955;
  assign tmp8971 = s6 ? tmp8093 : tmp8958;
  assign tmp8970 = s7 ? tmp7996 : tmp8971;
  assign tmp8969 = s8 ? tmp8956 : tmp8970;
  assign tmp8968 = s9 ? tmp7951 : tmp8969;
  assign tmp8953 = ~(s10 ? tmp8954 : tmp8968);
  assign tmp8930 = s11 ? tmp8931 : tmp8953;
  assign tmp8981 = s2 ? tmp8581 : tmp8600;
  assign tmp8982 = s2 ? tmp8583 : tmp8033;
  assign tmp8980 = ~(s3 ? tmp8981 : tmp8982);
  assign tmp8979 = s4 ? tmp8570 : tmp8980;
  assign tmp8978 = s5 ? tmp8564 : tmp8979;
  assign tmp8977 = s6 ? tmp8978 : tmp7997;
  assign tmp8976 = s7 ? tmp8561 : tmp8977;
  assign tmp8987 = ~(s3 ? tmp8981 : tmp8583);
  assign tmp8986 = s4 ? tmp8570 : tmp8987;
  assign tmp8985 = s5 ? tmp8564 : tmp8986;
  assign tmp8984 = s6 ? tmp8594 : tmp8985;
  assign tmp8983 = s7 ? tmp8585 : tmp8984;
  assign tmp8975 = s8 ? tmp8976 : tmp8983;
  assign tmp8974 = s9 ? tmp8531 : tmp8975;
  assign tmp8991 = s6 ? tmp8607 : tmp8978;
  assign tmp8990 = s7 ? tmp8561 : tmp8991;
  assign tmp8989 = s8 ? tmp8976 : tmp8990;
  assign tmp8988 = s9 ? tmp8531 : tmp8989;
  assign tmp8973 = ~(s10 ? tmp8974 : tmp8988);
  assign tmp8972 = s11 ? tmp8447 : tmp8973;
  assign tmp8929 = ~(s12 ? tmp8930 : tmp8972);
  assign tmp8848 = ~(s13 ? tmp8849 : tmp8929);
  assign tmp8615 = ~(s15 ? tmp8616 : tmp8848);
  assign tmp7945 = s16 ? tmp7946 : tmp8615;
  assign s0n = tmp7945;

  initial
   begin
    s0 = 0;
    s1 = 0;
    s2 = 0;
    s3 = 0;
    s4 = 0;
    s5 = 0;
    s6 = 0;
    s7 = 0;
    s8 = 0;
    s9 = 0;
    s10 = 0;
    s11 = 0;
    s12 = 0;
    s13 = 0;
    s14 = 0;
    s15 = 0;
    s16 = 0;
   end

  always @(posedge clock)
   begin
    s0 = s0n;
    s1 = s1n;
    s2 = s2n;
    s3 = s3n;
    s4 = s4n;
    s5 = s5n;
    s6 = s6n;
    s7 = s7n;
    s8 = s8n;
    s9 = s9n;
    s10 = s10n;
    s11 = s11n;
    s12 = s12n;
    s13 = s13n;
    s14 = s14n;
    s15 = s15n;
    s16 = s16n;
   end
endmodule

